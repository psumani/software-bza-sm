// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 13 2021 17:23:46

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "zim" view "INTERFACE"

module zim (
    VAC_DRDY,
    IAC_FLT1,
    DDS_SCK,
    ICE_IOR_166,
    ICE_IOR_119,
    DDS_MOSI,
    VAC_MISO,
    DDS_MOSI1,
    ICE_IOR_146,
    VDC_CLK,
    ICE_IOT_222,
    IAC_CS,
    ICE_IOL_18B,
    ICE_IOL_13A,
    ICE_IOB_81,
    VAC_OSR1,
    IAC_MOSI,
    DDS_CS1,
    ICE_IOL_4B,
    ICE_IOB_94,
    VAC_CS,
    VAC_CLK,
    ICE_SPI_CE0,
    ICE_IOR_167,
    ICE_IOR_118,
    RTD_SDO,
    IAC_OSR0,
    VDC_SCLK,
    VAC_FLT1,
    ICE_SPI_MOSI,
    ICE_IOR_165,
    ICE_IOR_147,
    ICE_IOL_14A,
    ICE_IOL_13B,
    ICE_IOB_91,
    ICE_GPMO_0,
    DDS_RNG_0,
    VDC_RNG0,
    ICE_SPI_SCLK,
    ICE_IOR_152,
    ICE_IOL_12A,
    RTD_DRDY,
    ICE_SPI_MISO,
    ICE_IOT_177,
    ICE_IOR_141,
    ICE_IOB_80,
    ICE_IOB_102,
    ICE_GPMO_2,
    ICE_GPMI_0,
    IAC_MISO,
    VAC_OSR0,
    VAC_MOSI,
    TEST_LED,
    ICE_IOR_148,
    STAT_COMM,
    ICE_SYSCLK,
    ICE_IOR_161,
    ICE_IOB_95,
    ICE_IOB_82,
    ICE_IOB_104,
    IAC_CLK,
    DDS_CS,
    SELIRNG0,
    RTD_SDI,
    ICE_IOT_221,
    ICE_IOT_197,
    DDS_MCLK,
    RTD_SCLK,
    RTD_CS,
    ICE_IOR_137,
    IAC_OSR1,
    VAC_FLT0,
    ICE_IOR_144,
    ICE_IOR_128,
    ICE_GPMO_1,
    IAC_SCLK,
    EIS_SYNCCLK,
    ICE_IOR_139,
    ICE_IOL_4A,
    VAC_SCLK,
    THERMOSTAT,
    ICE_IOR_164,
    ICE_IOB_103,
    AMPV_POW,
    VDC_SDO,
    ICE_IOT_174,
    ICE_IOR_140,
    ICE_IOB_96,
    CONT_SD,
    AC_ADC_SYNC,
    SELIRNG1,
    ICE_IOL_12B,
    ICE_IOR_160,
    ICE_IOR_136,
    DDS_MCLK1,
    ICE_IOT_198,
    ICE_IOT_173,
    IAC_DRDY,
    ICE_IOT_178,
    ICE_IOR_138,
    ICE_IOR_120,
    IAC_FLT0,
    DDS_SCK1);

    input VAC_DRDY;
    output IAC_FLT1;
    output DDS_SCK;
    input ICE_IOR_166;
    input ICE_IOR_119;
    output DDS_MOSI;
    input VAC_MISO;
    output DDS_MOSI1;
    input ICE_IOR_146;
    output VDC_CLK;
    input ICE_IOT_222;
    output IAC_CS;
    input ICE_IOL_18B;
    input ICE_IOL_13A;
    input ICE_IOB_81;
    output VAC_OSR1;
    output IAC_MOSI;
    output DDS_CS1;
    input ICE_IOL_4B;
    input ICE_IOB_94;
    output VAC_CS;
    output VAC_CLK;
    input ICE_SPI_CE0;
    input ICE_IOR_167;
    input ICE_IOR_118;
    input RTD_SDO;
    output IAC_OSR0;
    output VDC_SCLK;
    output VAC_FLT1;
    input ICE_SPI_MOSI;
    input ICE_IOR_165;
    input ICE_IOR_147;
    input ICE_IOL_14A;
    input ICE_IOL_13B;
    input ICE_IOB_91;
    input ICE_GPMO_0;
    output DDS_RNG_0;
    output VDC_RNG0;
    input ICE_SPI_SCLK;
    input ICE_IOR_152;
    input ICE_IOL_12A;
    input RTD_DRDY;
    output ICE_SPI_MISO;
    input ICE_IOT_177;
    input ICE_IOR_141;
    input ICE_IOB_80;
    input ICE_IOB_102;
    input ICE_GPMO_2;
    output ICE_GPMI_0;
    input IAC_MISO;
    output VAC_OSR0;
    output VAC_MOSI;
    output TEST_LED;
    input ICE_IOR_148;
    output STAT_COMM;
    input ICE_SYSCLK;
    input ICE_IOR_161;
    input ICE_IOB_95;
    input ICE_IOB_82;
    input ICE_IOB_104;
    output IAC_CLK;
    output DDS_CS;
    output SELIRNG0;
    output RTD_SDI;
    input ICE_IOT_221;
    input ICE_IOT_197;
    output DDS_MCLK;
    output RTD_SCLK;
    output RTD_CS;
    input ICE_IOR_137;
    output IAC_OSR1;
    output VAC_FLT0;
    input ICE_IOR_144;
    input ICE_IOR_128;
    input ICE_GPMO_1;
    output IAC_SCLK;
    input EIS_SYNCCLK;
    input ICE_IOR_139;
    input ICE_IOL_4A;
    output VAC_SCLK;
    input THERMOSTAT;
    input ICE_IOR_164;
    input ICE_IOB_103;
    output AMPV_POW;
    input VDC_SDO;
    input ICE_IOT_174;
    input ICE_IOR_140;
    input ICE_IOB_96;
    output CONT_SD;
    output AC_ADC_SYNC;
    output SELIRNG1;
    input ICE_IOL_12B;
    input ICE_IOR_160;
    input ICE_IOR_136;
    output DDS_MCLK1;
    input ICE_IOT_198;
    input ICE_IOT_173;
    input IAC_DRDY;
    input ICE_IOT_178;
    input ICE_IOR_138;
    input ICE_IOR_120;
    output IAC_FLT0;
    output DDS_SCK1;

    wire N__65921;
    wire N__65920;
    wire N__65919;
    wire N__65912;
    wire N__65911;
    wire N__65910;
    wire N__65903;
    wire N__65902;
    wire N__65901;
    wire N__65894;
    wire N__65893;
    wire N__65892;
    wire N__65885;
    wire N__65884;
    wire N__65883;
    wire N__65876;
    wire N__65875;
    wire N__65874;
    wire N__65867;
    wire N__65866;
    wire N__65865;
    wire N__65858;
    wire N__65857;
    wire N__65856;
    wire N__65849;
    wire N__65848;
    wire N__65847;
    wire N__65840;
    wire N__65839;
    wire N__65838;
    wire N__65831;
    wire N__65830;
    wire N__65829;
    wire N__65822;
    wire N__65821;
    wire N__65820;
    wire N__65813;
    wire N__65812;
    wire N__65811;
    wire N__65804;
    wire N__65803;
    wire N__65802;
    wire N__65795;
    wire N__65794;
    wire N__65793;
    wire N__65786;
    wire N__65785;
    wire N__65784;
    wire N__65777;
    wire N__65776;
    wire N__65775;
    wire N__65768;
    wire N__65767;
    wire N__65766;
    wire N__65759;
    wire N__65758;
    wire N__65757;
    wire N__65750;
    wire N__65749;
    wire N__65748;
    wire N__65741;
    wire N__65740;
    wire N__65739;
    wire N__65732;
    wire N__65731;
    wire N__65730;
    wire N__65723;
    wire N__65722;
    wire N__65721;
    wire N__65714;
    wire N__65713;
    wire N__65712;
    wire N__65705;
    wire N__65704;
    wire N__65703;
    wire N__65696;
    wire N__65695;
    wire N__65694;
    wire N__65687;
    wire N__65686;
    wire N__65685;
    wire N__65678;
    wire N__65677;
    wire N__65676;
    wire N__65669;
    wire N__65668;
    wire N__65667;
    wire N__65660;
    wire N__65659;
    wire N__65658;
    wire N__65651;
    wire N__65650;
    wire N__65649;
    wire N__65642;
    wire N__65641;
    wire N__65640;
    wire N__65633;
    wire N__65632;
    wire N__65631;
    wire N__65624;
    wire N__65623;
    wire N__65622;
    wire N__65615;
    wire N__65614;
    wire N__65613;
    wire N__65606;
    wire N__65605;
    wire N__65604;
    wire N__65597;
    wire N__65596;
    wire N__65595;
    wire N__65588;
    wire N__65587;
    wire N__65586;
    wire N__65579;
    wire N__65578;
    wire N__65577;
    wire N__65570;
    wire N__65569;
    wire N__65568;
    wire N__65561;
    wire N__65560;
    wire N__65559;
    wire N__65552;
    wire N__65551;
    wire N__65550;
    wire N__65543;
    wire N__65542;
    wire N__65541;
    wire N__65534;
    wire N__65533;
    wire N__65532;
    wire N__65525;
    wire N__65524;
    wire N__65523;
    wire N__65516;
    wire N__65515;
    wire N__65514;
    wire N__65507;
    wire N__65506;
    wire N__65505;
    wire N__65498;
    wire N__65497;
    wire N__65496;
    wire N__65489;
    wire N__65488;
    wire N__65487;
    wire N__65480;
    wire N__65479;
    wire N__65478;
    wire N__65471;
    wire N__65470;
    wire N__65469;
    wire N__65462;
    wire N__65461;
    wire N__65460;
    wire N__65453;
    wire N__65452;
    wire N__65451;
    wire N__65444;
    wire N__65443;
    wire N__65442;
    wire N__65435;
    wire N__65434;
    wire N__65433;
    wire N__65426;
    wire N__65425;
    wire N__65424;
    wire N__65417;
    wire N__65416;
    wire N__65415;
    wire N__65408;
    wire N__65407;
    wire N__65406;
    wire N__65399;
    wire N__65398;
    wire N__65397;
    wire N__65390;
    wire N__65389;
    wire N__65388;
    wire N__65381;
    wire N__65380;
    wire N__65379;
    wire N__65372;
    wire N__65371;
    wire N__65370;
    wire N__65363;
    wire N__65362;
    wire N__65361;
    wire N__65354;
    wire N__65353;
    wire N__65352;
    wire N__65345;
    wire N__65344;
    wire N__65343;
    wire N__65336;
    wire N__65335;
    wire N__65334;
    wire N__65327;
    wire N__65326;
    wire N__65325;
    wire N__65318;
    wire N__65317;
    wire N__65316;
    wire N__65309;
    wire N__65308;
    wire N__65307;
    wire N__65300;
    wire N__65299;
    wire N__65298;
    wire N__65291;
    wire N__65290;
    wire N__65289;
    wire N__65282;
    wire N__65281;
    wire N__65280;
    wire N__65273;
    wire N__65272;
    wire N__65271;
    wire N__65264;
    wire N__65263;
    wire N__65262;
    wire N__65255;
    wire N__65254;
    wire N__65253;
    wire N__65246;
    wire N__65245;
    wire N__65244;
    wire N__65237;
    wire N__65236;
    wire N__65235;
    wire N__65228;
    wire N__65227;
    wire N__65226;
    wire N__65219;
    wire N__65218;
    wire N__65217;
    wire N__65210;
    wire N__65209;
    wire N__65208;
    wire N__65201;
    wire N__65200;
    wire N__65199;
    wire N__65192;
    wire N__65191;
    wire N__65190;
    wire N__65183;
    wire N__65182;
    wire N__65181;
    wire N__65174;
    wire N__65173;
    wire N__65172;
    wire N__65165;
    wire N__65164;
    wire N__65163;
    wire N__65156;
    wire N__65155;
    wire N__65154;
    wire N__65147;
    wire N__65146;
    wire N__65145;
    wire N__65138;
    wire N__65137;
    wire N__65136;
    wire N__65129;
    wire N__65128;
    wire N__65127;
    wire N__65120;
    wire N__65119;
    wire N__65118;
    wire N__65111;
    wire N__65110;
    wire N__65109;
    wire N__65102;
    wire N__65101;
    wire N__65100;
    wire N__65093;
    wire N__65092;
    wire N__65091;
    wire N__65084;
    wire N__65083;
    wire N__65082;
    wire N__65075;
    wire N__65074;
    wire N__65073;
    wire N__65066;
    wire N__65065;
    wire N__65064;
    wire N__65057;
    wire N__65056;
    wire N__65055;
    wire N__65048;
    wire N__65047;
    wire N__65046;
    wire N__65039;
    wire N__65038;
    wire N__65037;
    wire N__65030;
    wire N__65029;
    wire N__65028;
    wire N__65021;
    wire N__65020;
    wire N__65019;
    wire N__65012;
    wire N__65011;
    wire N__65010;
    wire N__65003;
    wire N__65002;
    wire N__65001;
    wire N__64984;
    wire N__64981;
    wire N__64980;
    wire N__64977;
    wire N__64974;
    wire N__64971;
    wire N__64966;
    wire N__64963;
    wire N__64962;
    wire N__64959;
    wire N__64956;
    wire N__64951;
    wire N__64948;
    wire N__64947;
    wire N__64944;
    wire N__64941;
    wire N__64936;
    wire N__64933;
    wire N__64932;
    wire N__64929;
    wire N__64926;
    wire N__64921;
    wire N__64918;
    wire N__64917;
    wire N__64914;
    wire N__64911;
    wire N__64906;
    wire N__64903;
    wire N__64902;
    wire N__64899;
    wire N__64896;
    wire N__64891;
    wire N__64888;
    wire N__64887;
    wire N__64884;
    wire N__64881;
    wire N__64876;
    wire N__64873;
    wire N__64870;
    wire N__64869;
    wire N__64868;
    wire N__64865;
    wire N__64862;
    wire N__64859;
    wire N__64858;
    wire N__64857;
    wire N__64856;
    wire N__64855;
    wire N__64854;
    wire N__64853;
    wire N__64852;
    wire N__64851;
    wire N__64850;
    wire N__64849;
    wire N__64848;
    wire N__64847;
    wire N__64846;
    wire N__64845;
    wire N__64844;
    wire N__64841;
    wire N__64836;
    wire N__64833;
    wire N__64830;
    wire N__64829;
    wire N__64828;
    wire N__64825;
    wire N__64824;
    wire N__64823;
    wire N__64820;
    wire N__64819;
    wire N__64816;
    wire N__64815;
    wire N__64812;
    wire N__64811;
    wire N__64808;
    wire N__64807;
    wire N__64804;
    wire N__64803;
    wire N__64800;
    wire N__64799;
    wire N__64796;
    wire N__64795;
    wire N__64792;
    wire N__64789;
    wire N__64788;
    wire N__64785;
    wire N__64784;
    wire N__64781;
    wire N__64780;
    wire N__64777;
    wire N__64774;
    wire N__64767;
    wire N__64764;
    wire N__64761;
    wire N__64758;
    wire N__64755;
    wire N__64752;
    wire N__64749;
    wire N__64734;
    wire N__64733;
    wire N__64732;
    wire N__64731;
    wire N__64730;
    wire N__64729;
    wire N__64728;
    wire N__64727;
    wire N__64712;
    wire N__64697;
    wire N__64696;
    wire N__64695;
    wire N__64694;
    wire N__64693;
    wire N__64684;
    wire N__64677;
    wire N__64676;
    wire N__64673;
    wire N__64670;
    wire N__64667;
    wire N__64666;
    wire N__64663;
    wire N__64660;
    wire N__64657;
    wire N__64654;
    wire N__64651;
    wire N__64648;
    wire N__64645;
    wire N__64642;
    wire N__64641;
    wire N__64638;
    wire N__64637;
    wire N__64634;
    wire N__64633;
    wire N__64630;
    wire N__64629;
    wire N__64626;
    wire N__64621;
    wire N__64618;
    wire N__64617;
    wire N__64616;
    wire N__64613;
    wire N__64610;
    wire N__64601;
    wire N__64592;
    wire N__64587;
    wire N__64570;
    wire N__64567;
    wire N__64564;
    wire N__64561;
    wire N__64558;
    wire N__64557;
    wire N__64554;
    wire N__64551;
    wire N__64542;
    wire N__64537;
    wire N__64534;
    wire N__64531;
    wire N__64528;
    wire N__64521;
    wire N__64518;
    wire N__64513;
    wire N__64510;
    wire N__64501;
    wire N__64498;
    wire N__64497;
    wire N__64494;
    wire N__64491;
    wire N__64488;
    wire N__64483;
    wire N__64480;
    wire N__64479;
    wire N__64476;
    wire N__64473;
    wire N__64470;
    wire N__64467;
    wire N__64462;
    wire N__64459;
    wire N__64458;
    wire N__64457;
    wire N__64454;
    wire N__64451;
    wire N__64448;
    wire N__64447;
    wire N__64444;
    wire N__64441;
    wire N__64438;
    wire N__64435;
    wire N__64432;
    wire N__64427;
    wire N__64424;
    wire N__64417;
    wire N__64416;
    wire N__64413;
    wire N__64410;
    wire N__64407;
    wire N__64404;
    wire N__64401;
    wire N__64398;
    wire N__64393;
    wire N__64392;
    wire N__64389;
    wire N__64386;
    wire N__64381;
    wire N__64378;
    wire N__64377;
    wire N__64374;
    wire N__64371;
    wire N__64366;
    wire N__64363;
    wire N__64360;
    wire N__64359;
    wire N__64356;
    wire N__64353;
    wire N__64348;
    wire N__64345;
    wire N__64342;
    wire N__64341;
    wire N__64338;
    wire N__64335;
    wire N__64330;
    wire N__64327;
    wire N__64326;
    wire N__64323;
    wire N__64320;
    wire N__64317;
    wire N__64314;
    wire N__64311;
    wire N__64306;
    wire N__64303;
    wire N__64302;
    wire N__64299;
    wire N__64296;
    wire N__64291;
    wire N__64288;
    wire N__64285;
    wire N__64284;
    wire N__64281;
    wire N__64278;
    wire N__64273;
    wire N__64270;
    wire N__64269;
    wire N__64266;
    wire N__64263;
    wire N__64260;
    wire N__64255;
    wire N__64252;
    wire N__64249;
    wire N__64246;
    wire N__64243;
    wire N__64240;
    wire N__64237;
    wire N__64234;
    wire N__64231;
    wire N__64228;
    wire N__64227;
    wire N__64224;
    wire N__64221;
    wire N__64220;
    wire N__64219;
    wire N__64218;
    wire N__64217;
    wire N__64216;
    wire N__64211;
    wire N__64206;
    wire N__64203;
    wire N__64198;
    wire N__64189;
    wire N__64186;
    wire N__64183;
    wire N__64180;
    wire N__64179;
    wire N__64176;
    wire N__64173;
    wire N__64168;
    wire N__64167;
    wire N__64164;
    wire N__64163;
    wire N__64162;
    wire N__64161;
    wire N__64154;
    wire N__64151;
    wire N__64148;
    wire N__64143;
    wire N__64138;
    wire N__64135;
    wire N__64132;
    wire N__64129;
    wire N__64126;
    wire N__64123;
    wire N__64120;
    wire N__64117;
    wire N__64114;
    wire N__64111;
    wire N__64110;
    wire N__64109;
    wire N__64102;
    wire N__64101;
    wire N__64098;
    wire N__64097;
    wire N__64096;
    wire N__64095;
    wire N__64092;
    wire N__64091;
    wire N__64090;
    wire N__64089;
    wire N__64088;
    wire N__64085;
    wire N__64080;
    wire N__64079;
    wire N__64078;
    wire N__64077;
    wire N__64076;
    wire N__64067;
    wire N__64066;
    wire N__64065;
    wire N__64062;
    wire N__64059;
    wire N__64054;
    wire N__64051;
    wire N__64050;
    wire N__64049;
    wire N__64048;
    wire N__64041;
    wire N__64038;
    wire N__64035;
    wire N__64034;
    wire N__64033;
    wire N__64032;
    wire N__64031;
    wire N__64030;
    wire N__64029;
    wire N__64026;
    wire N__64025;
    wire N__64024;
    wire N__64023;
    wire N__64022;
    wire N__64017;
    wire N__64012;
    wire N__64011;
    wire N__64008;
    wire N__64007;
    wire N__64006;
    wire N__64001;
    wire N__63998;
    wire N__63995;
    wire N__63994;
    wire N__63993;
    wire N__63992;
    wire N__63991;
    wire N__63990;
    wire N__63989;
    wire N__63988;
    wire N__63987;
    wire N__63986;
    wire N__63985;
    wire N__63980;
    wire N__63973;
    wire N__63970;
    wire N__63967;
    wire N__63966;
    wire N__63963;
    wire N__63960;
    wire N__63959;
    wire N__63956;
    wire N__63951;
    wire N__63946;
    wire N__63941;
    wire N__63936;
    wire N__63931;
    wire N__63928;
    wire N__63923;
    wire N__63920;
    wire N__63911;
    wire N__63910;
    wire N__63909;
    wire N__63908;
    wire N__63905;
    wire N__63902;
    wire N__63899;
    wire N__63896;
    wire N__63893;
    wire N__63890;
    wire N__63889;
    wire N__63888;
    wire N__63885;
    wire N__63882;
    wire N__63879;
    wire N__63876;
    wire N__63873;
    wire N__63868;
    wire N__63865;
    wire N__63860;
    wire N__63853;
    wire N__63848;
    wire N__63845;
    wire N__63836;
    wire N__63827;
    wire N__63822;
    wire N__63815;
    wire N__63802;
    wire N__63799;
    wire N__63784;
    wire N__63783;
    wire N__63782;
    wire N__63781;
    wire N__63780;
    wire N__63779;
    wire N__63778;
    wire N__63777;
    wire N__63774;
    wire N__63771;
    wire N__63770;
    wire N__63769;
    wire N__63768;
    wire N__63767;
    wire N__63766;
    wire N__63765;
    wire N__63764;
    wire N__63763;
    wire N__63762;
    wire N__63761;
    wire N__63760;
    wire N__63757;
    wire N__63756;
    wire N__63753;
    wire N__63752;
    wire N__63749;
    wire N__63748;
    wire N__63745;
    wire N__63744;
    wire N__63743;
    wire N__63742;
    wire N__63741;
    wire N__63740;
    wire N__63739;
    wire N__63738;
    wire N__63737;
    wire N__63736;
    wire N__63735;
    wire N__63732;
    wire N__63727;
    wire N__63726;
    wire N__63725;
    wire N__63724;
    wire N__63723;
    wire N__63722;
    wire N__63719;
    wire N__63718;
    wire N__63717;
    wire N__63714;
    wire N__63711;
    wire N__63708;
    wire N__63705;
    wire N__63702;
    wire N__63699;
    wire N__63696;
    wire N__63693;
    wire N__63690;
    wire N__63687;
    wire N__63670;
    wire N__63667;
    wire N__63656;
    wire N__63655;
    wire N__63654;
    wire N__63651;
    wire N__63650;
    wire N__63649;
    wire N__63648;
    wire N__63645;
    wire N__63644;
    wire N__63643;
    wire N__63642;
    wire N__63637;
    wire N__63634;
    wire N__63631;
    wire N__63628;
    wire N__63625;
    wire N__63622;
    wire N__63619;
    wire N__63618;
    wire N__63617;
    wire N__63614;
    wire N__63613;
    wire N__63612;
    wire N__63611;
    wire N__63610;
    wire N__63609;
    wire N__63608;
    wire N__63607;
    wire N__63606;
    wire N__63605;
    wire N__63604;
    wire N__63603;
    wire N__63602;
    wire N__63601;
    wire N__63598;
    wire N__63597;
    wire N__63596;
    wire N__63595;
    wire N__63594;
    wire N__63589;
    wire N__63580;
    wire N__63571;
    wire N__63568;
    wire N__63559;
    wire N__63554;
    wire N__63551;
    wire N__63548;
    wire N__63545;
    wire N__63542;
    wire N__63541;
    wire N__63540;
    wire N__63539;
    wire N__63536;
    wire N__63529;
    wire N__63528;
    wire N__63527;
    wire N__63526;
    wire N__63525;
    wire N__63514;
    wire N__63511;
    wire N__63506;
    wire N__63505;
    wire N__63504;
    wire N__63501;
    wire N__63498;
    wire N__63495;
    wire N__63494;
    wire N__63493;
    wire N__63492;
    wire N__63491;
    wire N__63490;
    wire N__63489;
    wire N__63488;
    wire N__63487;
    wire N__63486;
    wire N__63485;
    wire N__63484;
    wire N__63483;
    wire N__63482;
    wire N__63479;
    wire N__63474;
    wire N__63469;
    wire N__63466;
    wire N__63457;
    wire N__63454;
    wire N__63451;
    wire N__63448;
    wire N__63445;
    wire N__63438;
    wire N__63421;
    wire N__63418;
    wire N__63415;
    wire N__63412;
    wire N__63407;
    wire N__63402;
    wire N__63397;
    wire N__63394;
    wire N__63393;
    wire N__63390;
    wire N__63383;
    wire N__63382;
    wire N__63381;
    wire N__63380;
    wire N__63379;
    wire N__63378;
    wire N__63373;
    wire N__63366;
    wire N__63359;
    wire N__63358;
    wire N__63357;
    wire N__63354;
    wire N__63349;
    wire N__63346;
    wire N__63341;
    wire N__63338;
    wire N__63331;
    wire N__63320;
    wire N__63317;
    wire N__63314;
    wire N__63305;
    wire N__63300;
    wire N__63291;
    wire N__63288;
    wire N__63285;
    wire N__63282;
    wire N__63279;
    wire N__63270;
    wire N__63267;
    wire N__63260;
    wire N__63255;
    wire N__63240;
    wire N__63229;
    wire N__63218;
    wire N__63205;
    wire N__63204;
    wire N__63201;
    wire N__63200;
    wire N__63197;
    wire N__63196;
    wire N__63195;
    wire N__63194;
    wire N__63191;
    wire N__63190;
    wire N__63189;
    wire N__63188;
    wire N__63185;
    wire N__63182;
    wire N__63177;
    wire N__63174;
    wire N__63173;
    wire N__63170;
    wire N__63167;
    wire N__63164;
    wire N__63163;
    wire N__63162;
    wire N__63157;
    wire N__63152;
    wire N__63149;
    wire N__63146;
    wire N__63145;
    wire N__63140;
    wire N__63133;
    wire N__63128;
    wire N__63125;
    wire N__63122;
    wire N__63119;
    wire N__63114;
    wire N__63111;
    wire N__63110;
    wire N__63105;
    wire N__63100;
    wire N__63097;
    wire N__63094;
    wire N__63085;
    wire N__63084;
    wire N__63083;
    wire N__63082;
    wire N__63081;
    wire N__63080;
    wire N__63079;
    wire N__63078;
    wire N__63077;
    wire N__63076;
    wire N__63075;
    wire N__63074;
    wire N__63073;
    wire N__63072;
    wire N__63071;
    wire N__63070;
    wire N__63067;
    wire N__63066;
    wire N__63061;
    wire N__63060;
    wire N__63059;
    wire N__63058;
    wire N__63057;
    wire N__63056;
    wire N__63055;
    wire N__63052;
    wire N__63051;
    wire N__63050;
    wire N__63049;
    wire N__63048;
    wire N__63047;
    wire N__63046;
    wire N__63045;
    wire N__63042;
    wire N__63039;
    wire N__63034;
    wire N__63031;
    wire N__63030;
    wire N__63029;
    wire N__63028;
    wire N__63027;
    wire N__63024;
    wire N__63021;
    wire N__63018;
    wire N__63015;
    wire N__63012;
    wire N__63003;
    wire N__63000;
    wire N__62991;
    wire N__62986;
    wire N__62983;
    wire N__62980;
    wire N__62973;
    wire N__62970;
    wire N__62969;
    wire N__62964;
    wire N__62957;
    wire N__62954;
    wire N__62949;
    wire N__62944;
    wire N__62943;
    wire N__62940;
    wire N__62937;
    wire N__62936;
    wire N__62935;
    wire N__62934;
    wire N__62933;
    wire N__62932;
    wire N__62931;
    wire N__62930;
    wire N__62927;
    wire N__62924;
    wire N__62913;
    wire N__62908;
    wire N__62907;
    wire N__62906;
    wire N__62905;
    wire N__62902;
    wire N__62899;
    wire N__62896;
    wire N__62891;
    wire N__62884;
    wire N__62881;
    wire N__62878;
    wire N__62875;
    wire N__62872;
    wire N__62863;
    wire N__62858;
    wire N__62849;
    wire N__62844;
    wire N__62841;
    wire N__62836;
    wire N__62831;
    wire N__62822;
    wire N__62803;
    wire N__62800;
    wire N__62797;
    wire N__62794;
    wire N__62791;
    wire N__62790;
    wire N__62789;
    wire N__62788;
    wire N__62785;
    wire N__62784;
    wire N__62781;
    wire N__62780;
    wire N__62779;
    wire N__62776;
    wire N__62775;
    wire N__62772;
    wire N__62769;
    wire N__62766;
    wire N__62763;
    wire N__62760;
    wire N__62757;
    wire N__62754;
    wire N__62751;
    wire N__62748;
    wire N__62743;
    wire N__62740;
    wire N__62737;
    wire N__62734;
    wire N__62731;
    wire N__62728;
    wire N__62727;
    wire N__62724;
    wire N__62721;
    wire N__62716;
    wire N__62713;
    wire N__62708;
    wire N__62705;
    wire N__62692;
    wire N__62691;
    wire N__62690;
    wire N__62689;
    wire N__62686;
    wire N__62685;
    wire N__62682;
    wire N__62679;
    wire N__62678;
    wire N__62677;
    wire N__62676;
    wire N__62675;
    wire N__62674;
    wire N__62673;
    wire N__62672;
    wire N__62671;
    wire N__62670;
    wire N__62667;
    wire N__62664;
    wire N__62663;
    wire N__62662;
    wire N__62661;
    wire N__62660;
    wire N__62659;
    wire N__62658;
    wire N__62657;
    wire N__62656;
    wire N__62655;
    wire N__62654;
    wire N__62653;
    wire N__62652;
    wire N__62649;
    wire N__62648;
    wire N__62647;
    wire N__62646;
    wire N__62645;
    wire N__62638;
    wire N__62637;
    wire N__62634;
    wire N__62633;
    wire N__62632;
    wire N__62631;
    wire N__62630;
    wire N__62629;
    wire N__62628;
    wire N__62627;
    wire N__62626;
    wire N__62625;
    wire N__62624;
    wire N__62623;
    wire N__62622;
    wire N__62621;
    wire N__62620;
    wire N__62619;
    wire N__62618;
    wire N__62617;
    wire N__62616;
    wire N__62615;
    wire N__62612;
    wire N__62611;
    wire N__62610;
    wire N__62609;
    wire N__62608;
    wire N__62607;
    wire N__62606;
    wire N__62605;
    wire N__62604;
    wire N__62603;
    wire N__62602;
    wire N__62601;
    wire N__62600;
    wire N__62599;
    wire N__62598;
    wire N__62597;
    wire N__62596;
    wire N__62595;
    wire N__62588;
    wire N__62585;
    wire N__62582;
    wire N__62579;
    wire N__62576;
    wire N__62573;
    wire N__62572;
    wire N__62571;
    wire N__62570;
    wire N__62569;
    wire N__62568;
    wire N__62567;
    wire N__62566;
    wire N__62565;
    wire N__62564;
    wire N__62561;
    wire N__62548;
    wire N__62531;
    wire N__62530;
    wire N__62529;
    wire N__62528;
    wire N__62527;
    wire N__62526;
    wire N__62525;
    wire N__62524;
    wire N__62523;
    wire N__62522;
    wire N__62521;
    wire N__62516;
    wire N__62513;
    wire N__62510;
    wire N__62507;
    wire N__62504;
    wire N__62487;
    wire N__62486;
    wire N__62485;
    wire N__62482;
    wire N__62481;
    wire N__62480;
    wire N__62463;
    wire N__62460;
    wire N__62451;
    wire N__62450;
    wire N__62449;
    wire N__62446;
    wire N__62443;
    wire N__62440;
    wire N__62435;
    wire N__62432;
    wire N__62429;
    wire N__62428;
    wire N__62427;
    wire N__62426;
    wire N__62423;
    wire N__62422;
    wire N__62421;
    wire N__62418;
    wire N__62411;
    wire N__62406;
    wire N__62403;
    wire N__62392;
    wire N__62385;
    wire N__62380;
    wire N__62373;
    wire N__62370;
    wire N__62369;
    wire N__62368;
    wire N__62361;
    wire N__62358;
    wire N__62355;
    wire N__62338;
    wire N__62335;
    wire N__62332;
    wire N__62327;
    wire N__62324;
    wire N__62321;
    wire N__62316;
    wire N__62313;
    wire N__62308;
    wire N__62301;
    wire N__62298;
    wire N__62297;
    wire N__62296;
    wire N__62295;
    wire N__62294;
    wire N__62293;
    wire N__62292;
    wire N__62291;
    wire N__62290;
    wire N__62285;
    wire N__62276;
    wire N__62273;
    wire N__62260;
    wire N__62243;
    wire N__62242;
    wire N__62241;
    wire N__62240;
    wire N__62237;
    wire N__62232;
    wire N__62227;
    wire N__62218;
    wire N__62215;
    wire N__62212;
    wire N__62205;
    wire N__62200;
    wire N__62197;
    wire N__62192;
    wire N__62187;
    wire N__62184;
    wire N__62179;
    wire N__62176;
    wire N__62171;
    wire N__62164;
    wire N__62157;
    wire N__62154;
    wire N__62145;
    wire N__62138;
    wire N__62113;
    wire N__62110;
    wire N__62107;
    wire N__62104;
    wire N__62101;
    wire N__62100;
    wire N__62097;
    wire N__62094;
    wire N__62093;
    wire N__62092;
    wire N__62087;
    wire N__62086;
    wire N__62083;
    wire N__62080;
    wire N__62079;
    wire N__62076;
    wire N__62073;
    wire N__62070;
    wire N__62065;
    wire N__62060;
    wire N__62057;
    wire N__62056;
    wire N__62053;
    wire N__62050;
    wire N__62047;
    wire N__62044;
    wire N__62041;
    wire N__62038;
    wire N__62033;
    wire N__62030;
    wire N__62025;
    wire N__62022;
    wire N__62019;
    wire N__62014;
    wire N__62013;
    wire N__62012;
    wire N__62011;
    wire N__62010;
    wire N__62009;
    wire N__62008;
    wire N__62007;
    wire N__62006;
    wire N__62005;
    wire N__62004;
    wire N__62003;
    wire N__62002;
    wire N__62001;
    wire N__62000;
    wire N__61999;
    wire N__61998;
    wire N__61997;
    wire N__61996;
    wire N__61995;
    wire N__61994;
    wire N__61993;
    wire N__61992;
    wire N__61991;
    wire N__61990;
    wire N__61989;
    wire N__61988;
    wire N__61987;
    wire N__61986;
    wire N__61985;
    wire N__61984;
    wire N__61983;
    wire N__61982;
    wire N__61981;
    wire N__61980;
    wire N__61979;
    wire N__61978;
    wire N__61977;
    wire N__61976;
    wire N__61975;
    wire N__61974;
    wire N__61973;
    wire N__61972;
    wire N__61971;
    wire N__61970;
    wire N__61969;
    wire N__61968;
    wire N__61967;
    wire N__61966;
    wire N__61965;
    wire N__61964;
    wire N__61963;
    wire N__61962;
    wire N__61961;
    wire N__61960;
    wire N__61959;
    wire N__61958;
    wire N__61957;
    wire N__61956;
    wire N__61955;
    wire N__61954;
    wire N__61953;
    wire N__61952;
    wire N__61951;
    wire N__61950;
    wire N__61949;
    wire N__61948;
    wire N__61947;
    wire N__61946;
    wire N__61945;
    wire N__61944;
    wire N__61943;
    wire N__61942;
    wire N__61941;
    wire N__61940;
    wire N__61939;
    wire N__61938;
    wire N__61937;
    wire N__61936;
    wire N__61935;
    wire N__61934;
    wire N__61933;
    wire N__61932;
    wire N__61931;
    wire N__61930;
    wire N__61929;
    wire N__61928;
    wire N__61927;
    wire N__61926;
    wire N__61925;
    wire N__61924;
    wire N__61923;
    wire N__61922;
    wire N__61921;
    wire N__61920;
    wire N__61919;
    wire N__61918;
    wire N__61917;
    wire N__61916;
    wire N__61915;
    wire N__61914;
    wire N__61913;
    wire N__61912;
    wire N__61911;
    wire N__61910;
    wire N__61909;
    wire N__61908;
    wire N__61907;
    wire N__61906;
    wire N__61905;
    wire N__61904;
    wire N__61903;
    wire N__61902;
    wire N__61901;
    wire N__61900;
    wire N__61899;
    wire N__61898;
    wire N__61897;
    wire N__61896;
    wire N__61895;
    wire N__61894;
    wire N__61893;
    wire N__61892;
    wire N__61891;
    wire N__61890;
    wire N__61889;
    wire N__61888;
    wire N__61887;
    wire N__61886;
    wire N__61885;
    wire N__61884;
    wire N__61883;
    wire N__61882;
    wire N__61881;
    wire N__61880;
    wire N__61879;
    wire N__61878;
    wire N__61877;
    wire N__61876;
    wire N__61875;
    wire N__61874;
    wire N__61873;
    wire N__61872;
    wire N__61871;
    wire N__61870;
    wire N__61869;
    wire N__61868;
    wire N__61867;
    wire N__61866;
    wire N__61865;
    wire N__61864;
    wire N__61863;
    wire N__61862;
    wire N__61861;
    wire N__61860;
    wire N__61859;
    wire N__61858;
    wire N__61857;
    wire N__61856;
    wire N__61855;
    wire N__61854;
    wire N__61853;
    wire N__61852;
    wire N__61851;
    wire N__61850;
    wire N__61849;
    wire N__61848;
    wire N__61847;
    wire N__61846;
    wire N__61845;
    wire N__61844;
    wire N__61843;
    wire N__61842;
    wire N__61841;
    wire N__61840;
    wire N__61839;
    wire N__61838;
    wire N__61837;
    wire N__61836;
    wire N__61835;
    wire N__61834;
    wire N__61833;
    wire N__61832;
    wire N__61831;
    wire N__61830;
    wire N__61829;
    wire N__61828;
    wire N__61827;
    wire N__61826;
    wire N__61825;
    wire N__61824;
    wire N__61441;
    wire N__61438;
    wire N__61437;
    wire N__61434;
    wire N__61431;
    wire N__61428;
    wire N__61425;
    wire N__61420;
    wire N__61417;
    wire N__61414;
    wire N__61413;
    wire N__61412;
    wire N__61411;
    wire N__61410;
    wire N__61409;
    wire N__61408;
    wire N__61407;
    wire N__61406;
    wire N__61405;
    wire N__61402;
    wire N__61401;
    wire N__61400;
    wire N__61399;
    wire N__61398;
    wire N__61397;
    wire N__61396;
    wire N__61395;
    wire N__61394;
    wire N__61391;
    wire N__61390;
    wire N__61387;
    wire N__61384;
    wire N__61383;
    wire N__61382;
    wire N__61381;
    wire N__61380;
    wire N__61379;
    wire N__61376;
    wire N__61375;
    wire N__61374;
    wire N__61373;
    wire N__61370;
    wire N__61367;
    wire N__61364;
    wire N__61363;
    wire N__61362;
    wire N__61359;
    wire N__61356;
    wire N__61353;
    wire N__61352;
    wire N__61349;
    wire N__61348;
    wire N__61347;
    wire N__61344;
    wire N__61339;
    wire N__61336;
    wire N__61333;
    wire N__61330;
    wire N__61327;
    wire N__61322;
    wire N__61319;
    wire N__61316;
    wire N__61313;
    wire N__61310;
    wire N__61307;
    wire N__61304;
    wire N__61301;
    wire N__61300;
    wire N__61297;
    wire N__61292;
    wire N__61291;
    wire N__61288;
    wire N__61281;
    wire N__61276;
    wire N__61269;
    wire N__61268;
    wire N__61267;
    wire N__61264;
    wire N__61261;
    wire N__61260;
    wire N__61255;
    wire N__61254;
    wire N__61253;
    wire N__61248;
    wire N__61245;
    wire N__61242;
    wire N__61233;
    wire N__61232;
    wire N__61231;
    wire N__61226;
    wire N__61223;
    wire N__61218;
    wire N__61215;
    wire N__61212;
    wire N__61207;
    wire N__61204;
    wire N__61201;
    wire N__61194;
    wire N__61189;
    wire N__61184;
    wire N__61183;
    wire N__61182;
    wire N__61179;
    wire N__61178;
    wire N__61175;
    wire N__61172;
    wire N__61169;
    wire N__61160;
    wire N__61157;
    wire N__61154;
    wire N__61141;
    wire N__61130;
    wire N__61121;
    wire N__61102;
    wire N__61099;
    wire N__61096;
    wire N__61095;
    wire N__61092;
    wire N__61089;
    wire N__61086;
    wire N__61083;
    wire N__61080;
    wire N__61075;
    wire N__61072;
    wire N__61069;
    wire N__61066;
    wire N__61063;
    wire N__61060;
    wire N__61057;
    wire N__61056;
    wire N__61055;
    wire N__61054;
    wire N__61053;
    wire N__61052;
    wire N__61051;
    wire N__61048;
    wire N__61045;
    wire N__61042;
    wire N__61037;
    wire N__61036;
    wire N__61035;
    wire N__61034;
    wire N__61033;
    wire N__61032;
    wire N__61029;
    wire N__61026;
    wire N__61025;
    wire N__61024;
    wire N__61023;
    wire N__61022;
    wire N__61021;
    wire N__61020;
    wire N__61019;
    wire N__61018;
    wire N__61017;
    wire N__61014;
    wire N__61013;
    wire N__61010;
    wire N__61007;
    wire N__61004;
    wire N__60995;
    wire N__60994;
    wire N__60993;
    wire N__60992;
    wire N__60991;
    wire N__60990;
    wire N__60989;
    wire N__60986;
    wire N__60981;
    wire N__60980;
    wire N__60979;
    wire N__60978;
    wire N__60977;
    wire N__60976;
    wire N__60975;
    wire N__60970;
    wire N__60963;
    wire N__60958;
    wire N__60957;
    wire N__60956;
    wire N__60955;
    wire N__60954;
    wire N__60953;
    wire N__60952;
    wire N__60949;
    wire N__60948;
    wire N__60945;
    wire N__60942;
    wire N__60939;
    wire N__60932;
    wire N__60929;
    wire N__60926;
    wire N__60921;
    wire N__60918;
    wire N__60915;
    wire N__60912;
    wire N__60909;
    wire N__60906;
    wire N__60903;
    wire N__60902;
    wire N__60899;
    wire N__60894;
    wire N__60889;
    wire N__60884;
    wire N__60881;
    wire N__60880;
    wire N__60879;
    wire N__60876;
    wire N__60871;
    wire N__60866;
    wire N__60865;
    wire N__60862;
    wire N__60859;
    wire N__60856;
    wire N__60853;
    wire N__60850;
    wire N__60847;
    wire N__60842;
    wire N__60837;
    wire N__60834;
    wire N__60831;
    wire N__60822;
    wire N__60819;
    wire N__60810;
    wire N__60807;
    wire N__60804;
    wire N__60801;
    wire N__60794;
    wire N__60793;
    wire N__60792;
    wire N__60789;
    wire N__60786;
    wire N__60781;
    wire N__60778;
    wire N__60775;
    wire N__60770;
    wire N__60757;
    wire N__60750;
    wire N__60747;
    wire N__60742;
    wire N__60721;
    wire N__60718;
    wire N__60715;
    wire N__60712;
    wire N__60709;
    wire N__60706;
    wire N__60703;
    wire N__60700;
    wire N__60697;
    wire N__60694;
    wire N__60691;
    wire N__60690;
    wire N__60689;
    wire N__60686;
    wire N__60681;
    wire N__60676;
    wire N__60673;
    wire N__60670;
    wire N__60669;
    wire N__60668;
    wire N__60667;
    wire N__60666;
    wire N__60665;
    wire N__60664;
    wire N__60663;
    wire N__60660;
    wire N__60657;
    wire N__60650;
    wire N__60649;
    wire N__60648;
    wire N__60647;
    wire N__60646;
    wire N__60643;
    wire N__60642;
    wire N__60641;
    wire N__60640;
    wire N__60637;
    wire N__60636;
    wire N__60635;
    wire N__60632;
    wire N__60631;
    wire N__60628;
    wire N__60627;
    wire N__60624;
    wire N__60621;
    wire N__60620;
    wire N__60619;
    wire N__60616;
    wire N__60615;
    wire N__60612;
    wire N__60611;
    wire N__60610;
    wire N__60609;
    wire N__60604;
    wire N__60603;
    wire N__60602;
    wire N__60601;
    wire N__60600;
    wire N__60599;
    wire N__60598;
    wire N__60597;
    wire N__60596;
    wire N__60595;
    wire N__60594;
    wire N__60593;
    wire N__60592;
    wire N__60591;
    wire N__60590;
    wire N__60589;
    wire N__60588;
    wire N__60587;
    wire N__60584;
    wire N__60579;
    wire N__60576;
    wire N__60573;
    wire N__60568;
    wire N__60565;
    wire N__60564;
    wire N__60561;
    wire N__60558;
    wire N__60555;
    wire N__60550;
    wire N__60547;
    wire N__60546;
    wire N__60545;
    wire N__60544;
    wire N__60543;
    wire N__60540;
    wire N__60537;
    wire N__60534;
    wire N__60531;
    wire N__60528;
    wire N__60523;
    wire N__60522;
    wire N__60521;
    wire N__60520;
    wire N__60519;
    wire N__60518;
    wire N__60517;
    wire N__60516;
    wire N__60513;
    wire N__60510;
    wire N__60507;
    wire N__60502;
    wire N__60501;
    wire N__60500;
    wire N__60499;
    wire N__60498;
    wire N__60497;
    wire N__60496;
    wire N__60495;
    wire N__60490;
    wire N__60487;
    wire N__60480;
    wire N__60479;
    wire N__60478;
    wire N__60475;
    wire N__60470;
    wire N__60469;
    wire N__60468;
    wire N__60467;
    wire N__60464;
    wire N__60463;
    wire N__60462;
    wire N__60461;
    wire N__60458;
    wire N__60453;
    wire N__60446;
    wire N__60439;
    wire N__60436;
    wire N__60433;
    wire N__60426;
    wire N__60423;
    wire N__60416;
    wire N__60413;
    wire N__60410;
    wire N__60407;
    wire N__60398;
    wire N__60397;
    wire N__60396;
    wire N__60395;
    wire N__60392;
    wire N__60389;
    wire N__60386;
    wire N__60381;
    wire N__60376;
    wire N__60371;
    wire N__60366;
    wire N__60359;
    wire N__60358;
    wire N__60357;
    wire N__60354;
    wire N__60353;
    wire N__60352;
    wire N__60349;
    wire N__60344;
    wire N__60341;
    wire N__60336;
    wire N__60331;
    wire N__60326;
    wire N__60321;
    wire N__60318;
    wire N__60315;
    wire N__60314;
    wire N__60313;
    wire N__60310;
    wire N__60309;
    wire N__60304;
    wire N__60301;
    wire N__60294;
    wire N__60285;
    wire N__60282;
    wire N__60273;
    wire N__60270;
    wire N__60269;
    wire N__60266;
    wire N__60263;
    wire N__60262;
    wire N__60251;
    wire N__60250;
    wire N__60249;
    wire N__60248;
    wire N__60247;
    wire N__60240;
    wire N__60237;
    wire N__60234;
    wire N__60233;
    wire N__60230;
    wire N__60225;
    wire N__60212;
    wire N__60209;
    wire N__60204;
    wire N__60195;
    wire N__60186;
    wire N__60181;
    wire N__60176;
    wire N__60173;
    wire N__60170;
    wire N__60167;
    wire N__60164;
    wire N__60157;
    wire N__60154;
    wire N__60151;
    wire N__60148;
    wire N__60143;
    wire N__60132;
    wire N__60123;
    wire N__60100;
    wire N__60099;
    wire N__60098;
    wire N__60097;
    wire N__60096;
    wire N__60095;
    wire N__60094;
    wire N__60093;
    wire N__60092;
    wire N__60091;
    wire N__60090;
    wire N__60087;
    wire N__60084;
    wire N__60083;
    wire N__60082;
    wire N__60081;
    wire N__60080;
    wire N__60077;
    wire N__60076;
    wire N__60073;
    wire N__60072;
    wire N__60069;
    wire N__60066;
    wire N__60065;
    wire N__60064;
    wire N__60063;
    wire N__60060;
    wire N__60059;
    wire N__60058;
    wire N__60053;
    wire N__60052;
    wire N__60049;
    wire N__60048;
    wire N__60047;
    wire N__60046;
    wire N__60045;
    wire N__60044;
    wire N__60043;
    wire N__60042;
    wire N__60041;
    wire N__60040;
    wire N__60037;
    wire N__60036;
    wire N__60031;
    wire N__60026;
    wire N__60021;
    wire N__60018;
    wire N__60015;
    wire N__60014;
    wire N__60009;
    wire N__60008;
    wire N__60007;
    wire N__60006;
    wire N__60003;
    wire N__60002;
    wire N__60001;
    wire N__60000;
    wire N__59999;
    wire N__59996;
    wire N__59995;
    wire N__59994;
    wire N__59993;
    wire N__59992;
    wire N__59991;
    wire N__59988;
    wire N__59987;
    wire N__59986;
    wire N__59985;
    wire N__59984;
    wire N__59983;
    wire N__59982;
    wire N__59979;
    wire N__59978;
    wire N__59977;
    wire N__59976;
    wire N__59975;
    wire N__59974;
    wire N__59973;
    wire N__59970;
    wire N__59969;
    wire N__59966;
    wire N__59965;
    wire N__59964;
    wire N__59963;
    wire N__59962;
    wire N__59961;
    wire N__59960;
    wire N__59955;
    wire N__59954;
    wire N__59951;
    wire N__59944;
    wire N__59937;
    wire N__59936;
    wire N__59933;
    wire N__59930;
    wire N__59925;
    wire N__59922;
    wire N__59917;
    wire N__59912;
    wire N__59905;
    wire N__59904;
    wire N__59901;
    wire N__59900;
    wire N__59897;
    wire N__59894;
    wire N__59891;
    wire N__59888;
    wire N__59887;
    wire N__59884;
    wire N__59881;
    wire N__59874;
    wire N__59871;
    wire N__59868;
    wire N__59867;
    wire N__59862;
    wire N__59857;
    wire N__59854;
    wire N__59851;
    wire N__59846;
    wire N__59839;
    wire N__59836;
    wire N__59831;
    wire N__59828;
    wire N__59823;
    wire N__59822;
    wire N__59819;
    wire N__59816;
    wire N__59813;
    wire N__59812;
    wire N__59809;
    wire N__59802;
    wire N__59797;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59785;
    wire N__59780;
    wire N__59777;
    wire N__59772;
    wire N__59769;
    wire N__59764;
    wire N__59759;
    wire N__59756;
    wire N__59751;
    wire N__59748;
    wire N__59743;
    wire N__59740;
    wire N__59737;
    wire N__59734;
    wire N__59725;
    wire N__59722;
    wire N__59717;
    wire N__59704;
    wire N__59703;
    wire N__59702;
    wire N__59697;
    wire N__59692;
    wire N__59687;
    wire N__59684;
    wire N__59673;
    wire N__59672;
    wire N__59661;
    wire N__59654;
    wire N__59649;
    wire N__59644;
    wire N__59629;
    wire N__59624;
    wire N__59619;
    wire N__59612;
    wire N__59609;
    wire N__59606;
    wire N__59601;
    wire N__59584;
    wire N__59581;
    wire N__59578;
    wire N__59575;
    wire N__59572;
    wire N__59569;
    wire N__59566;
    wire N__59563;
    wire N__59560;
    wire N__59557;
    wire N__59554;
    wire N__59551;
    wire N__59548;
    wire N__59545;
    wire N__59542;
    wire N__59539;
    wire N__59536;
    wire N__59533;
    wire N__59530;
    wire N__59527;
    wire N__59524;
    wire N__59521;
    wire N__59518;
    wire N__59517;
    wire N__59516;
    wire N__59515;
    wire N__59514;
    wire N__59513;
    wire N__59510;
    wire N__59509;
    wire N__59508;
    wire N__59507;
    wire N__59506;
    wire N__59505;
    wire N__59504;
    wire N__59503;
    wire N__59502;
    wire N__59501;
    wire N__59498;
    wire N__59497;
    wire N__59496;
    wire N__59493;
    wire N__59492;
    wire N__59491;
    wire N__59490;
    wire N__59489;
    wire N__59488;
    wire N__59485;
    wire N__59484;
    wire N__59483;
    wire N__59480;
    wire N__59479;
    wire N__59476;
    wire N__59475;
    wire N__59472;
    wire N__59469;
    wire N__59468;
    wire N__59467;
    wire N__59466;
    wire N__59461;
    wire N__59458;
    wire N__59455;
    wire N__59450;
    wire N__59447;
    wire N__59446;
    wire N__59445;
    wire N__59444;
    wire N__59443;
    wire N__59442;
    wire N__59441;
    wire N__59440;
    wire N__59439;
    wire N__59438;
    wire N__59437;
    wire N__59436;
    wire N__59435;
    wire N__59434;
    wire N__59433;
    wire N__59432;
    wire N__59431;
    wire N__59430;
    wire N__59429;
    wire N__59428;
    wire N__59427;
    wire N__59426;
    wire N__59425;
    wire N__59424;
    wire N__59423;
    wire N__59422;
    wire N__59421;
    wire N__59420;
    wire N__59417;
    wire N__59414;
    wire N__59411;
    wire N__59410;
    wire N__59409;
    wire N__59408;
    wire N__59407;
    wire N__59406;
    wire N__59405;
    wire N__59402;
    wire N__59401;
    wire N__59400;
    wire N__59399;
    wire N__59398;
    wire N__59397;
    wire N__59394;
    wire N__59391;
    wire N__59388;
    wire N__59381;
    wire N__59378;
    wire N__59373;
    wire N__59372;
    wire N__59371;
    wire N__59368;
    wire N__59367;
    wire N__59366;
    wire N__59365;
    wire N__59364;
    wire N__59363;
    wire N__59362;
    wire N__59359;
    wire N__59356;
    wire N__59355;
    wire N__59354;
    wire N__59353;
    wire N__59352;
    wire N__59351;
    wire N__59350;
    wire N__59347;
    wire N__59342;
    wire N__59337;
    wire N__59336;
    wire N__59335;
    wire N__59332;
    wire N__59331;
    wire N__59330;
    wire N__59329;
    wire N__59328;
    wire N__59327;
    wire N__59326;
    wire N__59325;
    wire N__59324;
    wire N__59323;
    wire N__59322;
    wire N__59321;
    wire N__59320;
    wire N__59317;
    wire N__59308;
    wire N__59307;
    wire N__59306;
    wire N__59305;
    wire N__59298;
    wire N__59293;
    wire N__59288;
    wire N__59283;
    wire N__59278;
    wire N__59269;
    wire N__59268;
    wire N__59267;
    wire N__59266;
    wire N__59265;
    wire N__59264;
    wire N__59263;
    wire N__59262;
    wire N__59261;
    wire N__59258;
    wire N__59251;
    wire N__59250;
    wire N__59247;
    wire N__59246;
    wire N__59241;
    wire N__59238;
    wire N__59231;
    wire N__59228;
    wire N__59227;
    wire N__59226;
    wire N__59225;
    wire N__59218;
    wire N__59215;
    wire N__59210;
    wire N__59209;
    wire N__59206;
    wire N__59201;
    wire N__59198;
    wire N__59193;
    wire N__59192;
    wire N__59191;
    wire N__59190;
    wire N__59189;
    wire N__59186;
    wire N__59185;
    wire N__59182;
    wire N__59181;
    wire N__59178;
    wire N__59165;
    wire N__59160;
    wire N__59157;
    wire N__59148;
    wire N__59143;
    wire N__59138;
    wire N__59127;
    wire N__59124;
    wire N__59121;
    wire N__59116;
    wire N__59115;
    wire N__59114;
    wire N__59113;
    wire N__59112;
    wire N__59111;
    wire N__59106;
    wire N__59103;
    wire N__59094;
    wire N__59091;
    wire N__59082;
    wire N__59079;
    wire N__59074;
    wire N__59069;
    wire N__59066;
    wire N__59063;
    wire N__59060;
    wire N__59057;
    wire N__59050;
    wire N__59045;
    wire N__59042;
    wire N__59035;
    wire N__59026;
    wire N__59021;
    wire N__59020;
    wire N__59017;
    wire N__59016;
    wire N__59015;
    wire N__59014;
    wire N__59011;
    wire N__59010;
    wire N__59009;
    wire N__59006;
    wire N__58999;
    wire N__58996;
    wire N__58993;
    wire N__58988;
    wire N__58981;
    wire N__58978;
    wire N__58973;
    wire N__58968;
    wire N__58963;
    wire N__58960;
    wire N__58957;
    wire N__58954;
    wire N__58951;
    wire N__58950;
    wire N__58949;
    wire N__58948;
    wire N__58945;
    wire N__58942;
    wire N__58939;
    wire N__58934;
    wire N__58923;
    wire N__58916;
    wire N__58915;
    wire N__58908;
    wire N__58905;
    wire N__58902;
    wire N__58899;
    wire N__58896;
    wire N__58889;
    wire N__58870;
    wire N__58861;
    wire N__58858;
    wire N__58857;
    wire N__58856;
    wire N__58855;
    wire N__58852;
    wire N__58845;
    wire N__58844;
    wire N__58843;
    wire N__58842;
    wire N__58841;
    wire N__58840;
    wire N__58837;
    wire N__58836;
    wire N__58831;
    wire N__58828;
    wire N__58823;
    wire N__58814;
    wire N__58807;
    wire N__58798;
    wire N__58791;
    wire N__58784;
    wire N__58777;
    wire N__58774;
    wire N__58771;
    wire N__58766;
    wire N__58753;
    wire N__58746;
    wire N__58743;
    wire N__58740;
    wire N__58733;
    wire N__58730;
    wire N__58727;
    wire N__58724;
    wire N__58721;
    wire N__58716;
    wire N__58709;
    wire N__58700;
    wire N__58689;
    wire N__58666;
    wire N__58663;
    wire N__58660;
    wire N__58657;
    wire N__58654;
    wire N__58653;
    wire N__58652;
    wire N__58651;
    wire N__58650;
    wire N__58649;
    wire N__58648;
    wire N__58643;
    wire N__58642;
    wire N__58641;
    wire N__58638;
    wire N__58635;
    wire N__58630;
    wire N__58627;
    wire N__58626;
    wire N__58625;
    wire N__58624;
    wire N__58621;
    wire N__58616;
    wire N__58615;
    wire N__58614;
    wire N__58611;
    wire N__58610;
    wire N__58609;
    wire N__58608;
    wire N__58607;
    wire N__58602;
    wire N__58599;
    wire N__58594;
    wire N__58591;
    wire N__58586;
    wire N__58585;
    wire N__58584;
    wire N__58581;
    wire N__58578;
    wire N__58575;
    wire N__58572;
    wire N__58567;
    wire N__58564;
    wire N__58557;
    wire N__58552;
    wire N__58547;
    wire N__58528;
    wire N__58527;
    wire N__58526;
    wire N__58523;
    wire N__58522;
    wire N__58521;
    wire N__58516;
    wire N__58515;
    wire N__58512;
    wire N__58511;
    wire N__58508;
    wire N__58505;
    wire N__58502;
    wire N__58499;
    wire N__58496;
    wire N__58493;
    wire N__58492;
    wire N__58491;
    wire N__58488;
    wire N__58487;
    wire N__58484;
    wire N__58483;
    wire N__58482;
    wire N__58475;
    wire N__58470;
    wire N__58469;
    wire N__58466;
    wire N__58463;
    wire N__58460;
    wire N__58457;
    wire N__58452;
    wire N__58447;
    wire N__58442;
    wire N__58429;
    wire N__58426;
    wire N__58423;
    wire N__58420;
    wire N__58417;
    wire N__58414;
    wire N__58411;
    wire N__58408;
    wire N__58407;
    wire N__58404;
    wire N__58403;
    wire N__58400;
    wire N__58399;
    wire N__58396;
    wire N__58393;
    wire N__58390;
    wire N__58387;
    wire N__58378;
    wire N__58375;
    wire N__58372;
    wire N__58369;
    wire N__58366;
    wire N__58365;
    wire N__58362;
    wire N__58359;
    wire N__58356;
    wire N__58353;
    wire N__58348;
    wire N__58345;
    wire N__58342;
    wire N__58339;
    wire N__58336;
    wire N__58333;
    wire N__58330;
    wire N__58327;
    wire N__58324;
    wire N__58321;
    wire N__58318;
    wire N__58315;
    wire N__58312;
    wire N__58309;
    wire N__58306;
    wire N__58303;
    wire N__58300;
    wire N__58297;
    wire N__58294;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58282;
    wire N__58279;
    wire N__58276;
    wire N__58273;
    wire N__58270;
    wire N__58267;
    wire N__58264;
    wire N__58261;
    wire N__58258;
    wire N__58255;
    wire N__58252;
    wire N__58249;
    wire N__58246;
    wire N__58243;
    wire N__58240;
    wire N__58237;
    wire N__58234;
    wire N__58231;
    wire N__58228;
    wire N__58225;
    wire N__58222;
    wire N__58219;
    wire N__58216;
    wire N__58213;
    wire N__58210;
    wire N__58209;
    wire N__58208;
    wire N__58207;
    wire N__58206;
    wire N__58205;
    wire N__58204;
    wire N__58201;
    wire N__58194;
    wire N__58193;
    wire N__58192;
    wire N__58189;
    wire N__58188;
    wire N__58187;
    wire N__58186;
    wire N__58185;
    wire N__58182;
    wire N__58181;
    wire N__58178;
    wire N__58173;
    wire N__58170;
    wire N__58161;
    wire N__58154;
    wire N__58153;
    wire N__58152;
    wire N__58151;
    wire N__58148;
    wire N__58147;
    wire N__58144;
    wire N__58141;
    wire N__58138;
    wire N__58133;
    wire N__58132;
    wire N__58129;
    wire N__58126;
    wire N__58119;
    wire N__58118;
    wire N__58117;
    wire N__58114;
    wire N__58107;
    wire N__58104;
    wire N__58097;
    wire N__58092;
    wire N__58089;
    wire N__58086;
    wire N__58083;
    wire N__58080;
    wire N__58077;
    wire N__58074;
    wire N__58071;
    wire N__58068;
    wire N__58063;
    wire N__58060;
    wire N__58055;
    wire N__58052;
    wire N__58047;
    wire N__58042;
    wire N__58041;
    wire N__58040;
    wire N__58039;
    wire N__58038;
    wire N__58037;
    wire N__58036;
    wire N__58035;
    wire N__58034;
    wire N__58033;
    wire N__58032;
    wire N__58031;
    wire N__58030;
    wire N__58023;
    wire N__58022;
    wire N__58019;
    wire N__58018;
    wire N__58011;
    wire N__58002;
    wire N__57999;
    wire N__57996;
    wire N__57993;
    wire N__57990;
    wire N__57985;
    wire N__57970;
    wire N__57967;
    wire N__57964;
    wire N__57961;
    wire N__57958;
    wire N__57957;
    wire N__57954;
    wire N__57953;
    wire N__57950;
    wire N__57947;
    wire N__57942;
    wire N__57937;
    wire N__57934;
    wire N__57931;
    wire N__57928;
    wire N__57925;
    wire N__57922;
    wire N__57919;
    wire N__57916;
    wire N__57913;
    wire N__57910;
    wire N__57907;
    wire N__57906;
    wire N__57905;
    wire N__57900;
    wire N__57897;
    wire N__57892;
    wire N__57889;
    wire N__57886;
    wire N__57883;
    wire N__57880;
    wire N__57879;
    wire N__57878;
    wire N__57877;
    wire N__57876;
    wire N__57873;
    wire N__57872;
    wire N__57871;
    wire N__57870;
    wire N__57869;
    wire N__57864;
    wire N__57863;
    wire N__57862;
    wire N__57861;
    wire N__57860;
    wire N__57857;
    wire N__57856;
    wire N__57855;
    wire N__57854;
    wire N__57853;
    wire N__57852;
    wire N__57851;
    wire N__57850;
    wire N__57849;
    wire N__57848;
    wire N__57845;
    wire N__57844;
    wire N__57841;
    wire N__57838;
    wire N__57835;
    wire N__57834;
    wire N__57833;
    wire N__57830;
    wire N__57827;
    wire N__57824;
    wire N__57821;
    wire N__57814;
    wire N__57811;
    wire N__57808;
    wire N__57805;
    wire N__57802;
    wire N__57799;
    wire N__57794;
    wire N__57789;
    wire N__57786;
    wire N__57783;
    wire N__57780;
    wire N__57779;
    wire N__57778;
    wire N__57775;
    wire N__57772;
    wire N__57765;
    wire N__57764;
    wire N__57763;
    wire N__57760;
    wire N__57757;
    wire N__57754;
    wire N__57751;
    wire N__57748;
    wire N__57747;
    wire N__57746;
    wire N__57745;
    wire N__57742;
    wire N__57741;
    wire N__57740;
    wire N__57739;
    wire N__57736;
    wire N__57731;
    wire N__57730;
    wire N__57729;
    wire N__57728;
    wire N__57723;
    wire N__57716;
    wire N__57713;
    wire N__57712;
    wire N__57711;
    wire N__57710;
    wire N__57709;
    wire N__57708;
    wire N__57707;
    wire N__57706;
    wire N__57705;
    wire N__57704;
    wire N__57703;
    wire N__57702;
    wire N__57701;
    wire N__57700;
    wire N__57697;
    wire N__57694;
    wire N__57693;
    wire N__57692;
    wire N__57687;
    wire N__57684;
    wire N__57681;
    wire N__57678;
    wire N__57673;
    wire N__57666;
    wire N__57665;
    wire N__57662;
    wire N__57661;
    wire N__57658;
    wire N__57655;
    wire N__57652;
    wire N__57647;
    wire N__57644;
    wire N__57639;
    wire N__57632;
    wire N__57625;
    wire N__57622;
    wire N__57621;
    wire N__57620;
    wire N__57619;
    wire N__57618;
    wire N__57617;
    wire N__57614;
    wire N__57611;
    wire N__57610;
    wire N__57607;
    wire N__57604;
    wire N__57603;
    wire N__57600;
    wire N__57591;
    wire N__57588;
    wire N__57587;
    wire N__57584;
    wire N__57583;
    wire N__57582;
    wire N__57571;
    wire N__57566;
    wire N__57563;
    wire N__57560;
    wire N__57557;
    wire N__57554;
    wire N__57551;
    wire N__57546;
    wire N__57543;
    wire N__57540;
    wire N__57535;
    wire N__57532;
    wire N__57527;
    wire N__57522;
    wire N__57521;
    wire N__57520;
    wire N__57517;
    wire N__57514;
    wire N__57509;
    wire N__57506;
    wire N__57501;
    wire N__57498;
    wire N__57489;
    wire N__57484;
    wire N__57475;
    wire N__57472;
    wire N__57469;
    wire N__57468;
    wire N__57465;
    wire N__57462;
    wire N__57455;
    wire N__57450;
    wire N__57445;
    wire N__57438;
    wire N__57435;
    wire N__57432;
    wire N__57429;
    wire N__57408;
    wire N__57405;
    wire N__57400;
    wire N__57397;
    wire N__57394;
    wire N__57389;
    wire N__57380;
    wire N__57367;
    wire N__57364;
    wire N__57361;
    wire N__57358;
    wire N__57355;
    wire N__57354;
    wire N__57353;
    wire N__57350;
    wire N__57347;
    wire N__57344;
    wire N__57337;
    wire N__57334;
    wire N__57331;
    wire N__57328;
    wire N__57325;
    wire N__57322;
    wire N__57319;
    wire N__57316;
    wire N__57313;
    wire N__57310;
    wire N__57307;
    wire N__57304;
    wire N__57301;
    wire N__57300;
    wire N__57299;
    wire N__57296;
    wire N__57293;
    wire N__57290;
    wire N__57283;
    wire N__57280;
    wire N__57277;
    wire N__57274;
    wire N__57271;
    wire N__57268;
    wire N__57265;
    wire N__57262;
    wire N__57261;
    wire N__57258;
    wire N__57255;
    wire N__57252;
    wire N__57249;
    wire N__57244;
    wire N__57243;
    wire N__57240;
    wire N__57237;
    wire N__57232;
    wire N__57231;
    wire N__57228;
    wire N__57225;
    wire N__57222;
    wire N__57217;
    wire N__57216;
    wire N__57213;
    wire N__57210;
    wire N__57205;
    wire N__57202;
    wire N__57199;
    wire N__57196;
    wire N__57195;
    wire N__57192;
    wire N__57189;
    wire N__57186;
    wire N__57183;
    wire N__57178;
    wire N__57177;
    wire N__57176;
    wire N__57175;
    wire N__57174;
    wire N__57173;
    wire N__57172;
    wire N__57171;
    wire N__57170;
    wire N__57167;
    wire N__57164;
    wire N__57161;
    wire N__57148;
    wire N__57147;
    wire N__57138;
    wire N__57137;
    wire N__57136;
    wire N__57135;
    wire N__57132;
    wire N__57131;
    wire N__57130;
    wire N__57129;
    wire N__57126;
    wire N__57123;
    wire N__57122;
    wire N__57121;
    wire N__57120;
    wire N__57119;
    wire N__57118;
    wire N__57117;
    wire N__57116;
    wire N__57115;
    wire N__57114;
    wire N__57113;
    wire N__57112;
    wire N__57111;
    wire N__57110;
    wire N__57109;
    wire N__57100;
    wire N__57097;
    wire N__57096;
    wire N__57093;
    wire N__57092;
    wire N__57087;
    wire N__57084;
    wire N__57079;
    wire N__57078;
    wire N__57077;
    wire N__57074;
    wire N__57071;
    wire N__57070;
    wire N__57063;
    wire N__57058;
    wire N__57053;
    wire N__57050;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57040;
    wire N__57037;
    wire N__57034;
    wire N__57031;
    wire N__57028;
    wire N__57025;
    wire N__57022;
    wire N__57019;
    wire N__57016;
    wire N__57011;
    wire N__57008;
    wire N__57003;
    wire N__57000;
    wire N__56997;
    wire N__56994;
    wire N__56989;
    wire N__56984;
    wire N__56979;
    wire N__56972;
    wire N__56969;
    wire N__56962;
    wire N__56957;
    wire N__56950;
    wire N__56947;
    wire N__56938;
    wire N__56933;
    wire N__56926;
    wire N__56923;
    wire N__56920;
    wire N__56917;
    wire N__56914;
    wire N__56911;
    wire N__56908;
    wire N__56905;
    wire N__56902;
    wire N__56899;
    wire N__56896;
    wire N__56893;
    wire N__56890;
    wire N__56887;
    wire N__56884;
    wire N__56881;
    wire N__56878;
    wire N__56875;
    wire N__56872;
    wire N__56871;
    wire N__56868;
    wire N__56865;
    wire N__56862;
    wire N__56859;
    wire N__56854;
    wire N__56851;
    wire N__56850;
    wire N__56849;
    wire N__56846;
    wire N__56843;
    wire N__56840;
    wire N__56839;
    wire N__56838;
    wire N__56835;
    wire N__56834;
    wire N__56831;
    wire N__56828;
    wire N__56825;
    wire N__56822;
    wire N__56819;
    wire N__56816;
    wire N__56813;
    wire N__56810;
    wire N__56807;
    wire N__56804;
    wire N__56799;
    wire N__56796;
    wire N__56793;
    wire N__56790;
    wire N__56785;
    wire N__56776;
    wire N__56773;
    wire N__56770;
    wire N__56767;
    wire N__56764;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56752;
    wire N__56751;
    wire N__56748;
    wire N__56745;
    wire N__56740;
    wire N__56739;
    wire N__56736;
    wire N__56733;
    wire N__56730;
    wire N__56727;
    wire N__56722;
    wire N__56721;
    wire N__56718;
    wire N__56715;
    wire N__56710;
    wire N__56707;
    wire N__56706;
    wire N__56703;
    wire N__56700;
    wire N__56697;
    wire N__56692;
    wire N__56689;
    wire N__56688;
    wire N__56685;
    wire N__56682;
    wire N__56677;
    wire N__56676;
    wire N__56673;
    wire N__56670;
    wire N__56667;
    wire N__56662;
    wire N__56661;
    wire N__56658;
    wire N__56655;
    wire N__56650;
    wire N__56647;
    wire N__56644;
    wire N__56643;
    wire N__56640;
    wire N__56637;
    wire N__56632;
    wire N__56629;
    wire N__56628;
    wire N__56625;
    wire N__56622;
    wire N__56617;
    wire N__56616;
    wire N__56613;
    wire N__56610;
    wire N__56607;
    wire N__56602;
    wire N__56599;
    wire N__56598;
    wire N__56595;
    wire N__56592;
    wire N__56587;
    wire N__56584;
    wire N__56583;
    wire N__56582;
    wire N__56579;
    wire N__56578;
    wire N__56577;
    wire N__56574;
    wire N__56571;
    wire N__56570;
    wire N__56569;
    wire N__56566;
    wire N__56563;
    wire N__56560;
    wire N__56557;
    wire N__56554;
    wire N__56551;
    wire N__56548;
    wire N__56543;
    wire N__56540;
    wire N__56533;
    wire N__56532;
    wire N__56529;
    wire N__56526;
    wire N__56521;
    wire N__56518;
    wire N__56515;
    wire N__56508;
    wire N__56503;
    wire N__56502;
    wire N__56499;
    wire N__56496;
    wire N__56495;
    wire N__56490;
    wire N__56487;
    wire N__56484;
    wire N__56479;
    wire N__56478;
    wire N__56475;
    wire N__56474;
    wire N__56473;
    wire N__56470;
    wire N__56469;
    wire N__56466;
    wire N__56463;
    wire N__56462;
    wire N__56461;
    wire N__56460;
    wire N__56459;
    wire N__56458;
    wire N__56455;
    wire N__56452;
    wire N__56451;
    wire N__56448;
    wire N__56445;
    wire N__56442;
    wire N__56439;
    wire N__56434;
    wire N__56429;
    wire N__56426;
    wire N__56423;
    wire N__56420;
    wire N__56417;
    wire N__56414;
    wire N__56405;
    wire N__56396;
    wire N__56389;
    wire N__56386;
    wire N__56383;
    wire N__56380;
    wire N__56377;
    wire N__56376;
    wire N__56373;
    wire N__56370;
    wire N__56365;
    wire N__56362;
    wire N__56359;
    wire N__56356;
    wire N__56353;
    wire N__56350;
    wire N__56347;
    wire N__56344;
    wire N__56341;
    wire N__56338;
    wire N__56335;
    wire N__56332;
    wire N__56329;
    wire N__56328;
    wire N__56325;
    wire N__56322;
    wire N__56319;
    wire N__56316;
    wire N__56313;
    wire N__56310;
    wire N__56307;
    wire N__56304;
    wire N__56301;
    wire N__56298;
    wire N__56295;
    wire N__56292;
    wire N__56289;
    wire N__56286;
    wire N__56283;
    wire N__56280;
    wire N__56277;
    wire N__56274;
    wire N__56271;
    wire N__56268;
    wire N__56265;
    wire N__56260;
    wire N__56257;
    wire N__56254;
    wire N__56251;
    wire N__56248;
    wire N__56247;
    wire N__56244;
    wire N__56241;
    wire N__56236;
    wire N__56233;
    wire N__56232;
    wire N__56229;
    wire N__56228;
    wire N__56225;
    wire N__56222;
    wire N__56217;
    wire N__56212;
    wire N__56209;
    wire N__56206;
    wire N__56205;
    wire N__56202;
    wire N__56199;
    wire N__56196;
    wire N__56193;
    wire N__56190;
    wire N__56185;
    wire N__56184;
    wire N__56181;
    wire N__56178;
    wire N__56173;
    wire N__56170;
    wire N__56167;
    wire N__56164;
    wire N__56161;
    wire N__56158;
    wire N__56157;
    wire N__56154;
    wire N__56151;
    wire N__56148;
    wire N__56145;
    wire N__56142;
    wire N__56137;
    wire N__56134;
    wire N__56133;
    wire N__56132;
    wire N__56129;
    wire N__56126;
    wire N__56123;
    wire N__56120;
    wire N__56117;
    wire N__56110;
    wire N__56109;
    wire N__56106;
    wire N__56103;
    wire N__56100;
    wire N__56097;
    wire N__56096;
    wire N__56093;
    wire N__56090;
    wire N__56087;
    wire N__56086;
    wire N__56079;
    wire N__56078;
    wire N__56075;
    wire N__56074;
    wire N__56071;
    wire N__56070;
    wire N__56069;
    wire N__56066;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56056;
    wire N__56051;
    wire N__56048;
    wire N__56045;
    wire N__56042;
    wire N__56037;
    wire N__56030;
    wire N__56023;
    wire N__56022;
    wire N__56019;
    wire N__56016;
    wire N__56013;
    wire N__56010;
    wire N__56007;
    wire N__56004;
    wire N__55999;
    wire N__55996;
    wire N__55993;
    wire N__55990;
    wire N__55987;
    wire N__55984;
    wire N__55981;
    wire N__55978;
    wire N__55975;
    wire N__55972;
    wire N__55969;
    wire N__55966;
    wire N__55963;
    wire N__55960;
    wire N__55957;
    wire N__55954;
    wire N__55951;
    wire N__55948;
    wire N__55945;
    wire N__55942;
    wire N__55941;
    wire N__55938;
    wire N__55937;
    wire N__55936;
    wire N__55935;
    wire N__55932;
    wire N__55931;
    wire N__55928;
    wire N__55925;
    wire N__55922;
    wire N__55917;
    wire N__55914;
    wire N__55909;
    wire N__55906;
    wire N__55903;
    wire N__55900;
    wire N__55899;
    wire N__55896;
    wire N__55893;
    wire N__55888;
    wire N__55885;
    wire N__55884;
    wire N__55881;
    wire N__55878;
    wire N__55873;
    wire N__55870;
    wire N__55867;
    wire N__55862;
    wire N__55859;
    wire N__55852;
    wire N__55849;
    wire N__55848;
    wire N__55845;
    wire N__55842;
    wire N__55841;
    wire N__55838;
    wire N__55837;
    wire N__55834;
    wire N__55831;
    wire N__55828;
    wire N__55827;
    wire N__55824;
    wire N__55823;
    wire N__55822;
    wire N__55817;
    wire N__55814;
    wire N__55811;
    wire N__55808;
    wire N__55805;
    wire N__55802;
    wire N__55799;
    wire N__55792;
    wire N__55787;
    wire N__55784;
    wire N__55781;
    wire N__55774;
    wire N__55771;
    wire N__55770;
    wire N__55769;
    wire N__55768;
    wire N__55767;
    wire N__55764;
    wire N__55761;
    wire N__55758;
    wire N__55755;
    wire N__55752;
    wire N__55751;
    wire N__55746;
    wire N__55743;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55729;
    wire N__55724;
    wire N__55721;
    wire N__55714;
    wire N__55711;
    wire N__55710;
    wire N__55709;
    wire N__55708;
    wire N__55707;
    wire N__55704;
    wire N__55701;
    wire N__55700;
    wire N__55697;
    wire N__55694;
    wire N__55691;
    wire N__55686;
    wire N__55683;
    wire N__55678;
    wire N__55675;
    wire N__55670;
    wire N__55667;
    wire N__55664;
    wire N__55661;
    wire N__55658;
    wire N__55651;
    wire N__55650;
    wire N__55649;
    wire N__55646;
    wire N__55641;
    wire N__55640;
    wire N__55637;
    wire N__55636;
    wire N__55635;
    wire N__55634;
    wire N__55631;
    wire N__55630;
    wire N__55627;
    wire N__55626;
    wire N__55623;
    wire N__55616;
    wire N__55613;
    wire N__55610;
    wire N__55607;
    wire N__55604;
    wire N__55599;
    wire N__55598;
    wire N__55595;
    wire N__55592;
    wire N__55589;
    wire N__55584;
    wire N__55581;
    wire N__55576;
    wire N__55573;
    wire N__55570;
    wire N__55565;
    wire N__55558;
    wire N__55555;
    wire N__55552;
    wire N__55549;
    wire N__55548;
    wire N__55545;
    wire N__55542;
    wire N__55539;
    wire N__55536;
    wire N__55533;
    wire N__55530;
    wire N__55529;
    wire N__55526;
    wire N__55523;
    wire N__55520;
    wire N__55515;
    wire N__55510;
    wire N__55507;
    wire N__55504;
    wire N__55501;
    wire N__55498;
    wire N__55497;
    wire N__55494;
    wire N__55491;
    wire N__55490;
    wire N__55487;
    wire N__55482;
    wire N__55477;
    wire N__55474;
    wire N__55471;
    wire N__55470;
    wire N__55469;
    wire N__55466;
    wire N__55461;
    wire N__55456;
    wire N__55453;
    wire N__55450;
    wire N__55447;
    wire N__55444;
    wire N__55441;
    wire N__55438;
    wire N__55435;
    wire N__55432;
    wire N__55431;
    wire N__55430;
    wire N__55427;
    wire N__55424;
    wire N__55423;
    wire N__55420;
    wire N__55415;
    wire N__55412;
    wire N__55409;
    wire N__55404;
    wire N__55403;
    wire N__55402;
    wire N__55401;
    wire N__55400;
    wire N__55399;
    wire N__55394;
    wire N__55389;
    wire N__55388;
    wire N__55385;
    wire N__55382;
    wire N__55381;
    wire N__55380;
    wire N__55377;
    wire N__55372;
    wire N__55371;
    wire N__55370;
    wire N__55369;
    wire N__55368;
    wire N__55365;
    wire N__55362;
    wire N__55359;
    wire N__55356;
    wire N__55353;
    wire N__55348;
    wire N__55345;
    wire N__55338;
    wire N__55335;
    wire N__55332;
    wire N__55329;
    wire N__55326;
    wire N__55323;
    wire N__55320;
    wire N__55313;
    wire N__55310;
    wire N__55307;
    wire N__55304;
    wire N__55297;
    wire N__55288;
    wire N__55287;
    wire N__55284;
    wire N__55283;
    wire N__55280;
    wire N__55277;
    wire N__55276;
    wire N__55273;
    wire N__55270;
    wire N__55267;
    wire N__55264;
    wire N__55261;
    wire N__55258;
    wire N__55255;
    wire N__55252;
    wire N__55249;
    wire N__55246;
    wire N__55237;
    wire N__55234;
    wire N__55231;
    wire N__55228;
    wire N__55227;
    wire N__55224;
    wire N__55223;
    wire N__55220;
    wire N__55217;
    wire N__55214;
    wire N__55207;
    wire N__55206;
    wire N__55203;
    wire N__55200;
    wire N__55195;
    wire N__55194;
    wire N__55193;
    wire N__55190;
    wire N__55189;
    wire N__55186;
    wire N__55183;
    wire N__55180;
    wire N__55177;
    wire N__55174;
    wire N__55171;
    wire N__55170;
    wire N__55169;
    wire N__55164;
    wire N__55161;
    wire N__55160;
    wire N__55157;
    wire N__55154;
    wire N__55151;
    wire N__55148;
    wire N__55145;
    wire N__55142;
    wire N__55139;
    wire N__55136;
    wire N__55133;
    wire N__55132;
    wire N__55129;
    wire N__55124;
    wire N__55117;
    wire N__55114;
    wire N__55105;
    wire N__55102;
    wire N__55099;
    wire N__55096;
    wire N__55093;
    wire N__55090;
    wire N__55087;
    wire N__55084;
    wire N__55081;
    wire N__55078;
    wire N__55077;
    wire N__55076;
    wire N__55073;
    wire N__55072;
    wire N__55071;
    wire N__55068;
    wire N__55067;
    wire N__55064;
    wire N__55061;
    wire N__55060;
    wire N__55057;
    wire N__55054;
    wire N__55051;
    wire N__55048;
    wire N__55045;
    wire N__55042;
    wire N__55039;
    wire N__55038;
    wire N__55033;
    wire N__55028;
    wire N__55025;
    wire N__55020;
    wire N__55017;
    wire N__55016;
    wire N__55013;
    wire N__55010;
    wire N__55003;
    wire N__55000;
    wire N__54991;
    wire N__54988;
    wire N__54985;
    wire N__54982;
    wire N__54979;
    wire N__54976;
    wire N__54973;
    wire N__54970;
    wire N__54967;
    wire N__54964;
    wire N__54961;
    wire N__54958;
    wire N__54955;
    wire N__54952;
    wire N__54949;
    wire N__54946;
    wire N__54943;
    wire N__54940;
    wire N__54939;
    wire N__54938;
    wire N__54935;
    wire N__54932;
    wire N__54931;
    wire N__54930;
    wire N__54929;
    wire N__54926;
    wire N__54925;
    wire N__54920;
    wire N__54917;
    wire N__54914;
    wire N__54911;
    wire N__54908;
    wire N__54905;
    wire N__54900;
    wire N__54897;
    wire N__54896;
    wire N__54893;
    wire N__54888;
    wire N__54885;
    wire N__54882;
    wire N__54879;
    wire N__54878;
    wire N__54875;
    wire N__54872;
    wire N__54869;
    wire N__54864;
    wire N__54861;
    wire N__54850;
    wire N__54847;
    wire N__54844;
    wire N__54841;
    wire N__54838;
    wire N__54835;
    wire N__54832;
    wire N__54829;
    wire N__54826;
    wire N__54823;
    wire N__54820;
    wire N__54817;
    wire N__54816;
    wire N__54813;
    wire N__54810;
    wire N__54809;
    wire N__54804;
    wire N__54801;
    wire N__54800;
    wire N__54797;
    wire N__54796;
    wire N__54793;
    wire N__54792;
    wire N__54789;
    wire N__54788;
    wire N__54785;
    wire N__54782;
    wire N__54779;
    wire N__54776;
    wire N__54773;
    wire N__54770;
    wire N__54769;
    wire N__54764;
    wire N__54759;
    wire N__54754;
    wire N__54751;
    wire N__54750;
    wire N__54747;
    wire N__54744;
    wire N__54741;
    wire N__54738;
    wire N__54735;
    wire N__54724;
    wire N__54721;
    wire N__54718;
    wire N__54715;
    wire N__54712;
    wire N__54709;
    wire N__54706;
    wire N__54703;
    wire N__54700;
    wire N__54697;
    wire N__54694;
    wire N__54691;
    wire N__54688;
    wire N__54685;
    wire N__54682;
    wire N__54679;
    wire N__54676;
    wire N__54673;
    wire N__54672;
    wire N__54669;
    wire N__54666;
    wire N__54663;
    wire N__54658;
    wire N__54657;
    wire N__54654;
    wire N__54651;
    wire N__54650;
    wire N__54647;
    wire N__54644;
    wire N__54641;
    wire N__54638;
    wire N__54635;
    wire N__54628;
    wire N__54625;
    wire N__54622;
    wire N__54619;
    wire N__54616;
    wire N__54613;
    wire N__54612;
    wire N__54611;
    wire N__54610;
    wire N__54609;
    wire N__54608;
    wire N__54603;
    wire N__54602;
    wire N__54601;
    wire N__54600;
    wire N__54599;
    wire N__54596;
    wire N__54593;
    wire N__54590;
    wire N__54589;
    wire N__54588;
    wire N__54587;
    wire N__54586;
    wire N__54585;
    wire N__54584;
    wire N__54581;
    wire N__54578;
    wire N__54573;
    wire N__54572;
    wire N__54567;
    wire N__54562;
    wire N__54559;
    wire N__54550;
    wire N__54547;
    wire N__54546;
    wire N__54543;
    wire N__54542;
    wire N__54541;
    wire N__54540;
    wire N__54539;
    wire N__54538;
    wire N__54537;
    wire N__54534;
    wire N__54529;
    wire N__54528;
    wire N__54527;
    wire N__54526;
    wire N__54525;
    wire N__54522;
    wire N__54513;
    wire N__54510;
    wire N__54507;
    wire N__54504;
    wire N__54495;
    wire N__54490;
    wire N__54487;
    wire N__54484;
    wire N__54475;
    wire N__54468;
    wire N__54465;
    wire N__54458;
    wire N__54445;
    wire N__54444;
    wire N__54441;
    wire N__54438;
    wire N__54435;
    wire N__54430;
    wire N__54427;
    wire N__54424;
    wire N__54423;
    wire N__54422;
    wire N__54421;
    wire N__54420;
    wire N__54419;
    wire N__54418;
    wire N__54417;
    wire N__54416;
    wire N__54415;
    wire N__54414;
    wire N__54413;
    wire N__54410;
    wire N__54409;
    wire N__54408;
    wire N__54407;
    wire N__54406;
    wire N__54405;
    wire N__54402;
    wire N__54401;
    wire N__54400;
    wire N__54399;
    wire N__54398;
    wire N__54391;
    wire N__54388;
    wire N__54385;
    wire N__54382;
    wire N__54373;
    wire N__54372;
    wire N__54371;
    wire N__54370;
    wire N__54367;
    wire N__54364;
    wire N__54363;
    wire N__54362;
    wire N__54353;
    wire N__54350;
    wire N__54341;
    wire N__54338;
    wire N__54335;
    wire N__54332;
    wire N__54331;
    wire N__54330;
    wire N__54327;
    wire N__54326;
    wire N__54323;
    wire N__54316;
    wire N__54313;
    wire N__54312;
    wire N__54311;
    wire N__54310;
    wire N__54309;
    wire N__54308;
    wire N__54307;
    wire N__54306;
    wire N__54303;
    wire N__54298;
    wire N__54293;
    wire N__54290;
    wire N__54287;
    wire N__54282;
    wire N__54277;
    wire N__54274;
    wire N__54271;
    wire N__54264;
    wire N__54259;
    wire N__54254;
    wire N__54251;
    wire N__54246;
    wire N__54243;
    wire N__54234;
    wire N__54231;
    wire N__54220;
    wire N__54205;
    wire N__54202;
    wire N__54199;
    wire N__54198;
    wire N__54195;
    wire N__54192;
    wire N__54189;
    wire N__54184;
    wire N__54183;
    wire N__54182;
    wire N__54179;
    wire N__54176;
    wire N__54175;
    wire N__54172;
    wire N__54171;
    wire N__54168;
    wire N__54165;
    wire N__54162;
    wire N__54161;
    wire N__54160;
    wire N__54159;
    wire N__54156;
    wire N__54153;
    wire N__54150;
    wire N__54145;
    wire N__54142;
    wire N__54137;
    wire N__54136;
    wire N__54131;
    wire N__54128;
    wire N__54125;
    wire N__54122;
    wire N__54119;
    wire N__54116;
    wire N__54113;
    wire N__54110;
    wire N__54101;
    wire N__54098;
    wire N__54091;
    wire N__54088;
    wire N__54085;
    wire N__54082;
    wire N__54081;
    wire N__54078;
    wire N__54075;
    wire N__54072;
    wire N__54069;
    wire N__54068;
    wire N__54067;
    wire N__54066;
    wire N__54065;
    wire N__54060;
    wire N__54057;
    wire N__54052;
    wire N__54049;
    wire N__54044;
    wire N__54037;
    wire N__54034;
    wire N__54031;
    wire N__54028;
    wire N__54025;
    wire N__54024;
    wire N__54023;
    wire N__54022;
    wire N__54021;
    wire N__54020;
    wire N__54017;
    wire N__54016;
    wire N__54015;
    wire N__54012;
    wire N__54009;
    wire N__54006;
    wire N__54003;
    wire N__54000;
    wire N__53997;
    wire N__53994;
    wire N__53991;
    wire N__53990;
    wire N__53987;
    wire N__53984;
    wire N__53979;
    wire N__53970;
    wire N__53967;
    wire N__53964;
    wire N__53961;
    wire N__53958;
    wire N__53953;
    wire N__53948;
    wire N__53943;
    wire N__53938;
    wire N__53935;
    wire N__53932;
    wire N__53929;
    wire N__53926;
    wire N__53923;
    wire N__53920;
    wire N__53917;
    wire N__53914;
    wire N__53911;
    wire N__53908;
    wire N__53905;
    wire N__53902;
    wire N__53899;
    wire N__53896;
    wire N__53895;
    wire N__53894;
    wire N__53893;
    wire N__53890;
    wire N__53887;
    wire N__53884;
    wire N__53883;
    wire N__53880;
    wire N__53879;
    wire N__53874;
    wire N__53871;
    wire N__53868;
    wire N__53865;
    wire N__53862;
    wire N__53857;
    wire N__53856;
    wire N__53855;
    wire N__53852;
    wire N__53847;
    wire N__53844;
    wire N__53841;
    wire N__53838;
    wire N__53837;
    wire N__53834;
    wire N__53827;
    wire N__53824;
    wire N__53821;
    wire N__53812;
    wire N__53809;
    wire N__53806;
    wire N__53803;
    wire N__53800;
    wire N__53797;
    wire N__53794;
    wire N__53791;
    wire N__53788;
    wire N__53785;
    wire N__53782;
    wire N__53781;
    wire N__53780;
    wire N__53779;
    wire N__53778;
    wire N__53777;
    wire N__53776;
    wire N__53775;
    wire N__53772;
    wire N__53771;
    wire N__53756;
    wire N__53753;
    wire N__53750;
    wire N__53747;
    wire N__53740;
    wire N__53739;
    wire N__53738;
    wire N__53737;
    wire N__53736;
    wire N__53735;
    wire N__53734;
    wire N__53733;
    wire N__53730;
    wire N__53715;
    wire N__53710;
    wire N__53707;
    wire N__53706;
    wire N__53703;
    wire N__53700;
    wire N__53699;
    wire N__53698;
    wire N__53697;
    wire N__53692;
    wire N__53691;
    wire N__53690;
    wire N__53689;
    wire N__53688;
    wire N__53685;
    wire N__53682;
    wire N__53679;
    wire N__53678;
    wire N__53677;
    wire N__53674;
    wire N__53671;
    wire N__53670;
    wire N__53667;
    wire N__53666;
    wire N__53665;
    wire N__53662;
    wire N__53659;
    wire N__53656;
    wire N__53653;
    wire N__53650;
    wire N__53647;
    wire N__53644;
    wire N__53639;
    wire N__53638;
    wire N__53635;
    wire N__53634;
    wire N__53631;
    wire N__53628;
    wire N__53627;
    wire N__53624;
    wire N__53621;
    wire N__53618;
    wire N__53617;
    wire N__53614;
    wire N__53609;
    wire N__53606;
    wire N__53603;
    wire N__53602;
    wire N__53601;
    wire N__53598;
    wire N__53595;
    wire N__53592;
    wire N__53589;
    wire N__53588;
    wire N__53583;
    wire N__53580;
    wire N__53577;
    wire N__53572;
    wire N__53569;
    wire N__53568;
    wire N__53561;
    wire N__53558;
    wire N__53555;
    wire N__53552;
    wire N__53547;
    wire N__53542;
    wire N__53539;
    wire N__53534;
    wire N__53531;
    wire N__53526;
    wire N__53523;
    wire N__53520;
    wire N__53517;
    wire N__53514;
    wire N__53511;
    wire N__53504;
    wire N__53501;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53485;
    wire N__53480;
    wire N__53473;
    wire N__53464;
    wire N__53461;
    wire N__53458;
    wire N__53455;
    wire N__53452;
    wire N__53449;
    wire N__53446;
    wire N__53443;
    wire N__53440;
    wire N__53439;
    wire N__53438;
    wire N__53435;
    wire N__53432;
    wire N__53429;
    wire N__53426;
    wire N__53419;
    wire N__53416;
    wire N__53413;
    wire N__53410;
    wire N__53409;
    wire N__53406;
    wire N__53403;
    wire N__53398;
    wire N__53395;
    wire N__53392;
    wire N__53391;
    wire N__53388;
    wire N__53385;
    wire N__53380;
    wire N__53377;
    wire N__53374;
    wire N__53371;
    wire N__53368;
    wire N__53365;
    wire N__53364;
    wire N__53361;
    wire N__53358;
    wire N__53353;
    wire N__53350;
    wire N__53349;
    wire N__53346;
    wire N__53343;
    wire N__53338;
    wire N__53335;
    wire N__53332;
    wire N__53329;
    wire N__53326;
    wire N__53323;
    wire N__53320;
    wire N__53317;
    wire N__53314;
    wire N__53313;
    wire N__53310;
    wire N__53307;
    wire N__53302;
    wire N__53301;
    wire N__53298;
    wire N__53295;
    wire N__53290;
    wire N__53287;
    wire N__53286;
    wire N__53283;
    wire N__53280;
    wire N__53277;
    wire N__53272;
    wire N__53271;
    wire N__53268;
    wire N__53265;
    wire N__53260;
    wire N__53259;
    wire N__53256;
    wire N__53253;
    wire N__53250;
    wire N__53245;
    wire N__53244;
    wire N__53241;
    wire N__53238;
    wire N__53233;
    wire N__53230;
    wire N__53229;
    wire N__53226;
    wire N__53223;
    wire N__53218;
    wire N__53217;
    wire N__53212;
    wire N__53209;
    wire N__53206;
    wire N__53203;
    wire N__53200;
    wire N__53197;
    wire N__53194;
    wire N__53191;
    wire N__53188;
    wire N__53185;
    wire N__53182;
    wire N__53179;
    wire N__53176;
    wire N__53173;
    wire N__53170;
    wire N__53167;
    wire N__53164;
    wire N__53161;
    wire N__53158;
    wire N__53155;
    wire N__53152;
    wire N__53151;
    wire N__53148;
    wire N__53145;
    wire N__53142;
    wire N__53139;
    wire N__53136;
    wire N__53133;
    wire N__53130;
    wire N__53127;
    wire N__53122;
    wire N__53119;
    wire N__53116;
    wire N__53113;
    wire N__53110;
    wire N__53107;
    wire N__53104;
    wire N__53101;
    wire N__53098;
    wire N__53095;
    wire N__53092;
    wire N__53089;
    wire N__53086;
    wire N__53083;
    wire N__53082;
    wire N__53079;
    wire N__53076;
    wire N__53073;
    wire N__53070;
    wire N__53067;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53052;
    wire N__53049;
    wire N__53046;
    wire N__53043;
    wire N__53038;
    wire N__53035;
    wire N__53032;
    wire N__53029;
    wire N__53026;
    wire N__53023;
    wire N__53020;
    wire N__53017;
    wire N__53014;
    wire N__53011;
    wire N__53008;
    wire N__53005;
    wire N__53002;
    wire N__52999;
    wire N__52996;
    wire N__52993;
    wire N__52990;
    wire N__52987;
    wire N__52984;
    wire N__52981;
    wire N__52978;
    wire N__52975;
    wire N__52972;
    wire N__52969;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52957;
    wire N__52954;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52939;
    wire N__52936;
    wire N__52935;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52927;
    wire N__52926;
    wire N__52925;
    wire N__52922;
    wire N__52919;
    wire N__52916;
    wire N__52913;
    wire N__52910;
    wire N__52909;
    wire N__52906;
    wire N__52901;
    wire N__52896;
    wire N__52893;
    wire N__52890;
    wire N__52889;
    wire N__52888;
    wire N__52885;
    wire N__52880;
    wire N__52875;
    wire N__52870;
    wire N__52867;
    wire N__52864;
    wire N__52859;
    wire N__52856;
    wire N__52853;
    wire N__52850;
    wire N__52843;
    wire N__52842;
    wire N__52839;
    wire N__52836;
    wire N__52833;
    wire N__52832;
    wire N__52829;
    wire N__52826;
    wire N__52823;
    wire N__52816;
    wire N__52813;
    wire N__52812;
    wire N__52811;
    wire N__52808;
    wire N__52805;
    wire N__52802;
    wire N__52799;
    wire N__52796;
    wire N__52793;
    wire N__52786;
    wire N__52783;
    wire N__52780;
    wire N__52779;
    wire N__52776;
    wire N__52773;
    wire N__52770;
    wire N__52767;
    wire N__52764;
    wire N__52763;
    wire N__52760;
    wire N__52757;
    wire N__52754;
    wire N__52751;
    wire N__52744;
    wire N__52743;
    wire N__52742;
    wire N__52739;
    wire N__52736;
    wire N__52733;
    wire N__52730;
    wire N__52727;
    wire N__52720;
    wire N__52717;
    wire N__52716;
    wire N__52713;
    wire N__52710;
    wire N__52705;
    wire N__52704;
    wire N__52701;
    wire N__52698;
    wire N__52695;
    wire N__52690;
    wire N__52687;
    wire N__52684;
    wire N__52681;
    wire N__52678;
    wire N__52675;
    wire N__52672;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52660;
    wire N__52659;
    wire N__52658;
    wire N__52655;
    wire N__52652;
    wire N__52649;
    wire N__52642;
    wire N__52639;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52626;
    wire N__52625;
    wire N__52622;
    wire N__52619;
    wire N__52616;
    wire N__52613;
    wire N__52606;
    wire N__52603;
    wire N__52600;
    wire N__52597;
    wire N__52594;
    wire N__52591;
    wire N__52588;
    wire N__52587;
    wire N__52584;
    wire N__52581;
    wire N__52578;
    wire N__52575;
    wire N__52572;
    wire N__52567;
    wire N__52564;
    wire N__52563;
    wire N__52560;
    wire N__52557;
    wire N__52554;
    wire N__52549;
    wire N__52546;
    wire N__52545;
    wire N__52542;
    wire N__52541;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52525;
    wire N__52522;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52512;
    wire N__52509;
    wire N__52506;
    wire N__52505;
    wire N__52502;
    wire N__52499;
    wire N__52496;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52482;
    wire N__52481;
    wire N__52478;
    wire N__52475;
    wire N__52472;
    wire N__52467;
    wire N__52462;
    wire N__52459;
    wire N__52456;
    wire N__52453;
    wire N__52450;
    wire N__52447;
    wire N__52444;
    wire N__52441;
    wire N__52438;
    wire N__52435;
    wire N__52432;
    wire N__52429;
    wire N__52426;
    wire N__52423;
    wire N__52420;
    wire N__52419;
    wire N__52416;
    wire N__52413;
    wire N__52408;
    wire N__52405;
    wire N__52402;
    wire N__52399;
    wire N__52398;
    wire N__52397;
    wire N__52394;
    wire N__52391;
    wire N__52388;
    wire N__52385;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52366;
    wire N__52363;
    wire N__52360;
    wire N__52357;
    wire N__52354;
    wire N__52351;
    wire N__52348;
    wire N__52345;
    wire N__52342;
    wire N__52341;
    wire N__52338;
    wire N__52335;
    wire N__52332;
    wire N__52329;
    wire N__52326;
    wire N__52323;
    wire N__52320;
    wire N__52319;
    wire N__52316;
    wire N__52313;
    wire N__52310;
    wire N__52307;
    wire N__52304;
    wire N__52297;
    wire N__52294;
    wire N__52291;
    wire N__52288;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52276;
    wire N__52273;
    wire N__52272;
    wire N__52269;
    wire N__52266;
    wire N__52263;
    wire N__52258;
    wire N__52257;
    wire N__52254;
    wire N__52251;
    wire N__52248;
    wire N__52247;
    wire N__52242;
    wire N__52239;
    wire N__52234;
    wire N__52233;
    wire N__52230;
    wire N__52229;
    wire N__52226;
    wire N__52223;
    wire N__52220;
    wire N__52215;
    wire N__52212;
    wire N__52207;
    wire N__52206;
    wire N__52205;
    wire N__52202;
    wire N__52199;
    wire N__52196;
    wire N__52193;
    wire N__52190;
    wire N__52183;
    wire N__52180;
    wire N__52177;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52156;
    wire N__52153;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52143;
    wire N__52142;
    wire N__52139;
    wire N__52138;
    wire N__52135;
    wire N__52134;
    wire N__52131;
    wire N__52128;
    wire N__52125;
    wire N__52122;
    wire N__52121;
    wire N__52118;
    wire N__52115;
    wire N__52108;
    wire N__52107;
    wire N__52104;
    wire N__52101;
    wire N__52098;
    wire N__52095;
    wire N__52092;
    wire N__52091;
    wire N__52090;
    wire N__52087;
    wire N__52084;
    wire N__52077;
    wire N__52072;
    wire N__52069;
    wire N__52066;
    wire N__52063;
    wire N__52060;
    wire N__52057;
    wire N__52054;
    wire N__52051;
    wire N__52048;
    wire N__52039;
    wire N__52036;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52024;
    wire N__52021;
    wire N__52018;
    wire N__52015;
    wire N__52012;
    wire N__52009;
    wire N__52006;
    wire N__52003;
    wire N__52000;
    wire N__51999;
    wire N__51996;
    wire N__51993;
    wire N__51990;
    wire N__51985;
    wire N__51982;
    wire N__51981;
    wire N__51980;
    wire N__51977;
    wire N__51974;
    wire N__51971;
    wire N__51968;
    wire N__51965;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51949;
    wire N__51948;
    wire N__51945;
    wire N__51944;
    wire N__51941;
    wire N__51938;
    wire N__51933;
    wire N__51928;
    wire N__51925;
    wire N__51924;
    wire N__51921;
    wire N__51918;
    wire N__51917;
    wire N__51914;
    wire N__51911;
    wire N__51908;
    wire N__51901;
    wire N__51898;
    wire N__51895;
    wire N__51892;
    wire N__51889;
    wire N__51886;
    wire N__51883;
    wire N__51880;
    wire N__51877;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51865;
    wire N__51862;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51850;
    wire N__51847;
    wire N__51844;
    wire N__51841;
    wire N__51838;
    wire N__51837;
    wire N__51834;
    wire N__51831;
    wire N__51830;
    wire N__51829;
    wire N__51824;
    wire N__51823;
    wire N__51822;
    wire N__51821;
    wire N__51818;
    wire N__51815;
    wire N__51812;
    wire N__51809;
    wire N__51808;
    wire N__51807;
    wire N__51804;
    wire N__51801;
    wire N__51800;
    wire N__51797;
    wire N__51792;
    wire N__51789;
    wire N__51786;
    wire N__51785;
    wire N__51784;
    wire N__51781;
    wire N__51780;
    wire N__51779;
    wire N__51774;
    wire N__51771;
    wire N__51768;
    wire N__51765;
    wire N__51762;
    wire N__51755;
    wire N__51752;
    wire N__51747;
    wire N__51730;
    wire N__51729;
    wire N__51726;
    wire N__51725;
    wire N__51722;
    wire N__51719;
    wire N__51716;
    wire N__51713;
    wire N__51708;
    wire N__51703;
    wire N__51700;
    wire N__51699;
    wire N__51696;
    wire N__51693;
    wire N__51690;
    wire N__51685;
    wire N__51682;
    wire N__51679;
    wire N__51676;
    wire N__51673;
    wire N__51670;
    wire N__51667;
    wire N__51664;
    wire N__51661;
    wire N__51658;
    wire N__51655;
    wire N__51652;
    wire N__51649;
    wire N__51646;
    wire N__51645;
    wire N__51642;
    wire N__51639;
    wire N__51636;
    wire N__51633;
    wire N__51630;
    wire N__51625;
    wire N__51624;
    wire N__51623;
    wire N__51620;
    wire N__51615;
    wire N__51614;
    wire N__51609;
    wire N__51606;
    wire N__51601;
    wire N__51598;
    wire N__51595;
    wire N__51592;
    wire N__51589;
    wire N__51586;
    wire N__51585;
    wire N__51582;
    wire N__51579;
    wire N__51574;
    wire N__51571;
    wire N__51568;
    wire N__51567;
    wire N__51566;
    wire N__51563;
    wire N__51560;
    wire N__51557;
    wire N__51554;
    wire N__51547;
    wire N__51546;
    wire N__51543;
    wire N__51542;
    wire N__51539;
    wire N__51536;
    wire N__51531;
    wire N__51528;
    wire N__51525;
    wire N__51522;
    wire N__51519;
    wire N__51514;
    wire N__51511;
    wire N__51508;
    wire N__51505;
    wire N__51502;
    wire N__51501;
    wire N__51498;
    wire N__51495;
    wire N__51492;
    wire N__51489;
    wire N__51486;
    wire N__51483;
    wire N__51478;
    wire N__51475;
    wire N__51472;
    wire N__51471;
    wire N__51470;
    wire N__51469;
    wire N__51462;
    wire N__51459;
    wire N__51454;
    wire N__51451;
    wire N__51450;
    wire N__51447;
    wire N__51446;
    wire N__51445;
    wire N__51444;
    wire N__51441;
    wire N__51432;
    wire N__51429;
    wire N__51424;
    wire N__51423;
    wire N__51422;
    wire N__51417;
    wire N__51414;
    wire N__51409;
    wire N__51406;
    wire N__51403;
    wire N__51400;
    wire N__51397;
    wire N__51396;
    wire N__51393;
    wire N__51390;
    wire N__51387;
    wire N__51384;
    wire N__51381;
    wire N__51380;
    wire N__51377;
    wire N__51374;
    wire N__51371;
    wire N__51364;
    wire N__51363;
    wire N__51362;
    wire N__51361;
    wire N__51360;
    wire N__51355;
    wire N__51354;
    wire N__51353;
    wire N__51352;
    wire N__51349;
    wire N__51348;
    wire N__51343;
    wire N__51340;
    wire N__51339;
    wire N__51338;
    wire N__51331;
    wire N__51328;
    wire N__51325;
    wire N__51324;
    wire N__51323;
    wire N__51320;
    wire N__51317;
    wire N__51314;
    wire N__51311;
    wire N__51310;
    wire N__51307;
    wire N__51302;
    wire N__51299;
    wire N__51296;
    wire N__51289;
    wire N__51284;
    wire N__51283;
    wire N__51280;
    wire N__51277;
    wire N__51268;
    wire N__51265;
    wire N__51262;
    wire N__51259;
    wire N__51256;
    wire N__51247;
    wire N__51244;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51225;
    wire N__51224;
    wire N__51223;
    wire N__51220;
    wire N__51219;
    wire N__51216;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51204;
    wire N__51197;
    wire N__51192;
    wire N__51189;
    wire N__51184;
    wire N__51181;
    wire N__51178;
    wire N__51175;
    wire N__51172;
    wire N__51169;
    wire N__51168;
    wire N__51167;
    wire N__51166;
    wire N__51165;
    wire N__51164;
    wire N__51161;
    wire N__51158;
    wire N__51153;
    wire N__51148;
    wire N__51141;
    wire N__51136;
    wire N__51133;
    wire N__51130;
    wire N__51127;
    wire N__51124;
    wire N__51121;
    wire N__51118;
    wire N__51115;
    wire N__51114;
    wire N__51111;
    wire N__51108;
    wire N__51103;
    wire N__51100;
    wire N__51097;
    wire N__51094;
    wire N__51093;
    wire N__51090;
    wire N__51087;
    wire N__51082;
    wire N__51079;
    wire N__51076;
    wire N__51075;
    wire N__51072;
    wire N__51069;
    wire N__51066;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51052;
    wire N__51049;
    wire N__51046;
    wire N__51045;
    wire N__51042;
    wire N__51039;
    wire N__51036;
    wire N__51033;
    wire N__51028;
    wire N__51025;
    wire N__51022;
    wire N__51019;
    wire N__51016;
    wire N__51013;
    wire N__51010;
    wire N__51007;
    wire N__51004;
    wire N__51001;
    wire N__50998;
    wire N__50995;
    wire N__50992;
    wire N__50989;
    wire N__50986;
    wire N__50983;
    wire N__50980;
    wire N__50977;
    wire N__50974;
    wire N__50971;
    wire N__50968;
    wire N__50965;
    wire N__50962;
    wire N__50959;
    wire N__50956;
    wire N__50953;
    wire N__50950;
    wire N__50949;
    wire N__50946;
    wire N__50943;
    wire N__50938;
    wire N__50937;
    wire N__50934;
    wire N__50933;
    wire N__50930;
    wire N__50927;
    wire N__50924;
    wire N__50917;
    wire N__50914;
    wire N__50911;
    wire N__50908;
    wire N__50905;
    wire N__50902;
    wire N__50899;
    wire N__50896;
    wire N__50893;
    wire N__50892;
    wire N__50891;
    wire N__50890;
    wire N__50889;
    wire N__50888;
    wire N__50887;
    wire N__50886;
    wire N__50885;
    wire N__50880;
    wire N__50877;
    wire N__50872;
    wire N__50865;
    wire N__50862;
    wire N__50859;
    wire N__50858;
    wire N__50853;
    wire N__50850;
    wire N__50847;
    wire N__50844;
    wire N__50841;
    wire N__50836;
    wire N__50833;
    wire N__50828;
    wire N__50825;
    wire N__50820;
    wire N__50815;
    wire N__50814;
    wire N__50809;
    wire N__50808;
    wire N__50807;
    wire N__50804;
    wire N__50801;
    wire N__50798;
    wire N__50797;
    wire N__50794;
    wire N__50791;
    wire N__50788;
    wire N__50785;
    wire N__50776;
    wire N__50775;
    wire N__50772;
    wire N__50771;
    wire N__50770;
    wire N__50769;
    wire N__50768;
    wire N__50765;
    wire N__50764;
    wire N__50763;
    wire N__50760;
    wire N__50755;
    wire N__50754;
    wire N__50753;
    wire N__50748;
    wire N__50745;
    wire N__50742;
    wire N__50739;
    wire N__50738;
    wire N__50737;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50723;
    wire N__50722;
    wire N__50719;
    wire N__50716;
    wire N__50711;
    wire N__50704;
    wire N__50697;
    wire N__50694;
    wire N__50689;
    wire N__50688;
    wire N__50685;
    wire N__50682;
    wire N__50679;
    wire N__50676;
    wire N__50669;
    wire N__50666;
    wire N__50659;
    wire N__50656;
    wire N__50653;
    wire N__50644;
    wire N__50641;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50633;
    wire N__50630;
    wire N__50627;
    wire N__50624;
    wire N__50621;
    wire N__50614;
    wire N__50611;
    wire N__50610;
    wire N__50609;
    wire N__50608;
    wire N__50605;
    wire N__50600;
    wire N__50599;
    wire N__50596;
    wire N__50595;
    wire N__50594;
    wire N__50593;
    wire N__50592;
    wire N__50587;
    wire N__50584;
    wire N__50581;
    wire N__50578;
    wire N__50573;
    wire N__50570;
    wire N__50567;
    wire N__50554;
    wire N__50553;
    wire N__50552;
    wire N__50551;
    wire N__50550;
    wire N__50549;
    wire N__50548;
    wire N__50547;
    wire N__50546;
    wire N__50545;
    wire N__50544;
    wire N__50543;
    wire N__50542;
    wire N__50541;
    wire N__50540;
    wire N__50539;
    wire N__50538;
    wire N__50537;
    wire N__50536;
    wire N__50535;
    wire N__50532;
    wire N__50521;
    wire N__50510;
    wire N__50507;
    wire N__50498;
    wire N__50495;
    wire N__50492;
    wire N__50491;
    wire N__50490;
    wire N__50485;
    wire N__50480;
    wire N__50477;
    wire N__50474;
    wire N__50471;
    wire N__50466;
    wire N__50461;
    wire N__50460;
    wire N__50459;
    wire N__50456;
    wire N__50455;
    wire N__50452;
    wire N__50449;
    wire N__50440;
    wire N__50435;
    wire N__50432;
    wire N__50429;
    wire N__50416;
    wire N__50415;
    wire N__50414;
    wire N__50413;
    wire N__50412;
    wire N__50411;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50407;
    wire N__50406;
    wire N__50405;
    wire N__50404;
    wire N__50403;
    wire N__50390;
    wire N__50379;
    wire N__50376;
    wire N__50375;
    wire N__50374;
    wire N__50373;
    wire N__50372;
    wire N__50369;
    wire N__50368;
    wire N__50365;
    wire N__50364;
    wire N__50363;
    wire N__50360;
    wire N__50357;
    wire N__50354;
    wire N__50345;
    wire N__50342;
    wire N__50339;
    wire N__50336;
    wire N__50331;
    wire N__50330;
    wire N__50329;
    wire N__50326;
    wire N__50319;
    wire N__50318;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50311;
    wire N__50304;
    wire N__50301;
    wire N__50298;
    wire N__50293;
    wire N__50288;
    wire N__50281;
    wire N__50276;
    wire N__50263;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50203;
    wire N__50200;
    wire N__50199;
    wire N__50198;
    wire N__50195;
    wire N__50192;
    wire N__50189;
    wire N__50188;
    wire N__50185;
    wire N__50180;
    wire N__50177;
    wire N__50174;
    wire N__50169;
    wire N__50168;
    wire N__50165;
    wire N__50162;
    wire N__50159;
    wire N__50156;
    wire N__50153;
    wire N__50150;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50127;
    wire N__50124;
    wire N__50121;
    wire N__50118;
    wire N__50117;
    wire N__50114;
    wire N__50111;
    wire N__50108;
    wire N__50105;
    wire N__50102;
    wire N__50097;
    wire N__50092;
    wire N__50089;
    wire N__50086;
    wire N__50083;
    wire N__50082;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50068;
    wire N__50065;
    wire N__50062;
    wire N__50059;
    wire N__50058;
    wire N__50055;
    wire N__50052;
    wire N__50049;
    wire N__50044;
    wire N__50041;
    wire N__50038;
    wire N__50035;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50020;
    wire N__50019;
    wire N__50018;
    wire N__50017;
    wire N__50014;
    wire N__50013;
    wire N__50010;
    wire N__50007;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49995;
    wire N__49992;
    wire N__49989;
    wire N__49986;
    wire N__49983;
    wire N__49978;
    wire N__49973;
    wire N__49970;
    wire N__49967;
    wire N__49964;
    wire N__49957;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49947;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49939;
    wire N__49936;
    wire N__49933;
    wire N__49930;
    wire N__49925;
    wire N__49922;
    wire N__49919;
    wire N__49912;
    wire N__49909;
    wire N__49906;
    wire N__49903;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49888;
    wire N__49885;
    wire N__49884;
    wire N__49881;
    wire N__49878;
    wire N__49875;
    wire N__49872;
    wire N__49867;
    wire N__49866;
    wire N__49863;
    wire N__49860;
    wire N__49857;
    wire N__49852;
    wire N__49849;
    wire N__49848;
    wire N__49845;
    wire N__49844;
    wire N__49841;
    wire N__49838;
    wire N__49835;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49819;
    wire N__49816;
    wire N__49815;
    wire N__49812;
    wire N__49811;
    wire N__49808;
    wire N__49805;
    wire N__49802;
    wire N__49795;
    wire N__49792;
    wire N__49789;
    wire N__49786;
    wire N__49783;
    wire N__49782;
    wire N__49779;
    wire N__49778;
    wire N__49775;
    wire N__49772;
    wire N__49769;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49753;
    wire N__49750;
    wire N__49747;
    wire N__49746;
    wire N__49743;
    wire N__49742;
    wire N__49739;
    wire N__49736;
    wire N__49733;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49719;
    wire N__49716;
    wire N__49713;
    wire N__49710;
    wire N__49705;
    wire N__49702;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49687;
    wire N__49684;
    wire N__49683;
    wire N__49682;
    wire N__49679;
    wire N__49674;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49656;
    wire N__49655;
    wire N__49652;
    wire N__49647;
    wire N__49642;
    wire N__49639;
    wire N__49636;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49624;
    wire N__49621;
    wire N__49618;
    wire N__49615;
    wire N__49612;
    wire N__49609;
    wire N__49606;
    wire N__49605;
    wire N__49602;
    wire N__49599;
    wire N__49596;
    wire N__49591;
    wire N__49588;
    wire N__49585;
    wire N__49582;
    wire N__49579;
    wire N__49576;
    wire N__49573;
    wire N__49570;
    wire N__49569;
    wire N__49568;
    wire N__49567;
    wire N__49564;
    wire N__49563;
    wire N__49562;
    wire N__49561;
    wire N__49560;
    wire N__49559;
    wire N__49552;
    wire N__49549;
    wire N__49546;
    wire N__49543;
    wire N__49538;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49522;
    wire N__49519;
    wire N__49518;
    wire N__49515;
    wire N__49510;
    wire N__49507;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49499;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49479;
    wire N__49474;
    wire N__49471;
    wire N__49462;
    wire N__49459;
    wire N__49458;
    wire N__49457;
    wire N__49454;
    wire N__49451;
    wire N__49448;
    wire N__49443;
    wire N__49438;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49424;
    wire N__49421;
    wire N__49418;
    wire N__49413;
    wire N__49412;
    wire N__49409;
    wire N__49406;
    wire N__49403;
    wire N__49396;
    wire N__49393;
    wire N__49392;
    wire N__49389;
    wire N__49388;
    wire N__49385;
    wire N__49382;
    wire N__49379;
    wire N__49372;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49362;
    wire N__49359;
    wire N__49356;
    wire N__49351;
    wire N__49348;
    wire N__49345;
    wire N__49342;
    wire N__49339;
    wire N__49336;
    wire N__49333;
    wire N__49330;
    wire N__49327;
    wire N__49326;
    wire N__49323;
    wire N__49322;
    wire N__49319;
    wire N__49318;
    wire N__49315;
    wire N__49312;
    wire N__49311;
    wire N__49308;
    wire N__49305;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49293;
    wire N__49292;
    wire N__49289;
    wire N__49286;
    wire N__49283;
    wire N__49280;
    wire N__49277;
    wire N__49274;
    wire N__49273;
    wire N__49268;
    wire N__49261;
    wire N__49258;
    wire N__49255;
    wire N__49250;
    wire N__49243;
    wire N__49240;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49232;
    wire N__49231;
    wire N__49230;
    wire N__49225;
    wire N__49222;
    wire N__49221;
    wire N__49218;
    wire N__49215;
    wire N__49214;
    wire N__49211;
    wire N__49208;
    wire N__49205;
    wire N__49202;
    wire N__49199;
    wire N__49196;
    wire N__49193;
    wire N__49188;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49165;
    wire N__49162;
    wire N__49159;
    wire N__49150;
    wire N__49147;
    wire N__49146;
    wire N__49143;
    wire N__49142;
    wire N__49141;
    wire N__49140;
    wire N__49137;
    wire N__49134;
    wire N__49133;
    wire N__49130;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49106;
    wire N__49103;
    wire N__49100;
    wire N__49097;
    wire N__49094;
    wire N__49091;
    wire N__49088;
    wire N__49087;
    wire N__49082;
    wire N__49079;
    wire N__49076;
    wire N__49073;
    wire N__49066;
    wire N__49063;
    wire N__49060;
    wire N__49057;
    wire N__49052;
    wire N__49047;
    wire N__49042;
    wire N__49039;
    wire N__49030;
    wire N__49027;
    wire N__49026;
    wire N__49023;
    wire N__49020;
    wire N__49017;
    wire N__49012;
    wire N__49009;
    wire N__49006;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48993;
    wire N__48990;
    wire N__48987;
    wire N__48986;
    wire N__48983;
    wire N__48980;
    wire N__48977;
    wire N__48974;
    wire N__48971;
    wire N__48964;
    wire N__48961;
    wire N__48958;
    wire N__48957;
    wire N__48954;
    wire N__48951;
    wire N__48946;
    wire N__48943;
    wire N__48942;
    wire N__48941;
    wire N__48938;
    wire N__48935;
    wire N__48932;
    wire N__48929;
    wire N__48926;
    wire N__48923;
    wire N__48920;
    wire N__48917;
    wire N__48912;
    wire N__48909;
    wire N__48906;
    wire N__48901;
    wire N__48900;
    wire N__48897;
    wire N__48894;
    wire N__48889;
    wire N__48886;
    wire N__48883;
    wire N__48880;
    wire N__48879;
    wire N__48876;
    wire N__48873;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48867;
    wire N__48864;
    wire N__48861;
    wire N__48858;
    wire N__48857;
    wire N__48854;
    wire N__48849;
    wire N__48846;
    wire N__48843;
    wire N__48840;
    wire N__48833;
    wire N__48830;
    wire N__48827;
    wire N__48824;
    wire N__48821;
    wire N__48814;
    wire N__48811;
    wire N__48810;
    wire N__48809;
    wire N__48808;
    wire N__48807;
    wire N__48804;
    wire N__48801;
    wire N__48800;
    wire N__48799;
    wire N__48798;
    wire N__48791;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48777;
    wire N__48774;
    wire N__48771;
    wire N__48768;
    wire N__48765;
    wire N__48762;
    wire N__48759;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48734;
    wire N__48731;
    wire N__48724;
    wire N__48721;
    wire N__48720;
    wire N__48719;
    wire N__48716;
    wire N__48713;
    wire N__48710;
    wire N__48707;
    wire N__48706;
    wire N__48699;
    wire N__48696;
    wire N__48693;
    wire N__48692;
    wire N__48689;
    wire N__48686;
    wire N__48683;
    wire N__48680;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48642;
    wire N__48639;
    wire N__48636;
    wire N__48633;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48609;
    wire N__48606;
    wire N__48603;
    wire N__48602;
    wire N__48597;
    wire N__48594;
    wire N__48591;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48561;
    wire N__48558;
    wire N__48555;
    wire N__48552;
    wire N__48549;
    wire N__48544;
    wire N__48543;
    wire N__48542;
    wire N__48541;
    wire N__48540;
    wire N__48539;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48535;
    wire N__48534;
    wire N__48533;
    wire N__48532;
    wire N__48523;
    wire N__48514;
    wire N__48513;
    wire N__48512;
    wire N__48511;
    wire N__48510;
    wire N__48509;
    wire N__48508;
    wire N__48507;
    wire N__48506;
    wire N__48505;
    wire N__48504;
    wire N__48503;
    wire N__48502;
    wire N__48493;
    wire N__48490;
    wire N__48487;
    wire N__48484;
    wire N__48475;
    wire N__48466;
    wire N__48457;
    wire N__48452;
    wire N__48439;
    wire N__48436;
    wire N__48435;
    wire N__48432;
    wire N__48429;
    wire N__48426;
    wire N__48421;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48414;
    wire N__48413;
    wire N__48412;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48408;
    wire N__48407;
    wire N__48406;
    wire N__48405;
    wire N__48404;
    wire N__48403;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48397;
    wire N__48396;
    wire N__48395;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48345;
    wire N__48342;
    wire N__48339;
    wire N__48338;
    wire N__48337;
    wire N__48332;
    wire N__48329;
    wire N__48326;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48314;
    wire N__48311;
    wire N__48308;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48291;
    wire N__48288;
    wire N__48285;
    wire N__48282;
    wire N__48279;
    wire N__48276;
    wire N__48271;
    wire N__48268;
    wire N__48265;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48235;
    wire N__48234;
    wire N__48231;
    wire N__48228;
    wire N__48225;
    wire N__48220;
    wire N__48217;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48205;
    wire N__48202;
    wire N__48201;
    wire N__48198;
    wire N__48195;
    wire N__48192;
    wire N__48187;
    wire N__48184;
    wire N__48183;
    wire N__48180;
    wire N__48177;
    wire N__48174;
    wire N__48169;
    wire N__48166;
    wire N__48165;
    wire N__48162;
    wire N__48159;
    wire N__48154;
    wire N__48151;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48139;
    wire N__48136;
    wire N__48135;
    wire N__48132;
    wire N__48129;
    wire N__48124;
    wire N__48121;
    wire N__48120;
    wire N__48117;
    wire N__48114;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48088;
    wire N__48085;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48070;
    wire N__48067;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48055;
    wire N__48052;
    wire N__48051;
    wire N__48048;
    wire N__48045;
    wire N__48040;
    wire N__48037;
    wire N__48036;
    wire N__48033;
    wire N__48030;
    wire N__48025;
    wire N__48022;
    wire N__48021;
    wire N__48018;
    wire N__48015;
    wire N__48010;
    wire N__48007;
    wire N__48006;
    wire N__48003;
    wire N__48000;
    wire N__47995;
    wire N__47992;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47980;
    wire N__47977;
    wire N__47974;
    wire N__47973;
    wire N__47970;
    wire N__47967;
    wire N__47962;
    wire N__47959;
    wire N__47958;
    wire N__47955;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47945;
    wire N__47938;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47926;
    wire N__47923;
    wire N__47920;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47908;
    wire N__47905;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47893;
    wire N__47890;
    wire N__47887;
    wire N__47884;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47872;
    wire N__47869;
    wire N__47868;
    wire N__47865;
    wire N__47862;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47836;
    wire N__47833;
    wire N__47832;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47818;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47810;
    wire N__47807;
    wire N__47804;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47788;
    wire N__47785;
    wire N__47784;
    wire N__47783;
    wire N__47780;
    wire N__47777;
    wire N__47776;
    wire N__47775;
    wire N__47774;
    wire N__47773;
    wire N__47772;
    wire N__47771;
    wire N__47770;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47742;
    wire N__47739;
    wire N__47736;
    wire N__47733;
    wire N__47728;
    wire N__47719;
    wire N__47710;
    wire N__47707;
    wire N__47704;
    wire N__47699;
    wire N__47692;
    wire N__47691;
    wire N__47688;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47674;
    wire N__47671;
    wire N__47668;
    wire N__47665;
    wire N__47662;
    wire N__47661;
    wire N__47660;
    wire N__47659;
    wire N__47656;
    wire N__47655;
    wire N__47648;
    wire N__47645;
    wire N__47642;
    wire N__47637;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47614;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47584;
    wire N__47583;
    wire N__47582;
    wire N__47579;
    wire N__47576;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47555;
    wire N__47550;
    wire N__47547;
    wire N__47542;
    wire N__47541;
    wire N__47538;
    wire N__47535;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47518;
    wire N__47517;
    wire N__47516;
    wire N__47515;
    wire N__47512;
    wire N__47509;
    wire N__47506;
    wire N__47503;
    wire N__47498;
    wire N__47495;
    wire N__47492;
    wire N__47489;
    wire N__47486;
    wire N__47479;
    wire N__47476;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47451;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47424;
    wire N__47419;
    wire N__47416;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47402;
    wire N__47397;
    wire N__47392;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47380;
    wire N__47377;
    wire N__47374;
    wire N__47373;
    wire N__47368;
    wire N__47367;
    wire N__47364;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47356;
    wire N__47353;
    wire N__47352;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47329;
    wire N__47324;
    wire N__47317;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47296;
    wire N__47293;
    wire N__47290;
    wire N__47289;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47269;
    wire N__47268;
    wire N__47267;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47246;
    wire N__47243;
    wire N__47236;
    wire N__47233;
    wire N__47232;
    wire N__47229;
    wire N__47226;
    wire N__47223;
    wire N__47220;
    wire N__47219;
    wire N__47214;
    wire N__47211;
    wire N__47208;
    wire N__47203;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47175;
    wire N__47172;
    wire N__47169;
    wire N__47164;
    wire N__47161;
    wire N__47158;
    wire N__47155;
    wire N__47154;
    wire N__47151;
    wire N__47148;
    wire N__47145;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47124;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47099;
    wire N__47094;
    wire N__47091;
    wire N__47088;
    wire N__47085;
    wire N__47080;
    wire N__47077;
    wire N__47076;
    wire N__47073;
    wire N__47070;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47052;
    wire N__47047;
    wire N__47044;
    wire N__47041;
    wire N__47038;
    wire N__47035;
    wire N__47032;
    wire N__47031;
    wire N__47030;
    wire N__47027;
    wire N__47022;
    wire N__47017;
    wire N__47014;
    wire N__47013;
    wire N__47010;
    wire N__47009;
    wire N__47006;
    wire N__47003;
    wire N__47000;
    wire N__46997;
    wire N__46990;
    wire N__46987;
    wire N__46984;
    wire N__46981;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46934;
    wire N__46931;
    wire N__46924;
    wire N__46921;
    wire N__46920;
    wire N__46917;
    wire N__46914;
    wire N__46911;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46889;
    wire N__46886;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46851;
    wire N__46850;
    wire N__46849;
    wire N__46848;
    wire N__46847;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46843;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46831;
    wire N__46826;
    wire N__46821;
    wire N__46820;
    wire N__46819;
    wire N__46818;
    wire N__46817;
    wire N__46814;
    wire N__46811;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46799;
    wire N__46794;
    wire N__46791;
    wire N__46788;
    wire N__46785;
    wire N__46782;
    wire N__46775;
    wire N__46768;
    wire N__46765;
    wire N__46750;
    wire N__46749;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46739;
    wire N__46738;
    wire N__46737;
    wire N__46736;
    wire N__46733;
    wire N__46730;
    wire N__46727;
    wire N__46720;
    wire N__46717;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46701;
    wire N__46698;
    wire N__46695;
    wire N__46690;
    wire N__46687;
    wire N__46684;
    wire N__46681;
    wire N__46678;
    wire N__46675;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46662;
    wire N__46659;
    wire N__46658;
    wire N__46655;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46647;
    wire N__46646;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46636;
    wire N__46633;
    wire N__46630;
    wire N__46629;
    wire N__46626;
    wire N__46623;
    wire N__46622;
    wire N__46621;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46602;
    wire N__46599;
    wire N__46596;
    wire N__46593;
    wire N__46588;
    wire N__46585;
    wire N__46582;
    wire N__46575;
    wire N__46572;
    wire N__46569;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46555;
    wire N__46552;
    wire N__46541;
    wire N__46534;
    wire N__46531;
    wire N__46530;
    wire N__46527;
    wire N__46524;
    wire N__46521;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46511;
    wire N__46504;
    wire N__46501;
    wire N__46498;
    wire N__46495;
    wire N__46492;
    wire N__46489;
    wire N__46486;
    wire N__46483;
    wire N__46482;
    wire N__46481;
    wire N__46478;
    wire N__46475;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46462;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46431;
    wire N__46428;
    wire N__46427;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46408;
    wire N__46405;
    wire N__46404;
    wire N__46403;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46391;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46354;
    wire N__46353;
    wire N__46352;
    wire N__46351;
    wire N__46350;
    wire N__46349;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46306;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46290;
    wire N__46285;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46237;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46219;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46204;
    wire N__46203;
    wire N__46202;
    wire N__46201;
    wire N__46200;
    wire N__46199;
    wire N__46196;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46164;
    wire N__46163;
    wire N__46160;
    wire N__46157;
    wire N__46150;
    wire N__46145;
    wire N__46142;
    wire N__46139;
    wire N__46132;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46109;
    wire N__46106;
    wire N__46101;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46058;
    wire N__46053;
    wire N__46050;
    wire N__46045;
    wire N__46042;
    wire N__46039;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46009;
    wire N__46008;
    wire N__46007;
    wire N__46002;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45996;
    wire N__45995;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45981;
    wire N__45978;
    wire N__45977;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45955;
    wire N__45954;
    wire N__45953;
    wire N__45950;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45942;
    wire N__45941;
    wire N__45940;
    wire N__45937;
    wire N__45934;
    wire N__45933;
    wire N__45930;
    wire N__45925;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45911;
    wire N__45904;
    wire N__45901;
    wire N__45898;
    wire N__45891;
    wire N__45886;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45874;
    wire N__45871;
    wire N__45868;
    wire N__45865;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45838;
    wire N__45835;
    wire N__45832;
    wire N__45829;
    wire N__45826;
    wire N__45823;
    wire N__45820;
    wire N__45817;
    wire N__45814;
    wire N__45811;
    wire N__45810;
    wire N__45809;
    wire N__45806;
    wire N__45801;
    wire N__45800;
    wire N__45799;
    wire N__45798;
    wire N__45797;
    wire N__45794;
    wire N__45791;
    wire N__45790;
    wire N__45789;
    wire N__45788;
    wire N__45787;
    wire N__45784;
    wire N__45783;
    wire N__45782;
    wire N__45781;
    wire N__45774;
    wire N__45769;
    wire N__45760;
    wire N__45757;
    wire N__45754;
    wire N__45749;
    wire N__45736;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45700;
    wire N__45699;
    wire N__45696;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45658;
    wire N__45657;
    wire N__45654;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45641;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45616;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45601;
    wire N__45598;
    wire N__45595;
    wire N__45592;
    wire N__45589;
    wire N__45586;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45569;
    wire N__45566;
    wire N__45563;
    wire N__45562;
    wire N__45559;
    wire N__45558;
    wire N__45557;
    wire N__45556;
    wire N__45553;
    wire N__45550;
    wire N__45547;
    wire N__45544;
    wire N__45537;
    wire N__45532;
    wire N__45527;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45496;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45455;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45437;
    wire N__45430;
    wire N__45427;
    wire N__45426;
    wire N__45423;
    wire N__45422;
    wire N__45421;
    wire N__45418;
    wire N__45415;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45401;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45380;
    wire N__45373;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45349;
    wire N__45340;
    wire N__45339;
    wire N__45336;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45328;
    wire N__45327;
    wire N__45326;
    wire N__45325;
    wire N__45322;
    wire N__45319;
    wire N__45316;
    wire N__45313;
    wire N__45312;
    wire N__45309;
    wire N__45304;
    wire N__45301;
    wire N__45298;
    wire N__45295;
    wire N__45292;
    wire N__45289;
    wire N__45284;
    wire N__45283;
    wire N__45276;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45259;
    wire N__45254;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45223;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45211;
    wire N__45208;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45169;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45154;
    wire N__45151;
    wire N__45148;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45136;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45112;
    wire N__45111;
    wire N__45106;
    wire N__45103;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45079;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45007;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44999;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44974;
    wire N__44971;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44941;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44926;
    wire N__44925;
    wire N__44920;
    wire N__44917;
    wire N__44916;
    wire N__44911;
    wire N__44908;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44875;
    wire N__44872;
    wire N__44869;
    wire N__44866;
    wire N__44863;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44803;
    wire N__44800;
    wire N__44797;
    wire N__44794;
    wire N__44791;
    wire N__44788;
    wire N__44785;
    wire N__44784;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44774;
    wire N__44769;
    wire N__44764;
    wire N__44763;
    wire N__44760;
    wire N__44759;
    wire N__44756;
    wire N__44751;
    wire N__44748;
    wire N__44743;
    wire N__44742;
    wire N__44739;
    wire N__44738;
    wire N__44737;
    wire N__44734;
    wire N__44729;
    wire N__44726;
    wire N__44719;
    wire N__44716;
    wire N__44715;
    wire N__44714;
    wire N__44711;
    wire N__44708;
    wire N__44707;
    wire N__44704;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44684;
    wire N__44681;
    wire N__44678;
    wire N__44677;
    wire N__44674;
    wire N__44665;
    wire N__44662;
    wire N__44657;
    wire N__44654;
    wire N__44647;
    wire N__44646;
    wire N__44643;
    wire N__44642;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44632;
    wire N__44631;
    wire N__44630;
    wire N__44627;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44617;
    wire N__44614;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44592;
    wire N__44589;
    wire N__44586;
    wire N__44583;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44569;
    wire N__44566;
    wire N__44565;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44540;
    wire N__44527;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44508;
    wire N__44505;
    wire N__44502;
    wire N__44497;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44484;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44464;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44383;
    wire N__44382;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44340;
    wire N__44337;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44296;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44288;
    wire N__44285;
    wire N__44280;
    wire N__44277;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44248;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44230;
    wire N__44229;
    wire N__44228;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44181;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44156;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44140;
    wire N__44137;
    wire N__44134;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44105;
    wire N__44100;
    wire N__44097;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44079;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44044;
    wire N__44041;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44017;
    wire N__44014;
    wire N__44011;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43957;
    wire N__43956;
    wire N__43955;
    wire N__43952;
    wire N__43949;
    wire N__43948;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43940;
    wire N__43939;
    wire N__43934;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43914;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43894;
    wire N__43891;
    wire N__43886;
    wire N__43873;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43848;
    wire N__43843;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43818;
    wire N__43815;
    wire N__43808;
    wire N__43805;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43671;
    wire N__43668;
    wire N__43665;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43650;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43633;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43618;
    wire N__43617;
    wire N__43616;
    wire N__43613;
    wire N__43612;
    wire N__43611;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43578;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43497;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43285;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43240;
    wire N__43237;
    wire N__43234;
    wire N__43231;
    wire N__43228;
    wire N__43227;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43071;
    wire N__43068;
    wire N__43065;
    wire N__43060;
    wire N__43057;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43042;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42982;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42972;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42960;
    wire N__42957;
    wire N__42954;
    wire N__42949;
    wire N__42948;
    wire N__42945;
    wire N__42942;
    wire N__42937;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42922;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42892;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42880;
    wire N__42879;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42865;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42846;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42826;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42808;
    wire N__42805;
    wire N__42802;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42792;
    wire N__42789;
    wire N__42786;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42759;
    wire N__42758;
    wire N__42757;
    wire N__42754;
    wire N__42753;
    wire N__42750;
    wire N__42749;
    wire N__42748;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42740;
    wire N__42739;
    wire N__42738;
    wire N__42737;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42721;
    wire N__42720;
    wire N__42719;
    wire N__42718;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42698;
    wire N__42697;
    wire N__42696;
    wire N__42695;
    wire N__42694;
    wire N__42691;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42679;
    wire N__42676;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42617;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42584;
    wire N__42581;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42565;
    wire N__42560;
    wire N__42555;
    wire N__42548;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42520;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42499;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42491;
    wire N__42490;
    wire N__42489;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42469;
    wire N__42466;
    wire N__42463;
    wire N__42460;
    wire N__42453;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42430;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42418;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42406;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42391;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42379;
    wire N__42376;
    wire N__42373;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42351;
    wire N__42350;
    wire N__42347;
    wire N__42344;
    wire N__42341;
    wire N__42334;
    wire N__42333;
    wire N__42332;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42306;
    wire N__42301;
    wire N__42298;
    wire N__42295;
    wire N__42292;
    wire N__42289;
    wire N__42286;
    wire N__42283;
    wire N__42280;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42268;
    wire N__42265;
    wire N__42262;
    wire N__42259;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42208;
    wire N__42207;
    wire N__42206;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42190;
    wire N__42187;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42157;
    wire N__42154;
    wire N__42153;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42133;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42110;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42096;
    wire N__42095;
    wire N__42092;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42076;
    wire N__42073;
    wire N__42070;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42056;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42044;
    wire N__42041;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41986;
    wire N__41985;
    wire N__41982;
    wire N__41981;
    wire N__41980;
    wire N__41977;
    wire N__41974;
    wire N__41971;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41963;
    wire N__41958;
    wire N__41955;
    wire N__41950;
    wire N__41947;
    wire N__41940;
    wire N__41935;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41903;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41872;
    wire N__41871;
    wire N__41868;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41846;
    wire N__41843;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41790;
    wire N__41789;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41773;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41763;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41728;
    wire N__41725;
    wire N__41722;
    wire N__41719;
    wire N__41718;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41656;
    wire N__41653;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41641;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41626;
    wire N__41625;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41615;
    wire N__41608;
    wire N__41605;
    wire N__41602;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41548;
    wire N__41545;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41533;
    wire N__41530;
    wire N__41527;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41512;
    wire N__41511;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41501;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41487;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41389;
    wire N__41386;
    wire N__41383;
    wire N__41380;
    wire N__41377;
    wire N__41374;
    wire N__41371;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41353;
    wire N__41350;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41273;
    wire N__41266;
    wire N__41265;
    wire N__41262;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41209;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41187;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41172;
    wire N__41169;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41148;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41134;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41067;
    wire N__41066;
    wire N__41063;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41020;
    wire N__41019;
    wire N__41016;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41005;
    wire N__41002;
    wire N__40997;
    wire N__40994;
    wire N__40991;
    wire N__40986;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40974;
    wire N__40973;
    wire N__40970;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40948;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40940;
    wire N__40939;
    wire N__40936;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40925;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40907;
    wire N__40904;
    wire N__40899;
    wire N__40894;
    wire N__40891;
    wire N__40890;
    wire N__40887;
    wire N__40884;
    wire N__40879;
    wire N__40876;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40854;
    wire N__40849;
    wire N__40846;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40834;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40643;
    wire N__40640;
    wire N__40635;
    wire N__40630;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40569;
    wire N__40568;
    wire N__40565;
    wire N__40564;
    wire N__40563;
    wire N__40562;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40539;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40526;
    wire N__40523;
    wire N__40518;
    wire N__40517;
    wire N__40514;
    wire N__40509;
    wire N__40504;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40484;
    wire N__40481;
    wire N__40476;
    wire N__40465;
    wire N__40462;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40432;
    wire N__40429;
    wire N__40426;
    wire N__40425;
    wire N__40424;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40369;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40357;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40345;
    wire N__40342;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40327;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40227;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40204;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40196;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40180;
    wire N__40177;
    wire N__40174;
    wire N__40171;
    wire N__40170;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40120;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40069;
    wire N__40066;
    wire N__40065;
    wire N__40064;
    wire N__40061;
    wire N__40058;
    wire N__40055;
    wire N__40052;
    wire N__40045;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39969;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39931;
    wire N__39928;
    wire N__39927;
    wire N__39926;
    wire N__39923;
    wire N__39920;
    wire N__39917;
    wire N__39910;
    wire N__39909;
    wire N__39908;
    wire N__39905;
    wire N__39902;
    wire N__39899;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39879;
    wire N__39876;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39856;
    wire N__39855;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39840;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39820;
    wire N__39819;
    wire N__39818;
    wire N__39817;
    wire N__39816;
    wire N__39813;
    wire N__39812;
    wire N__39811;
    wire N__39810;
    wire N__39809;
    wire N__39808;
    wire N__39807;
    wire N__39806;
    wire N__39801;
    wire N__39800;
    wire N__39799;
    wire N__39798;
    wire N__39797;
    wire N__39794;
    wire N__39785;
    wire N__39782;
    wire N__39781;
    wire N__39780;
    wire N__39777;
    wire N__39776;
    wire N__39775;
    wire N__39774;
    wire N__39773;
    wire N__39772;
    wire N__39769;
    wire N__39768;
    wire N__39767;
    wire N__39766;
    wire N__39765;
    wire N__39764;
    wire N__39763;
    wire N__39762;
    wire N__39759;
    wire N__39758;
    wire N__39755;
    wire N__39754;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39746;
    wire N__39745;
    wire N__39738;
    wire N__39733;
    wire N__39732;
    wire N__39729;
    wire N__39728;
    wire N__39725;
    wire N__39716;
    wire N__39715;
    wire N__39714;
    wire N__39713;
    wire N__39712;
    wire N__39711;
    wire N__39704;
    wire N__39701;
    wire N__39690;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39664;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39652;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39637;
    wire N__39636;
    wire N__39633;
    wire N__39632;
    wire N__39631;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39623;
    wire N__39622;
    wire N__39621;
    wire N__39620;
    wire N__39619;
    wire N__39618;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39610;
    wire N__39609;
    wire N__39608;
    wire N__39605;
    wire N__39598;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39580;
    wire N__39573;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39557;
    wire N__39556;
    wire N__39555;
    wire N__39554;
    wire N__39553;
    wire N__39552;
    wire N__39551;
    wire N__39550;
    wire N__39549;
    wire N__39548;
    wire N__39545;
    wire N__39542;
    wire N__39537;
    wire N__39534;
    wire N__39523;
    wire N__39520;
    wire N__39513;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39483;
    wire N__39474;
    wire N__39465;
    wire N__39454;
    wire N__39421;
    wire N__39420;
    wire N__39419;
    wire N__39418;
    wire N__39415;
    wire N__39410;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39404;
    wire N__39403;
    wire N__39402;
    wire N__39401;
    wire N__39400;
    wire N__39399;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39387;
    wire N__39386;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39378;
    wire N__39377;
    wire N__39372;
    wire N__39371;
    wire N__39370;
    wire N__39365;
    wire N__39362;
    wire N__39361;
    wire N__39360;
    wire N__39357;
    wire N__39352;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39334;
    wire N__39329;
    wire N__39326;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39310;
    wire N__39305;
    wire N__39302;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39286;
    wire N__39283;
    wire N__39274;
    wire N__39271;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39241;
    wire N__39232;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39209;
    wire N__39206;
    wire N__39201;
    wire N__39196;
    wire N__39193;
    wire N__39192;
    wire N__39191;
    wire N__39188;
    wire N__39183;
    wire N__39178;
    wire N__39177;
    wire N__39174;
    wire N__39173;
    wire N__39172;
    wire N__39171;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39137;
    wire N__39134;
    wire N__39133;
    wire N__39132;
    wire N__39131;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39105;
    wire N__39102;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38983;
    wire N__38980;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38965;
    wire N__38962;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38947;
    wire N__38944;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38929;
    wire N__38926;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38872;
    wire N__38871;
    wire N__38868;
    wire N__38867;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38846;
    wire N__38839;
    wire N__38836;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38821;
    wire N__38818;
    wire N__38817;
    wire N__38816;
    wire N__38813;
    wire N__38808;
    wire N__38803;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38793;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38776;
    wire N__38775;
    wire N__38774;
    wire N__38773;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38759;
    wire N__38758;
    wire N__38757;
    wire N__38754;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38722;
    wire N__38719;
    wire N__38712;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38694;
    wire N__38691;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38676;
    wire N__38673;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38661;
    wire N__38658;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38628;
    wire N__38623;
    wire N__38620;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38584;
    wire N__38583;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38565;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38353;
    wire N__38352;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38334;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38311;
    wire N__38308;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38238;
    wire N__38237;
    wire N__38234;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38216;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38198;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38140;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38118;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38098;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38071;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38036;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38022;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37993;
    wire N__37990;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37941;
    wire N__37940;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37882;
    wire N__37879;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37871;
    wire N__37868;
    wire N__37865;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37839;
    wire N__37838;
    wire N__37837;
    wire N__37836;
    wire N__37833;
    wire N__37832;
    wire N__37831;
    wire N__37830;
    wire N__37825;
    wire N__37824;
    wire N__37823;
    wire N__37822;
    wire N__37821;
    wire N__37816;
    wire N__37815;
    wire N__37814;
    wire N__37811;
    wire N__37810;
    wire N__37807;
    wire N__37802;
    wire N__37801;
    wire N__37800;
    wire N__37797;
    wire N__37796;
    wire N__37795;
    wire N__37794;
    wire N__37793;
    wire N__37792;
    wire N__37791;
    wire N__37790;
    wire N__37789;
    wire N__37786;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37772;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37758;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37748;
    wire N__37747;
    wire N__37746;
    wire N__37745;
    wire N__37744;
    wire N__37743;
    wire N__37740;
    wire N__37737;
    wire N__37732;
    wire N__37723;
    wire N__37718;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37700;
    wire N__37697;
    wire N__37692;
    wire N__37689;
    wire N__37678;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37655;
    wire N__37650;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37599;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37513;
    wire N__37510;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37485;
    wire N__37480;
    wire N__37477;
    wire N__37476;
    wire N__37475;
    wire N__37472;
    wire N__37467;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37444;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37432;
    wire N__37429;
    wire N__37426;
    wire N__37423;
    wire N__37420;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37405;
    wire N__37404;
    wire N__37403;
    wire N__37398;
    wire N__37395;
    wire N__37394;
    wire N__37393;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37382;
    wire N__37381;
    wire N__37376;
    wire N__37373;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37351;
    wire N__37348;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37333;
    wire N__37330;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37315;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37300;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37285;
    wire N__37284;
    wire N__37281;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37258;
    wire N__37255;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37228;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37188;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37164;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37141;
    wire N__37138;
    wire N__37135;
    wire N__37134;
    wire N__37131;
    wire N__37130;
    wire N__37127;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37109;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37095;
    wire N__37092;
    wire N__37087;
    wire N__37084;
    wire N__37083;
    wire N__37080;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37047;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36978;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36955;
    wire N__36952;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36922;
    wire N__36919;
    wire N__36918;
    wire N__36915;
    wire N__36914;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36891;
    wire N__36888;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36846;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36834;
    wire N__36833;
    wire N__36830;
    wire N__36825;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36798;
    wire N__36795;
    wire N__36794;
    wire N__36791;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36777;
    wire N__36774;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36727;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36696;
    wire N__36695;
    wire N__36694;
    wire N__36693;
    wire N__36692;
    wire N__36675;
    wire N__36672;
    wire N__36671;
    wire N__36670;
    wire N__36669;
    wire N__36668;
    wire N__36667;
    wire N__36666;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36644;
    wire N__36641;
    wire N__36634;
    wire N__36631;
    wire N__36630;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36591;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36565;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36553;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36501;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36486;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36436;
    wire N__36433;
    wire N__36430;
    wire N__36425;
    wire N__36420;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36342;
    wire N__36341;
    wire N__36338;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36294;
    wire N__36289;
    wire N__36286;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36201;
    wire N__36200;
    wire N__36195;
    wire N__36192;
    wire N__36187;
    wire N__36184;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36172;
    wire N__36169;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36094;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36067;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36057;
    wire N__36056;
    wire N__36053;
    wire N__36048;
    wire N__36043;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36033;
    wire N__36030;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36013;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36009;
    wire N__36008;
    wire N__36007;
    wire N__36006;
    wire N__36005;
    wire N__36004;
    wire N__36003;
    wire N__36002;
    wire N__36001;
    wire N__36000;
    wire N__35999;
    wire N__35998;
    wire N__35997;
    wire N__35994;
    wire N__35993;
    wire N__35992;
    wire N__35991;
    wire N__35990;
    wire N__35989;
    wire N__35988;
    wire N__35977;
    wire N__35966;
    wire N__35965;
    wire N__35964;
    wire N__35963;
    wire N__35962;
    wire N__35959;
    wire N__35958;
    wire N__35947;
    wire N__35946;
    wire N__35943;
    wire N__35938;
    wire N__35933;
    wire N__35930;
    wire N__35929;
    wire N__35928;
    wire N__35927;
    wire N__35926;
    wire N__35925;
    wire N__35924;
    wire N__35923;
    wire N__35922;
    wire N__35921;
    wire N__35918;
    wire N__35917;
    wire N__35916;
    wire N__35915;
    wire N__35914;
    wire N__35913;
    wire N__35912;
    wire N__35911;
    wire N__35910;
    wire N__35909;
    wire N__35904;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35896;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35868;
    wire N__35867;
    wire N__35866;
    wire N__35865;
    wire N__35860;
    wire N__35855;
    wire N__35854;
    wire N__35851;
    wire N__35846;
    wire N__35843;
    wire N__35838;
    wire N__35835;
    wire N__35826;
    wire N__35819;
    wire N__35814;
    wire N__35809;
    wire N__35802;
    wire N__35799;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35779;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35775;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35763;
    wire N__35758;
    wire N__35755;
    wire N__35748;
    wire N__35745;
    wire N__35740;
    wire N__35737;
    wire N__35730;
    wire N__35727;
    wire N__35724;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35714;
    wire N__35713;
    wire N__35712;
    wire N__35711;
    wire N__35710;
    wire N__35709;
    wire N__35702;
    wire N__35697;
    wire N__35692;
    wire N__35687;
    wire N__35670;
    wire N__35667;
    wire N__35662;
    wire N__35653;
    wire N__35648;
    wire N__35629;
    wire N__35626;
    wire N__35625;
    wire N__35624;
    wire N__35623;
    wire N__35618;
    wire N__35617;
    wire N__35616;
    wire N__35611;
    wire N__35610;
    wire N__35609;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35601;
    wire N__35600;
    wire N__35599;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35591;
    wire N__35588;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35572;
    wire N__35571;
    wire N__35568;
    wire N__35567;
    wire N__35566;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35552;
    wire N__35547;
    wire N__35542;
    wire N__35539;
    wire N__35534;
    wire N__35531;
    wire N__35526;
    wire N__35523;
    wire N__35520;
    wire N__35517;
    wire N__35512;
    wire N__35507;
    wire N__35504;
    wire N__35499;
    wire N__35494;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35472;
    wire N__35467;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35448;
    wire N__35447;
    wire N__35444;
    wire N__35439;
    wire N__35434;
    wire N__35433;
    wire N__35430;
    wire N__35425;
    wire N__35422;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35410;
    wire N__35409;
    wire N__35406;
    wire N__35405;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35388;
    wire N__35385;
    wire N__35382;
    wire N__35379;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35355;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35326;
    wire N__35323;
    wire N__35318;
    wire N__35311;
    wire N__35308;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35275;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35155;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35131;
    wire N__35130;
    wire N__35129;
    wire N__35128;
    wire N__35125;
    wire N__35118;
    wire N__35117;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35101;
    wire N__35098;
    wire N__35097;
    wire N__35096;
    wire N__35091;
    wire N__35088;
    wire N__35083;
    wire N__35082;
    wire N__35081;
    wire N__35080;
    wire N__35073;
    wire N__35070;
    wire N__35065;
    wire N__35064;
    wire N__35063;
    wire N__35062;
    wire N__35061;
    wire N__35052;
    wire N__35049;
    wire N__35044;
    wire N__35043;
    wire N__35042;
    wire N__35039;
    wire N__35038;
    wire N__35035;
    wire N__35034;
    wire N__35031;
    wire N__35030;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35022;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35014;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35006;
    wire N__35003;
    wire N__35002;
    wire N__35001;
    wire N__35000;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34984;
    wire N__34981;
    wire N__34980;
    wire N__34977;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34956;
    wire N__34953;
    wire N__34948;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34932;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34909;
    wire N__34902;
    wire N__34895;
    wire N__34892;
    wire N__34887;
    wire N__34886;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34792;
    wire N__34791;
    wire N__34788;
    wire N__34787;
    wire N__34786;
    wire N__34785;
    wire N__34784;
    wire N__34783;
    wire N__34782;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34751;
    wire N__34744;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34723;
    wire N__34718;
    wire N__34705;
    wire N__34702;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34697;
    wire N__34696;
    wire N__34695;
    wire N__34692;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34678;
    wire N__34673;
    wire N__34672;
    wire N__34671;
    wire N__34670;
    wire N__34667;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34655;
    wire N__34648;
    wire N__34645;
    wire N__34640;
    wire N__34633;
    wire N__34618;
    wire N__34615;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34548;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34536;
    wire N__34535;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34524;
    wire N__34523;
    wire N__34522;
    wire N__34519;
    wire N__34518;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34504;
    wire N__34503;
    wire N__34500;
    wire N__34499;
    wire N__34498;
    wire N__34495;
    wire N__34492;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34465;
    wire N__34458;
    wire N__34451;
    wire N__34448;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34386;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34344;
    wire N__34343;
    wire N__34340;
    wire N__34335;
    wire N__34332;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34300;
    wire N__34299;
    wire N__34294;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34276;
    wire N__34275;
    wire N__34274;
    wire N__34271;
    wire N__34266;
    wire N__34261;
    wire N__34258;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34246;
    wire N__34245;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34179;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34169;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34136;
    wire N__34133;
    wire N__34128;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34077;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34051;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34024;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34002;
    wire N__34001;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33993;
    wire N__33992;
    wire N__33991;
    wire N__33990;
    wire N__33989;
    wire N__33988;
    wire N__33987;
    wire N__33986;
    wire N__33985;
    wire N__33982;
    wire N__33981;
    wire N__33980;
    wire N__33979;
    wire N__33978;
    wire N__33975;
    wire N__33974;
    wire N__33973;
    wire N__33972;
    wire N__33967;
    wire N__33962;
    wire N__33955;
    wire N__33954;
    wire N__33953;
    wire N__33952;
    wire N__33951;
    wire N__33950;
    wire N__33945;
    wire N__33940;
    wire N__33939;
    wire N__33938;
    wire N__33937;
    wire N__33936;
    wire N__33935;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33921;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33903;
    wire N__33902;
    wire N__33897;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33868;
    wire N__33861;
    wire N__33858;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33836;
    wire N__33823;
    wire N__33820;
    wire N__33815;
    wire N__33812;
    wire N__33805;
    wire N__33804;
    wire N__33801;
    wire N__33798;
    wire N__33797;
    wire N__33794;
    wire N__33789;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33690;
    wire N__33689;
    wire N__33686;
    wire N__33681;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33669;
    wire N__33668;
    wire N__33665;
    wire N__33660;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33645;
    wire N__33644;
    wire N__33641;
    wire N__33636;
    wire N__33631;
    wire N__33628;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33610;
    wire N__33607;
    wire N__33606;
    wire N__33603;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33586;
    wire N__33583;
    wire N__33582;
    wire N__33581;
    wire N__33580;
    wire N__33579;
    wire N__33578;
    wire N__33577;
    wire N__33576;
    wire N__33575;
    wire N__33574;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33556;
    wire N__33553;
    wire N__33552;
    wire N__33551;
    wire N__33550;
    wire N__33549;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33537;
    wire N__33536;
    wire N__33535;
    wire N__33534;
    wire N__33533;
    wire N__33532;
    wire N__33531;
    wire N__33526;
    wire N__33517;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33494;
    wire N__33485;
    wire N__33480;
    wire N__33475;
    wire N__33472;
    wire N__33467;
    wire N__33448;
    wire N__33447;
    wire N__33446;
    wire N__33445;
    wire N__33444;
    wire N__33443;
    wire N__33442;
    wire N__33441;
    wire N__33440;
    wire N__33439;
    wire N__33438;
    wire N__33437;
    wire N__33436;
    wire N__33433;
    wire N__33432;
    wire N__33431;
    wire N__33430;
    wire N__33429;
    wire N__33426;
    wire N__33411;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33403;
    wire N__33402;
    wire N__33399;
    wire N__33398;
    wire N__33397;
    wire N__33396;
    wire N__33395;
    wire N__33394;
    wire N__33393;
    wire N__33388;
    wire N__33387;
    wire N__33386;
    wire N__33385;
    wire N__33382;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33368;
    wire N__33363;
    wire N__33356;
    wire N__33355;
    wire N__33354;
    wire N__33353;
    wire N__33352;
    wire N__33349;
    wire N__33348;
    wire N__33333;
    wire N__33330;
    wire N__33327;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33315;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33303;
    wire N__33300;
    wire N__33295;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33285;
    wire N__33274;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33266;
    wire N__33261;
    wire N__33258;
    wire N__33253;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33233;
    wire N__33226;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33182;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33150;
    wire N__33147;
    wire N__33146;
    wire N__33145;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33130;
    wire N__33121;
    wire N__33118;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33096;
    wire N__33091;
    wire N__33088;
    wire N__33087;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33066;
    wire N__33063;
    wire N__33056;
    wire N__33053;
    wire N__33046;
    wire N__33043;
    wire N__33042;
    wire N__33041;
    wire N__33040;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33013;
    wire N__33010;
    wire N__33009;
    wire N__33008;
    wire N__33007;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32992;
    wire N__32989;
    wire N__32980;
    wire N__32977;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32965;
    wire N__32962;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32904;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32887;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32874;
    wire N__32873;
    wire N__32872;
    wire N__32869;
    wire N__32862;
    wire N__32857;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32845;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32833;
    wire N__32830;
    wire N__32829;
    wire N__32828;
    wire N__32825;
    wire N__32820;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32804;
    wire N__32801;
    wire N__32800;
    wire N__32795;
    wire N__32792;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32734;
    wire N__32733;
    wire N__32732;
    wire N__32731;
    wire N__32730;
    wire N__32729;
    wire N__32728;
    wire N__32727;
    wire N__32726;
    wire N__32725;
    wire N__32724;
    wire N__32723;
    wire N__32722;
    wire N__32719;
    wire N__32716;
    wire N__32715;
    wire N__32714;
    wire N__32713;
    wire N__32712;
    wire N__32711;
    wire N__32710;
    wire N__32709;
    wire N__32708;
    wire N__32707;
    wire N__32704;
    wire N__32703;
    wire N__32702;
    wire N__32701;
    wire N__32700;
    wire N__32697;
    wire N__32696;
    wire N__32689;
    wire N__32688;
    wire N__32679;
    wire N__32674;
    wire N__32665;
    wire N__32650;
    wire N__32647;
    wire N__32642;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32622;
    wire N__32621;
    wire N__32620;
    wire N__32619;
    wire N__32618;
    wire N__32617;
    wire N__32608;
    wire N__32607;
    wire N__32606;
    wire N__32605;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32597;
    wire N__32596;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32577;
    wire N__32564;
    wire N__32561;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32543;
    wire N__32536;
    wire N__32531;
    wire N__32528;
    wire N__32509;
    wire N__32508;
    wire N__32507;
    wire N__32506;
    wire N__32505;
    wire N__32498;
    wire N__32497;
    wire N__32496;
    wire N__32495;
    wire N__32494;
    wire N__32491;
    wire N__32490;
    wire N__32487;
    wire N__32486;
    wire N__32485;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32473;
    wire N__32472;
    wire N__32471;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32428;
    wire N__32421;
    wire N__32414;
    wire N__32411;
    wire N__32406;
    wire N__32403;
    wire N__32380;
    wire N__32377;
    wire N__32376;
    wire N__32373;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32313;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32283;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32235;
    wire N__32232;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32196;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32149;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32143;
    wire N__32142;
    wire N__32137;
    wire N__32132;
    wire N__32129;
    wire N__32122;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32114;
    wire N__32109;
    wire N__32106;
    wire N__32101;
    wire N__32100;
    wire N__32099;
    wire N__32096;
    wire N__32095;
    wire N__32094;
    wire N__32093;
    wire N__32092;
    wire N__32091;
    wire N__32090;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32073;
    wire N__32072;
    wire N__32071;
    wire N__32068;
    wire N__32067;
    wire N__32066;
    wire N__32061;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32039;
    wire N__32034;
    wire N__32029;
    wire N__32020;
    wire N__32011;
    wire N__32008;
    wire N__32005;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31993;
    wire N__31992;
    wire N__31991;
    wire N__31988;
    wire N__31981;
    wire N__31976;
    wire N__31973;
    wire N__31972;
    wire N__31971;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31963;
    wire N__31958;
    wire N__31953;
    wire N__31948;
    wire N__31945;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31918;
    wire N__31915;
    wire N__31914;
    wire N__31913;
    wire N__31912;
    wire N__31911;
    wire N__31906;
    wire N__31901;
    wire N__31898;
    wire N__31891;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31877;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31854;
    wire N__31853;
    wire N__31850;
    wire N__31845;
    wire N__31840;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31830;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31762;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31716;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31644;
    wire N__31643;
    wire N__31640;
    wire N__31635;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31595;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31551;
    wire N__31548;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31516;
    wire N__31513;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31485;
    wire N__31484;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31432;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31417;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31405;
    wire N__31402;
    wire N__31399;
    wire N__31396;
    wire N__31393;
    wire N__31390;
    wire N__31389;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31377;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31365;
    wire N__31360;
    wire N__31357;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31339;
    wire N__31336;
    wire N__31335;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31323;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31252;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31197;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31182;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31170;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31159;
    wire N__31158;
    wire N__31153;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31126;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31114;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31084;
    wire N__31083;
    wire N__31082;
    wire N__31081;
    wire N__31080;
    wire N__31079;
    wire N__31078;
    wire N__31077;
    wire N__31076;
    wire N__31075;
    wire N__31074;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31068;
    wire N__31067;
    wire N__31066;
    wire N__31065;
    wire N__31064;
    wire N__31063;
    wire N__31062;
    wire N__31061;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31037;
    wire N__31034;
    wire N__31033;
    wire N__31032;
    wire N__31017;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30982;
    wire N__30977;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30946;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30795;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30768;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30639;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30604;
    wire N__30603;
    wire N__30600;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30564;
    wire N__30561;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30510;
    wire N__30507;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30497;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30456;
    wire N__30453;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30436;
    wire N__30435;
    wire N__30434;
    wire N__30433;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30425;
    wire N__30424;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30411;
    wire N__30410;
    wire N__30405;
    wire N__30402;
    wire N__30395;
    wire N__30382;
    wire N__30373;
    wire N__30372;
    wire N__30371;
    wire N__30368;
    wire N__30367;
    wire N__30366;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30346;
    wire N__30345;
    wire N__30344;
    wire N__30343;
    wire N__30342;
    wire N__30341;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30315;
    wire N__30304;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30271;
    wire N__30268;
    wire N__30267;
    wire N__30264;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30147;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30039;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29850;
    wire N__29847;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29734;
    wire N__29733;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29184;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29097;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29067;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29010;
    wire N__29009;
    wire N__29008;
    wire N__29005;
    wire N__28998;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28966;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28954;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28942;
    wire N__28941;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28924;
    wire N__28923;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28901;
    wire N__28900;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28884;
    wire N__28879;
    wire N__28876;
    wire N__28875;
    wire N__28872;
    wire N__28869;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28789;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28769;
    wire N__28764;
    wire N__28761;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28723;
    wire N__28722;
    wire N__28719;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28696;
    wire N__28693;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28675;
    wire N__28672;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28642;
    wire N__28639;
    wire N__28638;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28626;
    wire N__28625;
    wire N__28622;
    wire N__28621;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28593;
    wire N__28590;
    wire N__28589;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28564;
    wire N__28563;
    wire N__28562;
    wire N__28561;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28553;
    wire N__28550;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28497;
    wire N__28492;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28467;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28426;
    wire N__28425;
    wire N__28422;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28402;
    wire N__28401;
    wire N__28398;
    wire N__28397;
    wire N__28396;
    wire N__28395;
    wire N__28394;
    wire N__28393;
    wire N__28392;
    wire N__28391;
    wire N__28390;
    wire N__28387;
    wire N__28386;
    wire N__28385;
    wire N__28382;
    wire N__28381;
    wire N__28380;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28372;
    wire N__28371;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28348;
    wire N__28345;
    wire N__28344;
    wire N__28343;
    wire N__28342;
    wire N__28339;
    wire N__28338;
    wire N__28337;
    wire N__28328;
    wire N__28315;
    wire N__28310;
    wire N__28297;
    wire N__28292;
    wire N__28285;
    wire N__28282;
    wire N__28281;
    wire N__28278;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28258;
    wire N__28255;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28243;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28231;
    wire N__28228;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28195;
    wire N__28192;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28180;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28122;
    wire N__28121;
    wire N__28118;
    wire N__28113;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28089;
    wire N__28088;
    wire N__28085;
    wire N__28080;
    wire N__28075;
    wire N__28074;
    wire N__28073;
    wire N__28070;
    wire N__28065;
    wire N__28060;
    wire N__28059;
    wire N__28056;
    wire N__28055;
    wire N__28048;
    wire N__28045;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28033;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28021;
    wire N__28018;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27993;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27970;
    wire N__27969;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27927;
    wire N__27926;
    wire N__27923;
    wire N__27918;
    wire N__27913;
    wire N__27910;
    wire N__27909;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27889;
    wire N__27886;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27854;
    wire N__27851;
    wire N__27846;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27828;
    wire N__27825;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27706;
    wire N__27703;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27691;
    wire N__27688;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27676;
    wire N__27673;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27636;
    wire N__27635;
    wire N__27632;
    wire N__27627;
    wire N__27624;
    wire N__27619;
    wire N__27616;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27604;
    wire N__27601;
    wire N__27600;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27577;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27523;
    wire N__27520;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27501;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27475;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27463;
    wire N__27460;
    wire N__27459;
    wire N__27458;
    wire N__27455;
    wire N__27450;
    wire N__27447;
    wire N__27442;
    wire N__27439;
    wire N__27438;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27415;
    wire N__27412;
    wire N__27411;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27379;
    wire N__27376;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27364;
    wire N__27361;
    wire N__27360;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27340;
    wire N__27337;
    wire N__27336;
    wire N__27333;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27313;
    wire N__27310;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27298;
    wire N__27295;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27285;
    wire N__27282;
    wire N__27277;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27265;
    wire N__27262;
    wire N__27261;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27238;
    wire N__27235;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27223;
    wire N__27220;
    wire N__27219;
    wire N__27218;
    wire N__27215;
    wire N__27210;
    wire N__27207;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27192;
    wire N__27189;
    wire N__27188;
    wire N__27185;
    wire N__27180;
    wire N__27177;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27159;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27129;
    wire N__27128;
    wire N__27125;
    wire N__27120;
    wire N__27117;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27084;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27054;
    wire N__27053;
    wire N__27050;
    wire N__27045;
    wire N__27042;
    wire N__27037;
    wire N__27034;
    wire N__27033;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27006;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26991;
    wire N__26988;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26970;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26940;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26925;
    wire N__26922;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26866;
    wire N__26865;
    wire N__26864;
    wire N__26863;
    wire N__26862;
    wire N__26859;
    wire N__26858;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26853;
    wire N__26852;
    wire N__26849;
    wire N__26848;
    wire N__26847;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26839;
    wire N__26838;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26823;
    wire N__26822;
    wire N__26819;
    wire N__26818;
    wire N__26817;
    wire N__26814;
    wire N__26805;
    wire N__26800;
    wire N__26799;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26787;
    wire N__26786;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26772;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26738;
    wire N__26733;
    wire N__26726;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26710;
    wire N__26701;
    wire N__26680;
    wire N__26677;
    wire N__26676;
    wire N__26675;
    wire N__26674;
    wire N__26673;
    wire N__26672;
    wire N__26671;
    wire N__26670;
    wire N__26669;
    wire N__26668;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26654;
    wire N__26653;
    wire N__26652;
    wire N__26651;
    wire N__26650;
    wire N__26647;
    wire N__26646;
    wire N__26643;
    wire N__26632;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26618;
    wire N__26617;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26609;
    wire N__26608;
    wire N__26607;
    wire N__26606;
    wire N__26605;
    wire N__26604;
    wire N__26599;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26581;
    wire N__26574;
    wire N__26569;
    wire N__26566;
    wire N__26561;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26536;
    wire N__26521;
    wire N__26520;
    wire N__26519;
    wire N__26518;
    wire N__26517;
    wire N__26516;
    wire N__26515;
    wire N__26514;
    wire N__26511;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26503;
    wire N__26502;
    wire N__26501;
    wire N__26500;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26496;
    wire N__26495;
    wire N__26494;
    wire N__26493;
    wire N__26492;
    wire N__26491;
    wire N__26490;
    wire N__26487;
    wire N__26486;
    wire N__26483;
    wire N__26476;
    wire N__26475;
    wire N__26474;
    wire N__26473;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26459;
    wire N__26456;
    wire N__26441;
    wire N__26438;
    wire N__26437;
    wire N__26436;
    wire N__26435;
    wire N__26434;
    wire N__26433;
    wire N__26432;
    wire N__26431;
    wire N__26430;
    wire N__26425;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26399;
    wire N__26398;
    wire N__26395;
    wire N__26394;
    wire N__26393;
    wire N__26392;
    wire N__26389;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26375;
    wire N__26374;
    wire N__26373;
    wire N__26372;
    wire N__26367;
    wire N__26356;
    wire N__26349;
    wire N__26340;
    wire N__26337;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26318;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26298;
    wire N__26291;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26252;
    wire N__26251;
    wire N__26250;
    wire N__26249;
    wire N__26248;
    wire N__26239;
    wire N__26236;
    wire N__26235;
    wire N__26234;
    wire N__26233;
    wire N__26230;
    wire N__26229;
    wire N__26226;
    wire N__26225;
    wire N__26224;
    wire N__26223;
    wire N__26222;
    wire N__26217;
    wire N__26214;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26191;
    wire N__26190;
    wire N__26189;
    wire N__26188;
    wire N__26187;
    wire N__26186;
    wire N__26185;
    wire N__26182;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26174;
    wire N__26169;
    wire N__26166;
    wire N__26165;
    wire N__26160;
    wire N__26157;
    wire N__26152;
    wire N__26147;
    wire N__26146;
    wire N__26145;
    wire N__26144;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26092;
    wire N__26089;
    wire N__26082;
    wire N__26077;
    wire N__26072;
    wire N__26069;
    wire N__26060;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25972;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25954;
    wire N__25951;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25939;
    wire N__25936;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25906;
    wire N__25903;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25875;
    wire N__25870;
    wire N__25869;
    wire N__25868;
    wire N__25867;
    wire N__25864;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25818;
    wire N__25817;
    wire N__25816;
    wire N__25813;
    wire N__25812;
    wire N__25807;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25782;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25753;
    wire N__25752;
    wire N__25747;
    wire N__25744;
    wire N__25743;
    wire N__25738;
    wire N__25735;
    wire N__25734;
    wire N__25731;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25708;
    wire N__25705;
    wire N__25704;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25636;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25624;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25609;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25597;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25585;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25573;
    wire N__25570;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25558;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25446;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25428;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25389;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25377;
    wire N__25372;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25360;
    wire N__25357;
    wire N__25356;
    wire N__25351;
    wire N__25348;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25225;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25217;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25198;
    wire N__25197;
    wire N__25196;
    wire N__25193;
    wire N__25188;
    wire N__25183;
    wire N__25180;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25162;
    wire N__25159;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25141;
    wire N__25138;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25108;
    wire N__25105;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25077;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25059;
    wire N__25056;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25027;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24961;
    wire N__24958;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24933;
    wire N__24930;
    wire N__24929;
    wire N__24928;
    wire N__24925;
    wire N__24924;
    wire N__24923;
    wire N__24922;
    wire N__24919;
    wire N__24914;
    wire N__24905;
    wire N__24902;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24762;
    wire N__24761;
    wire N__24760;
    wire N__24759;
    wire N__24758;
    wire N__24757;
    wire N__24756;
    wire N__24755;
    wire N__24754;
    wire N__24753;
    wire N__24752;
    wire N__24751;
    wire N__24750;
    wire N__24749;
    wire N__24748;
    wire N__24731;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24707;
    wire N__24706;
    wire N__24705;
    wire N__24704;
    wire N__24703;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24691;
    wire N__24690;
    wire N__24689;
    wire N__24688;
    wire N__24685;
    wire N__24684;
    wire N__24679;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24656;
    wire N__24647;
    wire N__24640;
    wire N__24639;
    wire N__24636;
    wire N__24635;
    wire N__24634;
    wire N__24633;
    wire N__24632;
    wire N__24631;
    wire N__24630;
    wire N__24629;
    wire N__24628;
    wire N__24627;
    wire N__24626;
    wire N__24625;
    wire N__24624;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24620;
    wire N__24619;
    wire N__24618;
    wire N__24615;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24611;
    wire N__24610;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24588;
    wire N__24585;
    wire N__24568;
    wire N__24565;
    wire N__24560;
    wire N__24557;
    wire N__24550;
    wire N__24547;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24530;
    wire N__24523;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24496;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24343;
    wire N__24340;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24322;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24262;
    wire N__24259;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24232;
    wire N__24229;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24204;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24192;
    wire N__24189;
    wire N__24186;
    wire N__24181;
    wire N__24180;
    wire N__24177;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24156;
    wire N__24155;
    wire N__24154;
    wire N__24151;
    wire N__24138;
    wire N__24133;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24118;
    wire N__24115;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24091;
    wire N__24090;
    wire N__24089;
    wire N__24088;
    wire N__24087;
    wire N__24084;
    wire N__24083;
    wire N__24080;
    wire N__24079;
    wire N__24078;
    wire N__24077;
    wire N__24076;
    wire N__24073;
    wire N__24068;
    wire N__24067;
    wire N__24062;
    wire N__24055;
    wire N__24054;
    wire N__24053;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24041;
    wire N__24038;
    wire N__24037;
    wire N__24032;
    wire N__24027;
    wire N__24024;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__23999;
    wire N__23986;
    wire N__23985;
    wire N__23984;
    wire N__23983;
    wire N__23982;
    wire N__23981;
    wire N__23980;
    wire N__23979;
    wire N__23978;
    wire N__23977;
    wire N__23976;
    wire N__23975;
    wire N__23974;
    wire N__23967;
    wire N__23960;
    wire N__23955;
    wire N__23950;
    wire N__23945;
    wire N__23942;
    wire N__23941;
    wire N__23940;
    wire N__23939;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23915;
    wire N__23912;
    wire N__23907;
    wire N__23902;
    wire N__23893;
    wire N__23892;
    wire N__23891;
    wire N__23888;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23835;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23823;
    wire N__23818;
    wire N__23817;
    wire N__23816;
    wire N__23815;
    wire N__23814;
    wire N__23813;
    wire N__23812;
    wire N__23811;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23792;
    wire N__23789;
    wire N__23784;
    wire N__23783;
    wire N__23782;
    wire N__23781;
    wire N__23780;
    wire N__23779;
    wire N__23772;
    wire N__23769;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23749;
    wire N__23746;
    wire N__23741;
    wire N__23736;
    wire N__23733;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23715;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23689;
    wire N__23688;
    wire N__23687;
    wire N__23686;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23650;
    wire N__23649;
    wire N__23648;
    wire N__23645;
    wire N__23640;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23584;
    wire N__23583;
    wire N__23578;
    wire N__23575;
    wire N__23574;
    wire N__23571;
    wire N__23566;
    wire N__23563;
    wire N__23562;
    wire N__23557;
    wire N__23554;
    wire N__23553;
    wire N__23548;
    wire N__23545;
    wire N__23544;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23502;
    wire N__23499;
    wire N__23492;
    wire N__23483;
    wire N__23476;
    wire N__23475;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23463;
    wire N__23462;
    wire N__23461;
    wire N__23460;
    wire N__23459;
    wire N__23458;
    wire N__23455;
    wire N__23446;
    wire N__23443;
    wire N__23436;
    wire N__23433;
    wire N__23428;
    wire N__23425;
    wire N__23416;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23404;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23364;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23349;
    wire N__23346;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23292;
    wire N__23291;
    wire N__23288;
    wire N__23283;
    wire N__23278;
    wire N__23275;
    wire N__23272;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23161;
    wire N__23160;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23138;
    wire N__23135;
    wire N__23130;
    wire N__23125;
    wire N__23124;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23091;
    wire N__23088;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23052;
    wire N__23049;
    wire N__23044;
    wire N__23041;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23022;
    wire N__23021;
    wire N__23018;
    wire N__23013;
    wire N__23008;
    wire N__23005;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22968;
    wire N__22967;
    wire N__22964;
    wire N__22959;
    wire N__22954;
    wire N__22951;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22943;
    wire N__22940;
    wire N__22935;
    wire N__22930;
    wire N__22927;
    wire N__22926;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22896;
    wire N__22895;
    wire N__22892;
    wire N__22887;
    wire N__22882;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22687;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22670;
    wire N__22665;
    wire N__22662;
    wire N__22657;
    wire N__22654;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22638;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22590;
    wire N__22585;
    wire N__22582;
    wire N__22581;
    wire N__22576;
    wire N__22573;
    wire N__22572;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22554;
    wire N__22549;
    wire N__22546;
    wire N__22545;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22526;
    wire N__22521;
    wire N__22516;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22508;
    wire N__22503;
    wire N__22500;
    wire N__22495;
    wire N__22492;
    wire N__22491;
    wire N__22486;
    wire N__22483;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22471;
    wire N__22468;
    wire N__22467;
    wire N__22464;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22452;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22375;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22363;
    wire N__22360;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22348;
    wire N__22345;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22311;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22296;
    wire N__22295;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22283;
    wire N__22280;
    wire N__22275;
    wire N__22272;
    wire N__22267;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22189;
    wire N__22186;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22178;
    wire N__22175;
    wire N__22170;
    wire N__22165;
    wire N__22162;
    wire N__22161;
    wire N__22158;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22120;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22108;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22093;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22062;
    wire N__22061;
    wire N__22058;
    wire N__22053;
    wire N__22048;
    wire N__22045;
    wire N__22044;
    wire N__22041;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22024;
    wire N__22021;
    wire N__22020;
    wire N__22019;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21984;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21961;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21953;
    wire N__21948;
    wire N__21943;
    wire N__21942;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21916;
    wire N__21915;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21886;
    wire N__21885;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21873;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21861;
    wire N__21858;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21841;
    wire N__21838;
    wire N__21837;
    wire N__21836;
    wire N__21833;
    wire N__21828;
    wire N__21823;
    wire N__21822;
    wire N__21819;
    wire N__21818;
    wire N__21815;
    wire N__21810;
    wire N__21807;
    wire N__21802;
    wire N__21799;
    wire N__21798;
    wire N__21797;
    wire N__21796;
    wire N__21793;
    wire N__21786;
    wire N__21783;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21774;
    wire N__21769;
    wire N__21768;
    wire N__21767;
    wire N__21764;
    wire N__21763;
    wire N__21758;
    wire N__21755;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21736;
    wire N__21733;
    wire N__21728;
    wire N__21725;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21705;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21687;
    wire N__21682;
    wire N__21681;
    wire N__21678;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21666;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21633;
    wire N__21630;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21546;
    wire N__21541;
    wire N__21538;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21512;
    wire N__21509;
    wire N__21504;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21453;
    wire N__21452;
    wire N__21451;
    wire N__21450;
    wire N__21447;
    wire N__21440;
    wire N__21437;
    wire N__21430;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21390;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire ICE_GPMO_2;
    wire VCCG0;
    wire INViac_raw_buf_vac_raw_buf_merged11WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged3WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged10WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged8WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged4WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged9WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged5WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged0WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged6WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged1WCLKN_net;
    wire ICE_SYSCLK;
    wire INViac_raw_buf_vac_raw_buf_merged7WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged2WCLKN_net;
    wire RTD_SCLK;
    wire \RTD.n8 ;
    wire RTD_SDI;
    wire \RTD.n21253 ;
    wire VAC_MISO;
    wire cmd_rdadctmp_0_adj_1548;
    wire VAC_SCLK;
    wire n14_cascade_;
    wire n21889;
    wire VAC_CS;
    wire DDS_SCK1;
    wire \RTD.n12262 ;
    wire RTD_SDO;
    wire \CLK_DDS.n18366 ;
    wire bit_cnt_0_adj_1512;
    wire bit_cnt_3;
    wire n22326;
    wire \CLK_DDS.n9 ;
    wire buf_adcdata_vac_4;
    wire cmd_rdadctmp_1_adj_1547;
    wire cmd_rdadctmp_14_adj_1534;
    wire bfn_2_14_0_;
    wire \ADC_VAC.n20683 ;
    wire \ADC_VAC.n20684 ;
    wire \ADC_VAC.n20685 ;
    wire \ADC_VAC.n20686 ;
    wire \ADC_VAC.n20687 ;
    wire \ADC_VAC.n20688 ;
    wire \ADC_VAC.n20689 ;
    wire \ADC_VAC.n13784 ;
    wire \ADC_VAC.n13784_cascade_ ;
    wire \ADC_VAC.n15660 ;
    wire \RTD.n22632_cascade_ ;
    wire DDS_CS1;
    wire \CLK_DDS.n9_adj_1489 ;
    wire read_buf_15;
    wire read_buf_10;
    wire bit_cnt_2;
    wire bit_cnt_1;
    wire dds_state_0_adj_1510;
    wire n8_adj_1686;
    wire read_buf_11;
    wire read_buf_12;
    wire read_buf_14;
    wire read_buf_3;
    wire read_buf_13;
    wire n19_adj_1690_cascade_;
    wire buf_adcdata_vac_6;
    wire n19_adj_1693_cascade_;
    wire buf_data_iac_5;
    wire buf_adcdata_iac_6;
    wire buf_adcdata_iac_7;
    wire cmd_rdadctmp_14;
    wire n19_adj_1700;
    wire buf_data_iac_4;
    wire n22_adj_1701_cascade_;
    wire buf_adcdata_vac_7;
    wire buf_adcdata_iac_4;
    wire n22_adj_1697;
    wire cmd_rdadctmp_15_adj_1533;
    wire cmd_rdadctmp_13;
    wire buf_adcdata_iac_5;
    wire \ADC_VAC.n13747_cascade_ ;
    wire \ADC_VAC.n13842 ;
    wire \ADC_VAC.bit_cnt_2 ;
    wire \ADC_VAC.bit_cnt_1 ;
    wire \ADC_VAC.bit_cnt_3 ;
    wire \ADC_VAC.bit_cnt_4 ;
    wire \ADC_VAC.bit_cnt_6 ;
    wire \ADC_VAC.bit_cnt_0 ;
    wire \ADC_VAC.n22109_cascade_ ;
    wire \ADC_VAC.bit_cnt_7 ;
    wire \ADC_VAC.n22126_cascade_ ;
    wire \ADC_VAC.bit_cnt_5 ;
    wire \ADC_VAC.n22389_cascade_ ;
    wire \ADC_VAC.n22030 ;
    wire \ADC_VAC.n17 ;
    wire VAC_DRDY;
    wire \ADC_VAC.n12 ;
    wire RTD_CS;
    wire \RTD.n22382 ;
    wire \RTD.n20051_cascade_ ;
    wire \RTD.n22079 ;
    wire \RTD.n22599_cascade_ ;
    wire \RTD.n23689 ;
    wire \RTD.n56_cascade_ ;
    wire \RTD.n5 ;
    wire \RTD.n71 ;
    wire \RTD.n71_cascade_ ;
    wire \RTD.n22623 ;
    wire \RTD.n20051 ;
    wire read_buf_0;
    wire \RTD.read_buf_4 ;
    wire n21989_cascade_;
    wire read_buf_1;
    wire read_buf_2;
    wire \RTD.n68_cascade_ ;
    wire \RTD.cfg_buf_4 ;
    wire \RTD.cfg_buf_2 ;
    wire \RTD.cfg_buf_0 ;
    wire \RTD.n10 ;
    wire \RTD.n9_cascade_ ;
    wire \RTD.cfg_buf_3 ;
    wire \RTD.adress_7 ;
    wire \RTD.n19_cascade_ ;
    wire \RTD.n15396 ;
    wire \RTD.n1 ;
    wire \RTD.n1_cascade_ ;
    wire \RTD.cfg_tmp_0 ;
    wire \RTD.cfg_tmp_1 ;
    wire \RTD.cfg_tmp_2 ;
    wire \RTD.cfg_tmp_3 ;
    wire \RTD.cfg_tmp_4 ;
    wire \RTD.cfg_tmp_5 ;
    wire \RTD.cfg_tmp_6 ;
    wire \RTD.cfg_tmp_7 ;
    wire buf_data_iac_6;
    wire n22_adj_1694;
    wire buf_readRTD_1;
    wire cmd_rdadctmp_2_adj_1546;
    wire cmd_rdadctmp_12;
    wire n19_adj_1696;
    wire buf_data_iac_7;
    wire n22_adj_1691;
    wire cmd_rdadctmp_16_adj_1532;
    wire cmd_rdadctmp_23_adj_1525;
    wire cmd_rdadctmp_24_adj_1524;
    wire cmd_rdadctmp_28_adj_1520;
    wire cmd_rdadctmp_15;
    wire cmd_rdadctmp_13_adj_1535;
    wire buf_adcdata_vac_5;
    wire cmd_rdadctmp_17_adj_1531;
    wire cmd_rdadctmp_18_adj_1530;
    wire n23543_cascade_;
    wire cmd_rdadctmp_31_adj_1517;
    wire cmd_rdadctmp_29_adj_1519;
    wire cmd_rdadctmp_30_adj_1518;
    wire n21948_cascade_;
    wire buf_adcdata_vac_22;
    wire AC_ADC_SYNC;
    wire \RTD.n21988 ;
    wire \RTD.n7_adj_1497_cascade_ ;
    wire n13603_cascade_;
    wire read_buf_5;
    wire \RTD.n62 ;
    wire \RTD.n12274 ;
    wire \RTD.n11_adj_1500 ;
    wire buf_adcdata_vac_23;
    wire n23435;
    wire \RTD.mode ;
    wire \RTD.cfg_buf_6 ;
    wire \RTD.cfg_buf_5 ;
    wire \RTD.n12 ;
    wire \RTD.cfg_buf_1 ;
    wire \RTD.n20093 ;
    wire \RTD.n13482 ;
    wire \RTD.n68 ;
    wire \RTD.cfg_buf_7 ;
    wire buf_readRTD_14;
    wire \RTD.n68_adj_1498 ;
    wire \RTD.n21954 ;
    wire RTD_DRDY;
    wire \RTD.n21954_cascade_ ;
    wire \RTD.n21955 ;
    wire \RTD.adress_7_N_1009_7 ;
    wire \RTD.n11 ;
    wire \RTD.n11_cascade_ ;
    wire \RTD.n13488 ;
    wire \RTD.n13488_cascade_ ;
    wire \RTD.n15585 ;
    wire \RTD.n22081 ;
    wire \RTD.adress_6 ;
    wire \RTD.adress_5 ;
    wire \RTD.adress_4 ;
    wire \RTD.adress_3 ;
    wire \RTD.adress_2 ;
    wire \RTD.adress_0 ;
    wire \RTD.n13441 ;
    wire \RTD.adress_1 ;
    wire read_buf_6;
    wire n21989;
    wire n13584;
    wire read_buf_7;
    wire buf_adcdata_vac_9;
    wire n19_adj_1752;
    wire read_buf_8;
    wire n13603;
    wire read_buf_9;
    wire buf_readRTD_2;
    wire cmd_rdadctmp_12_adj_1536;
    wire DDS_MOSI1;
    wire cmd_rdadctmp_22_adj_1526;
    wire buf_adcdata_vac_15;
    wire n19_adj_1714_cascade_;
    wire buf_readRTD_7;
    wire \CLK_DDS.tmp_buf_10 ;
    wire \CLK_DDS.tmp_buf_11 ;
    wire \CLK_DDS.tmp_buf_12 ;
    wire \CLK_DDS.tmp_buf_13 ;
    wire \CLK_DDS.tmp_buf_14 ;
    wire \CLK_DDS.tmp_buf_9 ;
    wire \CLK_DDS.tmp_buf_8 ;
    wire tmp_buf_15_adj_1511;
    wire \CLK_DDS.tmp_buf_0 ;
    wire \CLK_DDS.tmp_buf_1 ;
    wire \CLK_DDS.tmp_buf_2 ;
    wire \CLK_DDS.tmp_buf_3 ;
    wire \CLK_DDS.tmp_buf_4 ;
    wire \CLK_DDS.tmp_buf_5 ;
    wire dds_state_2_adj_1508;
    wire dds_state_1_adj_1509;
    wire \CLK_DDS.tmp_buf_6 ;
    wire \CLK_DDS.tmp_buf_7 ;
    wire \CLK_DDS.n13376 ;
    wire n19_adj_1765;
    wire n20_adj_1766;
    wire n21892_cascade_;
    wire IAC_MISO;
    wire GB_BUFFER_DDS_MCLK1_THRU_CO;
    wire n22388;
    wire VDC_SCLK;
    wire n12356;
    wire \RTD.n17 ;
    wire \RTD.n79 ;
    wire buf_adcdata_vdc_15;
    wire buf_adcdata_vdc_7;
    wire buf_adcdata_vdc_23;
    wire buf_adcdata_vdc_4;
    wire buf_adcdata_vdc_9;
    wire buf_adcdata_vdc_6;
    wire buf_adcdata_vdc_22;
    wire cmd_rdadctmp_26_adj_1522;
    wire n112_adj_1786_cascade_;
    wire buf_adcdata_vdc_10;
    wire buf_adcdata_vac_10;
    wire n19_adj_1747;
    wire comm_test_buf_24_22;
    wire buf_dds1_15;
    wire n111_adj_1771;
    wire buf_adcdata_vdc_8;
    wire buf_adcdata_vac_8;
    wire n30_adj_1695;
    wire buf_readRTD_11;
    wire buf_cfgRTD_3;
    wire n20_adj_1790;
    wire n23498_cascade_;
    wire buf_adcdata_vdc_20;
    wire buf_adcdata_vac_20;
    wire n16_adj_1787;
    wire n17_adj_1788;
    wire n23540;
    wire buf_adcdata_iac_23;
    wire cmd_rdadctmp_31;
    wire n19;
    wire buf_readRTD_0;
    wire n22041_cascade_;
    wire INVacadc_trig_303C_net;
    wire bfn_7_16_0_;
    wire \ADC_IAC.n20676 ;
    wire \ADC_IAC.n20677 ;
    wire \ADC_IAC.n20678 ;
    wire \ADC_IAC.n20679 ;
    wire \ADC_IAC.n20680 ;
    wire \ADC_IAC.n20681 ;
    wire \ADC_IAC.n20682 ;
    wire \ADC_IAC.n13667 ;
    wire \ADC_IAC.n15622 ;
    wire \ADC_IAC.n22031 ;
    wire \ADC_IAC.bit_cnt_4 ;
    wire \ADC_IAC.bit_cnt_3 ;
    wire \ADC_IAC.bit_cnt_1 ;
    wire \ADC_IAC.bit_cnt_2 ;
    wire \ADC_IAC.bit_cnt_6 ;
    wire \ADC_IAC.bit_cnt_0 ;
    wire \ADC_IAC.n22113_cascade_ ;
    wire \ADC_IAC.bit_cnt_7 ;
    wire \ADC_IAC.bit_cnt_5 ;
    wire \ADC_IAC.n22128_cascade_ ;
    wire \ADC_IAC.n22384_cascade_ ;
    wire \ADC_IAC.n22032 ;
    wire acadc_trig;
    wire \ADC_IAC.n17_cascade_ ;
    wire \ADC_IAC.n12 ;
    wire n21892;
    wire n14_adj_1578;
    wire IAC_DRDY;
    wire IAC_CS;
    wire cmd_rdadctmp_2;
    wire cmd_rdadctmp_3;
    wire cmd_rdadctmp_4;
    wire cmd_rdadctmp_0;
    wire cmd_rdadctmp_1;
    wire EIS_SYNCCLK;
    wire IAC_CLK;
    wire bfn_8_2_0_;
    wire \ADC_VDC.avg_cnt_1 ;
    wire \ADC_VDC.n20725 ;
    wire \ADC_VDC.avg_cnt_2 ;
    wire \ADC_VDC.n20726 ;
    wire \ADC_VDC.avg_cnt_3 ;
    wire \ADC_VDC.n20727 ;
    wire \ADC_VDC.avg_cnt_4 ;
    wire \ADC_VDC.n20728 ;
    wire \ADC_VDC.n20729 ;
    wire \ADC_VDC.avg_cnt_6 ;
    wire \ADC_VDC.n20730 ;
    wire \ADC_VDC.avg_cnt_7 ;
    wire \ADC_VDC.n20731 ;
    wire \ADC_VDC.n20732 ;
    wire bfn_8_3_0_;
    wire \ADC_VDC.avg_cnt_9 ;
    wire \ADC_VDC.n20733 ;
    wire \ADC_VDC.n20734 ;
    wire \ADC_VDC.n20735 ;
    wire \ADC_VDC.avg_cnt_11 ;
    wire \RTD.adc_state_3 ;
    wire \RTD.adc_state_1 ;
    wire adc_state_2;
    wire \RTD.adc_state_0 ;
    wire \ADC_VDC.n22071_cascade_ ;
    wire cmd_rdadctmp_0_adj_1574;
    wire \ADC_VDC.cmd_rdadcbuf_0 ;
    wire bfn_8_6_0_;
    wire cmd_rdadctmp_1_adj_1573;
    wire \ADC_VDC.cmd_rdadcbuf_1 ;
    wire \ADC_VDC.n20690 ;
    wire cmd_rdadctmp_2_adj_1572;
    wire \ADC_VDC.cmd_rdadcbuf_2 ;
    wire \ADC_VDC.n20691 ;
    wire cmd_rdadctmp_3_adj_1571;
    wire \ADC_VDC.cmd_rdadcbuf_3 ;
    wire \ADC_VDC.n20692 ;
    wire cmd_rdadctmp_4_adj_1570;
    wire \ADC_VDC.cmd_rdadcbuf_4 ;
    wire \ADC_VDC.n20693 ;
    wire cmd_rdadctmp_5_adj_1569;
    wire \ADC_VDC.cmd_rdadcbuf_5 ;
    wire \ADC_VDC.n20694 ;
    wire cmd_rdadctmp_6_adj_1568;
    wire \ADC_VDC.cmd_rdadcbuf_6 ;
    wire \ADC_VDC.n20695 ;
    wire cmd_rdadctmp_7_adj_1567;
    wire \ADC_VDC.cmd_rdadcbuf_7 ;
    wire \ADC_VDC.n20696 ;
    wire \ADC_VDC.n20697 ;
    wire \ADC_VDC.cmd_rdadcbuf_8 ;
    wire bfn_8_7_0_;
    wire \ADC_VDC.cmd_rdadcbuf_9 ;
    wire \ADC_VDC.n20698 ;
    wire cmd_rdadctmp_10_adj_1564;
    wire \ADC_VDC.cmd_rdadcbuf_10 ;
    wire \ADC_VDC.n20699 ;
    wire cmd_rdadctmp_11_adj_1563;
    wire \ADC_VDC.n20700 ;
    wire cmd_rdadctmp_12_adj_1562;
    wire cmd_rdadcbuf_12;
    wire \ADC_VDC.n20701 ;
    wire cmd_rdadctmp_13_adj_1561;
    wire \ADC_VDC.n20702 ;
    wire cmd_rdadctmp_14_adj_1560;
    wire \ADC_VDC.n20703 ;
    wire cmd_rdadctmp_15_adj_1559;
    wire cmd_rdadcbuf_15;
    wire \ADC_VDC.n20704 ;
    wire \ADC_VDC.n20705 ;
    wire cmd_rdadctmp_16_adj_1558;
    wire bfn_8_8_0_;
    wire cmd_rdadctmp_17_adj_1557;
    wire cmd_rdadcbuf_17;
    wire \ADC_VDC.n20706 ;
    wire cmd_rdadctmp_18_adj_1556;
    wire cmd_rdadcbuf_18;
    wire \ADC_VDC.n20707 ;
    wire cmd_rdadctmp_19_adj_1555;
    wire cmd_rdadcbuf_19;
    wire \ADC_VDC.n20708 ;
    wire cmd_rdadctmp_20_adj_1554;
    wire cmd_rdadcbuf_20;
    wire \ADC_VDC.n20709 ;
    wire cmd_rdadctmp_21_adj_1553;
    wire cmd_rdadcbuf_21;
    wire \ADC_VDC.n20710 ;
    wire \ADC_VDC.n20711 ;
    wire cmd_rdadcbuf_23;
    wire \ADC_VDC.n20712 ;
    wire \ADC_VDC.n20713 ;
    wire bfn_8_9_0_;
    wire cmd_rdadcbuf_25;
    wire \ADC_VDC.n20714 ;
    wire cmd_rdadcbuf_26;
    wire \ADC_VDC.n20715 ;
    wire \ADC_VDC.n20716 ;
    wire cmd_rdadcbuf_28;
    wire \ADC_VDC.n20717 ;
    wire cmd_rdadcbuf_29;
    wire \ADC_VDC.n20718 ;
    wire cmd_rdadcbuf_30;
    wire \ADC_VDC.n20719 ;
    wire cmd_rdadcbuf_31;
    wire \ADC_VDC.n20720 ;
    wire \ADC_VDC.n20721 ;
    wire bfn_8_10_0_;
    wire cmd_rdadcbuf_33;
    wire \ADC_VDC.n20722 ;
    wire \ADC_VDC.n20723 ;
    wire n23474_cascade_;
    wire n23477_cascade_;
    wire n30_adj_1784;
    wire n112_adj_1772;
    wire n30_adj_1768_cascade_;
    wire n19_adj_1780;
    wire n30_adj_1702;
    wire n22358;
    wire buf_adcdata_vdc_19;
    wire n19_adj_1789;
    wire n23426;
    wire n23429;
    wire cmd_rdadctmp_27_adj_1521;
    wire buf_adcdata_vac_19;
    wire buf_adcdata_iac_19;
    wire buf_dds1_12;
    wire n16_adj_1778;
    wire cmd_rdadctmp_26;
    wire buf_dds1_7;
    wire IAC_SCLK;
    wire cmd_rdadctmp_21;
    wire cmd_rdadctmp_22;
    wire cmd_rdadctmp_23;
    wire \ADC_VDC.avg_cnt_0 ;
    wire \ADC_VDC.avg_cnt_5 ;
    wire \ADC_VDC.avg_cnt_8 ;
    wire \ADC_VDC.avg_cnt_10 ;
    wire \ADC_VDC.n20 ;
    wire \ADC_VDC.n19_cascade_ ;
    wire \ADC_VDC.n21 ;
    wire \ADC_VDC.n28 ;
    wire \ADC_VDC.n21871 ;
    wire \ADC_VDC.n13865 ;
    wire \ADC_VDC.n9_cascade_ ;
    wire \ADC_VDC.n22071 ;
    wire \ADC_VDC.n5 ;
    wire cmd_rdadcbuf_14;
    wire cmd_rdadctmp_8_adj_1566;
    wire n13925;
    wire cmd_rdadctmp_9_adj_1565;
    wire cmd_rdadcbuf_22;
    wire cmd_rdadcbuf_13;
    wire cmd_rdadcbuf_16;
    wire buf_adcdata_vdc_5;
    wire cmd_rdadcbuf_27;
    wire buf_dds1_5;
    wire buf_adcdata_vdc_14;
    wire buf_adcdata_vac_14;
    wire \ADC_VDC.n14120 ;
    wire \ADC_VDC.n15721 ;
    wire \ADC_VDC.cmd_rdadcbuf_35_N_1344_34 ;
    wire \ADC_VDC.n4_cascade_ ;
    wire cmd_rdadcbuf_34;
    wire \ADC_VDC.n14092 ;
    wire \comm_spi.n24028 ;
    wire \comm_spi.n24028_cascade_ ;
    wire buf_readRTD_12;
    wire n20_adj_1781;
    wire cmd_rdadctmp_19_adj_1529;
    wire cmd_rdadctmp_20_adj_1528;
    wire n23309;
    wire buf_readRTD_10;
    wire n22164_cascade_;
    wire buf_dds1_14;
    wire n23366;
    wire n16_adj_1763_cascade_;
    wire n23369;
    wire n30_adj_1698;
    wire buf_cfgRTD_6;
    wire buf_cfgRTD_2;
    wire buf_cfgRTD_4;
    wire cmd_rdadctmp_18;
    wire buf_dds1_11;
    wire data_count_0;
    wire bfn_9_14_0_;
    wire data_count_1;
    wire n20613;
    wire data_count_2;
    wire n20614;
    wire data_count_3;
    wire n20615;
    wire data_count_4;
    wire n20616;
    wire data_count_5;
    wire n20617;
    wire data_count_6;
    wire n20618;
    wire data_count_7;
    wire n20619;
    wire n20620;
    wire INVdata_count_i0_i0C_net;
    wire data_count_8;
    wire bfn_9_15_0_;
    wire n20621;
    wire data_count_9;
    wire INVdata_count_i0_i8C_net;
    wire n11983;
    wire n24_adj_1598_cascade_;
    wire n24_adj_1506_cascade_;
    wire IAC_FLT1;
    wire n11982;
    wire cmd_rdadctmp_24;
    wire cmd_rdadctmp_5;
    wire n23468;
    wire cmd_rdadctmp_25;
    wire DTRIG_N_1182;
    wire adc_state_1;
    wire cmd_rdadctmp_27;
    wire buf_adcdata_iac_17;
    wire buf_dds1_10;
    wire n22160;
    wire buf_adcdata_iac_18;
    wire IAC_FLT0;
    wire n22161;
    wire \ADC_VDC.adc_state_3_N_1316_1 ;
    wire \ADC_VDC.n22404_cascade_ ;
    wire \ADC_VDC.n17 ;
    wire \ADC_VDC.n17_cascade_ ;
    wire \ADC_VDC.n22055 ;
    wire \ADC_VDC.n27_cascade_ ;
    wire \ADC_VDC.n10 ;
    wire \ADC_VDC.n21869 ;
    wire \ADC_VDC.n11923 ;
    wire \ADC_VDC.n11923_cascade_ ;
    wire \ADC_VDC.n20869_cascade_ ;
    wire \ADC_VDC.n8031 ;
    wire \ADC_VDC.n23531 ;
    wire \ADC_VDC.n20869 ;
    wire \ADC_VDC.n21991 ;
    wire \ADC_VDC.n22075_cascade_ ;
    wire \ADC_VDC.n44_adj_1487 ;
    wire \ADC_VDC.n39_adj_1488 ;
    wire \ADC_VDC.n6_adj_1485 ;
    wire \ADC_VDC.n21859_cascade_ ;
    wire \ADC_VDC.n22628_cascade_ ;
    wire \ADC_VDC.n21859 ;
    wire \ADC_VDC.n22625 ;
    wire \ADC_VDC.n6 ;
    wire cmd_rdadctmp_22_adj_1552;
    wire \ADC_VDC.n11183_cascade_ ;
    wire \ADC_VDC.cmd_rdadctmp_23 ;
    wire \ADC_VDC.n13957 ;
    wire \ADC_VDC.n21707 ;
    wire \INVcomm_spi.imiso_83_12612_12613_resetC_net ;
    wire \comm_spi.n15369 ;
    wire buf_readRTD_13;
    wire buf_adcdata_vac_21;
    wire buf_cfgRTD_5;
    wire n23384_cascade_;
    wire cmd_rdadcbuf_32;
    wire buf_adcdata_vdc_21;
    wire cmd_rdadcbuf_24;
    wire n12352;
    wire cmd_rdadcbuf_11;
    wire buf_adcdata_vdc_12;
    wire buf_adcdata_vac_12;
    wire buf_readRTD_4;
    wire n19_adj_1734_cascade_;
    wire cmd_rdadctmp_7_adj_1541;
    wire cmd_rdadctmp_6_adj_1542;
    wire cmd_rdadctmp_5_adj_1543;
    wire cmd_rdadctmp_3_adj_1545;
    wire cmd_rdadctmp_4_adj_1544;
    wire buf_dds1_6;
    wire buf_data_iac_0;
    wire cmd_rdadctmp_21_adj_1527;
    wire n30_adj_1692;
    wire cmd_rdadctmp_25_adj_1523;
    wire buf_adcdata_vdc_18;
    wire buf_adcdata_vac_18;
    wire n22163;
    wire \comm_spi.n15360 ;
    wire \comm_spi.data_tx_7__N_857 ;
    wire comm_test_buf_24_19;
    wire comm_test_buf_24_20;
    wire n111_adj_1785;
    wire n24_cascade_;
    wire buf_adcdata_iac_22;
    wire VAC_FLT0;
    wire n17_adj_1764;
    wire n11981_cascade_;
    wire VAC_FLT1;
    wire n24_adj_1576;
    wire n11986;
    wire n23510_cascade_;
    wire n22276;
    wire n23513_cascade_;
    wire n30_adj_1759_cascade_;
    wire n26_adj_1758;
    wire eis_end;
    wire INVeis_end_302C_net;
    wire n112_adj_1762;
    wire n21946_cascade_;
    wire n21880;
    wire n13_cascade_;
    wire INVeis_state_i2C_net;
    wire n22395;
    wire cmd_rdadctmp_30;
    wire n13_adj_1591;
    wire n11_adj_1592;
    wire cmd_rdadctmp_6;
    wire acadc_dtrig_i;
    wire cmd_rdadctmp_29;
    wire DTRIG_N_1182_adj_1549;
    wire adc_state_1_adj_1515;
    wire acadc_dtrig_v;
    wire buf_dds1_9;
    wire n23534;
    wire buf_dds0_10;
    wire buf_dds0_6;
    wire buf_dds0_5;
    wire \SIG_DDS.tmp_buf_4 ;
    wire \SIG_DDS.tmp_buf_5 ;
    wire \SIG_DDS.tmp_buf_9 ;
    wire \SIG_DDS.tmp_buf_6 ;
    wire buf_dds0_7;
    wire buf_dds0_12;
    wire \SIG_DDS.tmp_buf_12 ;
    wire \SIG_DDS.tmp_buf_13 ;
    wire buf_dds0_14;
    wire \SIG_DDS.tmp_buf_14 ;
    wire buf_dds0_15;
    wire \SIG_DDS.tmp_buf_7 ;
    wire \SIG_DDS.tmp_buf_8 ;
    wire \SIG_DDS.tmp_buf_10 ;
    wire buf_dds0_11;
    wire \SIG_DDS.tmp_buf_11 ;
    wire \ADC_VDC.n22063 ;
    wire \RTD.n20050 ;
    wire VDC_SDO;
    wire \ADC_VDC.n35_cascade_ ;
    wire \ADC_VDC.n45 ;
    wire \ADC_VDC.n22067 ;
    wire adc_state_3;
    wire adc_state_1_adj_1551;
    wire \ADC_VDC.adc_state_0 ;
    wire adc_state_2_adj_1550;
    wire \ADC_VDC.n11183 ;
    wire \ADC_VDC.n23528 ;
    wire \ADC_VDC.bit_cnt_0 ;
    wire bfn_11_6_0_;
    wire \ADC_VDC.bit_cnt_1 ;
    wire \ADC_VDC.n20812 ;
    wire \ADC_VDC.bit_cnt_2 ;
    wire \ADC_VDC.n20813 ;
    wire \ADC_VDC.bit_cnt_3 ;
    wire \ADC_VDC.n20814 ;
    wire \ADC_VDC.bit_cnt_4 ;
    wire \ADC_VDC.n20815 ;
    wire \ADC_VDC.bit_cnt_5 ;
    wire \ADC_VDC.n20816 ;
    wire \ADC_VDC.bit_cnt_6 ;
    wire \ADC_VDC.n20817 ;
    wire \ADC_VDC.n20818 ;
    wire \ADC_VDC.bit_cnt_7 ;
    wire \ADC_VDC.n17565 ;
    wire \ADC_VDC.n17542 ;
    wire \comm_spi.n15361 ;
    wire buf_adcdata_vdc_3;
    wire n19_adj_1703_cascade_;
    wire buf_data_iac_3;
    wire n22_adj_1704_cascade_;
    wire buf_adcdata_iac_3;
    wire cmd_rdadctmp_11_adj_1537;
    wire buf_adcdata_vac_3;
    wire buf_adcdata_vdc_1;
    wire buf_adcdata_vac_1;
    wire n19_adj_1710_cascade_;
    wire buf_data_iac_1;
    wire n22_adj_1711_cascade_;
    wire n30_adj_1712_cascade_;
    wire \comm_spi.n24031 ;
    wire n30_adj_1705;
    wire n13847;
    wire cmd_rdadctmp_9_adj_1539;
    wire n2_adj_1666_cascade_;
    wire n1_adj_1665;
    wire \comm_spi.data_tx_7__N_865 ;
    wire comm_test_buf_24_4;
    wire n13231;
    wire n13237;
    wire n22295;
    wire n4_adj_1667;
    wire n23294;
    wire n30_adj_1588;
    wire comm_test_buf_24_3;
    wire n111_adj_1794;
    wire n15545;
    wire buf_dds1_8;
    wire comm_test_buf_24_11;
    wire comm_test_buf_24_12;
    wire buf_adcdata_iac_16;
    wire n23324;
    wire req_data_cnt_8;
    wire n19_adj_1727_cascade_;
    wire n29_adj_1770_cascade_;
    wire comm_test_buf_24_14;
    wire comm_test_buf_24_6;
    wire n16_adj_1683;
    wire n17642_cascade_;
    wire n22312;
    wire n23330;
    wire n17633;
    wire iac_raw_buf_N_821;
    wire n17_adj_1742;
    wire INVeis_state_i0C_net;
    wire n12369;
    wire n24_adj_1503;
    wire n11980;
    wire eis_state_0;
    wire eis_state_2;
    wire n12450_cascade_;
    wire cmd_rdadctmp_16;
    wire bfn_11_18_0_;
    wire INVacadc_skipcnt_i0_i0C_net;
    wire n22120;
    wire n20637;
    wire n20637_THRU_CRY_0_THRU_CO;
    wire n20637_THRU_CRY_1_THRU_CO;
    wire n20637_THRU_CRY_2_THRU_CO;
    wire n20637_THRU_CRY_3_THRU_CO;
    wire n20637_THRU_CRY_4_THRU_CO;
    wire GNDG0;
    wire n20637_THRU_CRY_5_THRU_CO;
    wire n20637_THRU_CRY_6_THRU_CO;
    wire bfn_11_19_0_;
    wire n20638;
    wire n20639;
    wire n20640;
    wire n20641;
    wire n20642;
    wire n20643;
    wire n20644;
    wire n20645;
    wire INVacadc_skipcnt_i0_i1C_net;
    wire bfn_11_20_0_;
    wire n20646;
    wire n20647;
    wire n20648;
    wire n20649;
    wire n20650;
    wire n20651;
    wire INVacadc_skipcnt_i0_i9C_net;
    wire n12450;
    wire n15439;
    wire \RTD.bit_cnt_3 ;
    wire \RTD.bit_cnt_2 ;
    wire \RTD.bit_cnt_1 ;
    wire \RTD.bit_cnt_0 ;
    wire clk_RTD;
    wire \RTD.n18274 ;
    wire \RTD.n18275 ;
    wire buf_cfgRTD_7;
    wire buf_readRTD_15;
    wire n23432;
    wire n12610_cascade_;
    wire \comm_spi.data_tx_7__N_883 ;
    wire ICE_SPI_MISO;
    wire \comm_spi.data_tx_7__N_868 ;
    wire buf_adcdata_vdc_2;
    wire n19_adj_1706_cascade_;
    wire cmd_rdadctmp_8_adj_1540;
    wire buf_adcdata_iac_1;
    wire buf_adcdata_iac_2;
    wire cmd_rdadctmp_10_adj_1538;
    wire adc_state_0_adj_1516;
    wire n21948;
    wire buf_adcdata_vac_2;
    wire cmd_rdadctmp_9;
    wire cmd_rdadctmp_10;
    wire cmd_rdadctmp_11;
    wire \comm_spi.n24034_cascade_ ;
    wire \comm_spi.n15356 ;
    wire \comm_spi.data_tx_7__N_858 ;
    wire comm_tx_buf_6;
    wire \comm_spi.n24013 ;
    wire \comm_spi.data_tx_7__N_856 ;
    wire n2_adj_1669_cascade_;
    wire n4_adj_1670_cascade_;
    wire n23402;
    wire n22669;
    wire n1_adj_1668;
    wire n13219;
    wire comm_tx_buf_4;
    wire \comm_spi.data_tx_7__N_871 ;
    wire comm_buf_0_7_N_543_4;
    wire comm_buf_0_7_N_543_6;
    wire comm_buf_0_7_N_543_7;
    wire clk_cnt_1;
    wire clk_cnt_0;
    wire n18996;
    wire comm_buf_2_7_N_575_0;
    wire comm_buf_2_7_N_575_1;
    wire comm_buf_2_7_N_575_3;
    wire comm_buf_2_7_N_575_4;
    wire comm_buf_2_7_N_575_5;
    wire comm_buf_2_7_N_575_6;
    wire comm_buf_2_6;
    wire comm_buf_2_7_N_575_7;
    wire \comm_spi.data_tx_7__N_859 ;
    wire n6774;
    wire n111_adj_1796_cascade_;
    wire comm_test_buf_24_10;
    wire \comm_spi.n15365 ;
    wire \comm_spi.n24025 ;
    wire \comm_spi.n15364 ;
    wire \comm_spi.n15368 ;
    wire \comm_spi.data_tx_7__N_855 ;
    wire AMPV_POW;
    wire n111_adj_1761;
    wire buf_dds1_3;
    wire comm_buf_2_4;
    wire n11987_cascade_;
    wire n17_adj_1779;
    wire n11985_cascade_;
    wire n13117;
    wire n15538;
    wire IAC_OSR0;
    wire n24_adj_1575;
    wire IAC_OSR1;
    wire n24_adj_1601;
    wire n11984;
    wire n16_adj_1733;
    wire n23438;
    wire buf_adcdata_iac_12;
    wire comm_test_buf_24_21;
    wire comm_test_buf_24_13;
    wire comm_test_buf_24_5;
    wire n111_adj_1776_cascade_;
    wire n11979;
    wire acadc_skipcnt_15;
    wire acadc_skipcnt_9;
    wire acadc_skipcnt_14;
    wire acadc_skipcnt_11;
    wire cmd_rdadctmp_19;
    wire cmd_rdadctmp_20;
    wire buf_dds1_0;
    wire cmd_rdadctmp_28;
    wire buf_adcdata_iac_20;
    wire buf_control_6;
    wire acadc_skipCount_14;
    wire n23_adj_1767;
    wire \SIG_DDS.tmp_buf_0 ;
    wire \SIG_DDS.tmp_buf_3 ;
    wire \SIG_DDS.tmp_buf_1 ;
    wire \SIG_DDS.tmp_buf_2 ;
    wire \comm_spi.n15323 ;
    wire \comm_spi.data_tx_7__N_860 ;
    wire \comm_spi.n24040 ;
    wire \comm_spi.data_tx_7__N_880 ;
    wire \comm_spi.n24037 ;
    wire \comm_spi.n15348 ;
    wire \comm_spi.n15349 ;
    wire \comm_spi.n15335 ;
    wire \INVcomm_spi.MISO_48_12606_12607_resetC_net ;
    wire n23390;
    wire n1_adj_1674_cascade_;
    wire comm_tx_buf_1;
    wire n22341;
    wire n2_adj_1675;
    wire buf_adcdata_vdc_0;
    wire buf_adcdata_vac_0;
    wire n19_adj_1590_cascade_;
    wire n22_adj_1589;
    wire n21965_cascade_;
    wire n13746;
    wire cmd_rdadctmp_7;
    wire comm_buf_6_4;
    wire cmd_rdadctmp_8;
    wire buf_adcdata_iac_0;
    wire buf_adcdata_vdc_13;
    wire buf_adcdata_vac_13;
    wire buf_readRTD_5;
    wire n19_adj_1729_cascade_;
    wire comm_buf_6_6;
    wire n9_adj_1600_cascade_;
    wire n6776_cascade_;
    wire n18890;
    wire comm_test_buf_24_9;
    wire comm_buf_0_7_N_543_0;
    wire comm_test_buf_24_18;
    wire comm_test_buf_24_7;
    wire comm_test_buf_24_15;
    wire comm_buf_2_1;
    wire n13201;
    wire buf_readRTD_9;
    wire buf_cfgRTD_1;
    wire \comm_spi.n15337 ;
    wire \comm_spi.n15338 ;
    wire \INVcomm_spi.imiso_83_12612_12613_setC_net ;
    wire n15496;
    wire buf_data_iac_16;
    wire n22270_cascade_;
    wire n23450_cascade_;
    wire n23327;
    wire n23453;
    wire n112_adj_1583;
    wire n23522;
    wire n22267;
    wire n112_adj_1797;
    wire comm_buf_0_7_N_543_2;
    wire comm_test_buf_24_16;
    wire n111_adj_1584;
    wire n20_adj_1804;
    wire req_data_cnt_12;
    wire VAC_OSR1;
    wire buf_adcdata_iac_21;
    wire n9_adj_1600;
    wire bfn_13_15_0_;
    wire n20652;
    wire n20653;
    wire n20654;
    wire n20655;
    wire n20656;
    wire n20657;
    wire n20658;
    wire n20659;
    wire bfn_13_16_0_;
    wire n20660;
    wire eis_stop;
    wire acadc_skipcnt_13;
    wire acadc_skipCount_13;
    wire VAC_OSR0;
    wire n40;
    wire n24_adj_1505;
    wire req_data_cnt_10;
    wire acadc_rst;
    wire data_index_9_N_236_3;
    wire acadc_skipcnt_7;
    wire acadc_skipcnt_2;
    wire acadc_skipcnt_12;
    wire acadc_skipcnt_10;
    wire n23_adj_1514;
    wire n24_adj_1513;
    wire n21_cascade_;
    wire n22;
    wire n14_adj_1610_cascade_;
    wire acadc_skipcnt_0;
    wire acadc_skipcnt_6;
    wire SELIRNG0;
    wire acadc_skipCount_10;
    wire VDC_RNG0;
    wire acadc_skipCount_12;
    wire n23_adj_1783;
    wire adc_state_0;
    wire n21951;
    wire cmd_rdadctmp_17;
    wire buf_dds0_8;
    wire data_index_1;
    wire n8_adj_1630;
    wire n8_adj_1630_cascade_;
    wire n7_adj_1629;
    wire data_index_9_N_236_1;
    wire buf_dds0_3;
    wire tmp_buf_15;
    wire DDS_MOSI;
    wire \comm_spi.n24016 ;
    wire \comm_spi.n15326 ;
    wire \comm_spi.n24016_cascade_ ;
    wire \comm_spi.n15322 ;
    wire \comm_spi.data_tx_7__N_861 ;
    wire bfn_14_5_0_;
    wire n20790;
    wire n20791;
    wire n20792;
    wire n20793;
    wire n20794;
    wire n20795;
    wire n20796;
    wire n20797;
    wire bfn_14_6_0_;
    wire n20798;
    wire n20799;
    wire n20800;
    wire n20801;
    wire n20802;
    wire n20803;
    wire n20804;
    wire n20805;
    wire bfn_14_7_0_;
    wire n20806;
    wire n20807;
    wire n20808;
    wire n20809;
    wire n20810;
    wire n20811;
    wire secclk_cnt_19;
    wire secclk_cnt_21;
    wire secclk_cnt_12;
    wire secclk_cnt_22;
    wire comm_buf_0_6;
    wire comm_buf_6_1;
    wire buf_data_iac_2;
    wire n22_adj_1707;
    wire comm_buf_2_7;
    wire n22331_cascade_;
    wire n23360_cascade_;
    wire n2_adj_1663;
    wire n4_adj_1664;
    wire n1;
    wire comm_tx_buf_7;
    wire \comm_spi.data_tx_7__N_862 ;
    wire n4_adj_1673;
    wire n22342_cascade_;
    wire n23396;
    wire n1_adj_1671_cascade_;
    wire n2_adj_1672;
    wire comm_buf_2_2;
    wire comm_buf_0_2;
    wire n13207;
    wire comm_tx_buf_2;
    wire \comm_spi.data_tx_7__N_877 ;
    wire buf_data_vac_16;
    wire buf_data_vac_23;
    wire comm_buf_3_7;
    wire buf_data_vac_22;
    wire comm_buf_3_6;
    wire buf_data_vac_21;
    wire buf_data_vac_20;
    wire comm_buf_3_4;
    wire buf_data_vac_19;
    wire buf_data_vac_18;
    wire comm_buf_3_2;
    wire buf_data_vac_17;
    wire comm_buf_3_1;
    wire n15503;
    wire n30_adj_1708;
    wire comm_test_buf_24_2;
    wire comm_buf_2_7_N_575_2;
    wire n12880;
    wire n21886;
    wire n12_cascade_;
    wire n15553;
    wire n16_adj_1721;
    wire buf_adcdata_iac_14;
    wire n12015;
    wire n8_cascade_;
    wire buf_adcdata_vdc_11;
    wire buf_adcdata_vac_11;
    wire n22092;
    wire n13211;
    wire acadc_skipcnt_5;
    wire acadc_skipcnt_3;
    wire acadc_skipCount_15;
    wire n23_adj_1756;
    wire n21_adj_1803;
    wire n30_adj_1769;
    wire n22167;
    wire n22166;
    wire n23471;
    wire n23549_cascade_;
    wire n22174;
    wire n112;
    wire n30_adj_1805;
    wire n17650;
    wire n12;
    wire buf_data_iac_12;
    wire data_index_2;
    wire n8_adj_1628;
    wire n8_adj_1628_cascade_;
    wire n7_adj_1627;
    wire data_index_9_N_236_2;
    wire n18865;
    wire n7_adj_1626;
    wire data_index_3;
    wire acadc_skipcnt_8;
    wire n20;
    wire n14_adj_1599;
    wire n17;
    wire n26_cascade_;
    wire n30_adj_1743;
    wire n31;
    wire buf_dds0_1;
    wire buf_dds1_1;
    wire buf_dds1_2;
    wire buf_adcdata_iac_10;
    wire n16_adj_1746_cascade_;
    wire \comm_spi.n15341 ;
    wire \comm_spi.n15340 ;
    wire \comm_spi.n15333 ;
    wire \comm_spi.n15334 ;
    wire \INVcomm_spi.MISO_48_12606_12607_setC_net ;
    wire \comm_spi.data_tx_7__N_854 ;
    wire comm_test_buf_24_1;
    wire n111_adj_1798;
    wire n21965;
    wire n12056_cascade_;
    wire comm_test_buf_24_23;
    wire buf_dds0_2;
    wire data_index_9;
    wire n8_adj_1617_cascade_;
    wire data_index_9_N_236_8;
    wire \SIG_DDS.n13338 ;
    wire \comm_spi.iclk_N_850 ;
    wire \comm_spi.n15327 ;
    wire VDC_CLK;
    wire \INVADC_VDC.genclk.t_clk_24C_net ;
    wire n4_adj_1676;
    wire \comm_spi.DOUT_7__N_835 ;
    wire ICE_SPI_SCLK;
    wire \comm_spi.iclk_N_851 ;
    wire secclk_cnt_15;
    wire secclk_cnt_8;
    wire secclk_cnt_1;
    wire secclk_cnt_5;
    wire n25_adj_1717_cascade_;
    wire secclk_cnt_20;
    wire n20922_cascade_;
    wire n14_adj_1678;
    wire secclk_cnt_9;
    wire secclk_cnt_17;
    wire n10_adj_1679;
    wire secclk_cnt_6;
    wire secclk_cnt_14;
    wire secclk_cnt_10;
    wire secclk_cnt_3;
    wire n27;
    wire secclk_cnt_16;
    wire secclk_cnt_7;
    wire secclk_cnt_13;
    wire secclk_cnt_2;
    wire n26_adj_1715;
    wire n15420;
    wire TEST_LED;
    wire n9_adj_1596;
    wire comm_buf_6_7;
    wire comm_test_buf_24_17;
    wire comm_buf_6_0;
    wire n18818_cascade_;
    wire n23372_cascade_;
    wire n18816;
    wire comm_tx_buf_0;
    wire comm_buf_3_0;
    wire n22338;
    wire n18815;
    wire comm_buf_2_0;
    wire n18823;
    wire buf_data_vac_0;
    wire comm_buf_5_0;
    wire buf_data_vac_7;
    wire comm_buf_5_7;
    wire buf_data_vac_6;
    wire comm_buf_5_6;
    wire buf_data_vac_5;
    wire buf_data_vac_4;
    wire comm_buf_5_4;
    wire buf_data_vac_3;
    wire buf_data_vac_2;
    wire comm_buf_5_2;
    wire buf_data_vac_1;
    wire comm_buf_5_1;
    wire buf_readRTD_8;
    wire buf_adcdata_vdc_16;
    wire n23504_cascade_;
    wire buf_adcdata_vac_16;
    wire n22288;
    wire n12838;
    wire n23306;
    wire n8_adj_1504;
    wire n6_cascade_;
    wire n21938;
    wire n19_adj_1722;
    wire buf_readRTD_6;
    wire n23288;
    wire n22396_cascade_;
    wire n6;
    wire n22061;
    wire n21929;
    wire n22_adj_1801;
    wire n112_adj_1799;
    wire comm_buf_0_7_N_543_1;
    wire n18_adj_1699;
    wire n13257;
    wire acadc_skipcnt_1;
    wire acadc_skipcnt_4;
    wire n18;
    wire comm_buf_0_0;
    wire n11172;
    wire eis_start;
    wire n8_adj_1625_cascade_;
    wire data_index_9_N_236_4;
    wire n7_adj_1624;
    wire n8_adj_1625;
    wire data_index_4;
    wire n23546;
    wire n30;
    wire n17_adj_1594;
    wire acadc_skipCount_8;
    wire n24_adj_1800;
    wire req_data_cnt_9;
    wire req_data_cnt_15;
    wire n22314;
    wire n22169;
    wire req_data_cnt_3;
    wire n23312_cascade_;
    wire n23315_cascade_;
    wire n111_adj_1744;
    wire n30_adj_1741_cascade_;
    wire acadc_skipCount_3;
    wire n19_adj_1739;
    wire buf_readRTD_3;
    wire buf_adcdata_iac_11;
    wire n16_adj_1738;
    wire n23558_cascade_;
    wire n23561;
    wire \SIG_DDS.bit_cnt_2 ;
    wire \SIG_DDS.bit_cnt_1 ;
    wire comm_buf_0_4;
    wire comm_buf_0_1;
    wire \SIG_DDS.bit_cnt_3 ;
    wire n8_adj_1615;
    wire n7_adj_1614;
    wire data_index_9_N_236_9;
    wire data_index_6;
    wire n8_adj_1621;
    wire n8_adj_1621_cascade_;
    wire n7_adj_1620;
    wire data_index_9_N_236_6;
    wire data_index_7;
    wire n8_adj_1617;
    wire n7_adj_1616;
    wire data_index_8;
    wire n8_adj_1619;
    wire n7_adj_1618;
    wire data_index_9_N_236_7;
    wire \SIG_DDS.n22671 ;
    wire \SIG_DDS.n10 ;
    wire \comm_spi.imosi_N_841 ;
    wire \comm_spi.n15331 ;
    wire \comm_spi.imosi_cascade_ ;
    wire \comm_spi.n24019 ;
    wire \comm_spi.n15344 ;
    wire \comm_spi.n15345 ;
    wire \comm_spi.n24019_cascade_ ;
    wire secclk_cnt_0;
    wire secclk_cnt_18;
    wire secclk_cnt_11;
    wire secclk_cnt_4;
    wire n28;
    wire n12_adj_1760_cascade_;
    wire n20834_cascade_;
    wire n30_adj_1681;
    wire n33;
    wire n32;
    wire n34_cascade_;
    wire n31_adj_1680;
    wire n49_cascade_;
    wire \comm_spi.n24022 ;
    wire n8856_cascade_;
    wire n13273;
    wire comm_buf_0_5;
    wire comm_buf_3_5;
    wire comm_buf_6_5;
    wire comm_buf_2_5;
    wire n18882;
    wire n18883_cascade_;
    wire comm_tx_buf_5;
    wire comm_buf_5_5;
    wire n22371;
    wire n18885_cascade_;
    wire n23414;
    wire n22618;
    wire n8_adj_1755;
    wire n12976;
    wire n12976_cascade_;
    wire comm_buf_6_2;
    wire n22375_cascade_;
    wire buf_data_iac_22;
    wire n22297;
    wire \INVcomm_spi.bit_cnt_3787__i3C_net ;
    wire eis_state_1;
    wire n15517;
    wire n12585;
    wire n15238;
    wire n12958;
    wire n22397;
    wire n29_adj_1688;
    wire n11402_cascade_;
    wire comm_state_3_N_500_2;
    wire n18850_cascade_;
    wire n13076;
    wire n15531;
    wire comm_buf_3_3;
    wire comm_buf_6_3;
    wire n18851;
    wire comm_buf_5_3;
    wire n22346;
    wire n18853_cascade_;
    wire n23378;
    wire n6776;
    wire comm_buf_2_3;
    wire n18858;
    wire comm_tx_buf_3;
    wire THERMOSTAT;
    wire buf_control_7;
    wire n12021_cascade_;
    wire n12614;
    wire n25_cascade_;
    wire n12548;
    wire comm_buf_0_7;
    wire n21964;
    wire n11379;
    wire n9;
    wire n22059;
    wire n26_adj_1740;
    wire n26_adj_1580_cascade_;
    wire acadc_skipCount_0;
    wire n23552_cascade_;
    wire req_data_cnt_0;
    wire n16;
    wire n23300;
    wire buf_adcdata_iac_8;
    wire buf_adcdata_iac_15;
    wire n16_adj_1713;
    wire n22268;
    wire n13141;
    wire n12610;
    wire buf_dds0_4;
    wire buf_dds0_0;
    wire data_idxvec_0;
    wire bfn_16_16_0_;
    wire n14_adj_1613;
    wire n20661;
    wire n14_adj_1612;
    wire n20662;
    wire data_idxvec_3;
    wire n20663;
    wire n20664;
    wire n14_adj_1661;
    wire n20665;
    wire n14_adj_1610;
    wire n20666;
    wire n14_adj_1609;
    wire n20667;
    wire n20668;
    wire data_idxvec_8;
    wire bfn_16_17_0_;
    wire n20669;
    wire n14_adj_1655;
    wire data_idxvec_10;
    wire n20670;
    wire n20671;
    wire n14_adj_1653;
    wire n20672;
    wire n20673;
    wire n20674;
    wire n14_adj_1607;
    wire n20675;
    wire data_idxvec_15;
    wire data_index_0;
    wire n11254;
    wire n13052;
    wire n15562;
    wire n15562_cascade_;
    wire bit_cnt_0;
    wire \SIG_DDS.n9 ;
    wire DDS_SCK;
    wire trig_dds0;
    wire \comm_spi.imosi ;
    wire \comm_spi.DOUT_7__N_834 ;
    wire \comm_spi.n15330 ;
    wire wdtick_cnt_0;
    wire bfn_17_5_0_;
    wire wdtick_cnt_1;
    wire n20766;
    wire wdtick_cnt_2;
    wire n20767;
    wire wdtick_cnt_3;
    wire n20768;
    wire wdtick_cnt_4;
    wire n20769;
    wire wdtick_cnt_5;
    wire n20770;
    wire wdtick_cnt_6;
    wire n20771;
    wire wdtick_cnt_7;
    wire n20772;
    wire n20773;
    wire wdtick_cnt_8;
    wire bfn_17_6_0_;
    wire wdtick_cnt_9;
    wire n20774;
    wire wdtick_cnt_10;
    wire n20775;
    wire wdtick_cnt_11;
    wire n20776;
    wire wdtick_cnt_12;
    wire n20777;
    wire wdtick_cnt_13;
    wire n20778;
    wire wdtick_cnt_14;
    wire n20779;
    wire wdtick_cnt_15;
    wire n20780;
    wire n20781;
    wire wdtick_cnt_16;
    wire bfn_17_7_0_;
    wire wdtick_cnt_17;
    wire n20782;
    wire wdtick_cnt_18;
    wire n20783;
    wire wdtick_cnt_19;
    wire n20784;
    wire wdtick_cnt_20;
    wire n20785;
    wire wdtick_cnt_21;
    wire n20786;
    wire wdtick_cnt_22;
    wire n20787;
    wire wdtick_cnt_23;
    wire n20788;
    wire n20789;
    wire n49;
    wire bfn_17_8_0_;
    wire wdtick_cnt_24;
    wire DDS_MCLK1;
    wire n12366;
    wire n7_adj_1757;
    wire n2562_cascade_;
    wire n15378;
    wire n8_adj_1782;
    wire n12540;
    wire n14_adj_1606;
    wire n22238;
    wire n22240_cascade_;
    wire n23053;
    wire n11280_cascade_;
    wire n12509_cascade_;
    wire comm_length_2;
    wire comm_length_0;
    wire buf_adcdata_vac_17;
    wire n23486;
    wire buf_adcdata_vdc_17;
    wire n46_cascade_;
    wire comm_test_buf_24_0;
    wire comm_test_buf_24_8;
    wire n14_adj_1662;
    wire n4_adj_1749;
    wire n12_adj_1684;
    wire n14_adj_1608;
    wire n13129;
    wire buf_cfgRTD_0;
    wire n22351;
    wire n4_adj_1709_cascade_;
    wire n35;
    wire n12_adj_1802;
    wire comm_buf_1_7_N_559_3;
    wire comm_buf_1_3;
    wire comm_buf_1_6;
    wire comm_buf_1_0;
    wire data_idxvec_14;
    wire n22296;
    wire data_idxvec_12;
    wire n22499;
    wire acadc_skipCount_6;
    wire req_data_cnt_6;
    wire n23519_cascade_;
    wire n23291;
    wire n111_adj_1726;
    wire n30_adj_1724_cascade_;
    wire comm_buf_1_7_N_559_6;
    wire data_idxvec_6;
    wire n26_adj_1723_cascade_;
    wire n23516;
    wire n23303;
    wire n23555;
    wire n18363;
    wire buf_dds1_4;
    wire iac_raw_buf_N_823;
    wire data_cntvec_0;
    wire bfn_17_15_0_;
    wire n20622;
    wire n20623;
    wire data_cntvec_3;
    wire n20624;
    wire n20625;
    wire n20626;
    wire data_cntvec_6;
    wire n20627;
    wire n20628;
    wire n20629;
    wire INVdata_cntvec_i0_i0C_net;
    wire data_cntvec_8;
    wire bfn_17_16_0_;
    wire n20630;
    wire data_cntvec_10;
    wire n20631;
    wire n20632;
    wire data_cntvec_12;
    wire n20633;
    wire data_cntvec_13;
    wire n20634;
    wire n20635;
    wire n20636;
    wire data_cntvec_15;
    wire INVdata_cntvec_i0_i8C_net;
    wire n12394;
    wire n15431;
    wire n23480;
    wire DDS_RNG_0;
    wire acadc_skipCount_9;
    wire n22183_cascade_;
    wire n22177;
    wire n22180;
    wire n23462_cascade_;
    wire n23465;
    wire data_idxvec_9;
    wire data_cntvec_9;
    wire buf_data_iac_17;
    wire n22184_cascade_;
    wire n22186;
    wire n21997;
    wire n14_adj_1656;
    wire n13093;
    wire buf_dds0_9;
    wire dds_state_0;
    wire dds_state_2;
    wire dds_state_1;
    wire DDS_CS;
    wire \SIG_DDS.n9_adj_1490 ;
    wire buf_data_iac_23;
    wire n22595;
    wire ICE_SPI_MOSI;
    wire \comm_spi.imosi_N_840 ;
    wire \comm_spi.n24034 ;
    wire \comm_spi.n15352 ;
    wire \comm_spi.n15353 ;
    wire \comm_spi.n15357 ;
    wire \comm_spi.data_tx_7__N_874 ;
    wire n22489_cascade_;
    wire n20959_cascade_;
    wire n21883;
    wire n19241;
    wire n22033;
    wire n12064_cascade_;
    wire n21885;
    wire n22073_cascade_;
    wire flagcntwd;
    wire n12050;
    wire n10_adj_1602;
    wire comm_cmd_7;
    wire n29;
    wire n12951;
    wire n9714;
    wire n11_adj_1585;
    wire n14_adj_1652;
    wire \comm_spi.bit_cnt_1 ;
    wire \comm_spi.bit_cnt_0 ;
    wire \comm_spi.bit_cnt_2 ;
    wire n22487;
    wire n21983;
    wire n13171;
    wire n13171_cascade_;
    wire n22354;
    wire n22353;
    wire comm_length_1;
    wire n4_adj_1745;
    wire comm_index_1;
    wire req_data_cnt_14;
    wire data_cntvec_14;
    wire n23;
    wire n111;
    wire n30_adj_1579;
    wire comm_buf_1_7_N_559_0;
    wire n21271;
    wire n11258;
    wire n22089;
    wire n20318;
    wire n12_adj_1677_cascade_;
    wire n12892_cascade_;
    wire n37_cascade_;
    wire n12761_cascade_;
    wire data_idxvec_5;
    wire data_cntvec_5;
    wire n26_adj_1730_cascade_;
    wire req_data_cnt_5;
    wire n23336_cascade_;
    wire acadc_skipCount_5;
    wire n23339_cascade_;
    wire n30_adj_1731_cascade_;
    wire n111_adj_1732;
    wire comm_buf_1_7_N_559_5_cascade_;
    wire n16_adj_1728;
    wire buf_adcdata_iac_13;
    wire n23354;
    wire n23357;
    wire data_idxvec_1;
    wire data_cntvec_1;
    wire acadc_skipCount_1;
    wire req_data_cnt_1;
    wire n22142_cascade_;
    wire n22137;
    wire n23408_cascade_;
    wire n23411_cascade_;
    wire n111_adj_1754;
    wire comm_buf_1_7_N_559_1_cascade_;
    wire comm_buf_1_1;
    wire buf_data_iac_9;
    wire n26_adj_1753;
    wire n22143;
    wire data_idxvec_4;
    wire data_cntvec_4;
    wire n22301;
    wire n26_adj_1735_cascade_;
    wire acadc_skipCount_4;
    wire n23318_cascade_;
    wire req_data_cnt_4;
    wire n23441;
    wire n23321_cascade_;
    wire n111_adj_1737;
    wire n30_adj_1736_cascade_;
    wire comm_buf_1_7_N_559_4_cascade_;
    wire data_idxvec_2;
    wire data_cntvec_2;
    wire buf_data_iac_10;
    wire n26_adj_1748_cascade_;
    wire n22152_cascade_;
    wire n22149;
    wire n23444_cascade_;
    wire n22148;
    wire n111_adj_1750;
    wire n23447_cascade_;
    wire comm_buf_1_7_N_559_2_cascade_;
    wire comm_buf_1_2;
    wire req_data_cnt_2;
    wire acadc_skipCount_2;
    wire n22151;
    wire SELIRNG1;
    wire acadc_skipCount_11;
    wire buf_adcdata_iac_9;
    wire n16_adj_1751;
    wire n22136;
    wire wdtick_flag;
    wire buf_control_0;
    wire CONT_SD;
    wire n8_adj_1605;
    wire n7;
    wire data_index_9_N_236_0;
    wire buf_data_iac_20;
    wire n22500;
    wire bfn_19_5_0_;
    wire \ADC_VDC.genclk.n20751 ;
    wire \ADC_VDC.genclk.n20752 ;
    wire \ADC_VDC.genclk.n20753 ;
    wire \ADC_VDC.genclk.n20754 ;
    wire \ADC_VDC.genclk.n20755 ;
    wire \ADC_VDC.genclk.n20756 ;
    wire \ADC_VDC.genclk.n20757 ;
    wire \ADC_VDC.genclk.n20758 ;
    wire \INVADC_VDC.genclk.t0on_i0C_net ;
    wire bfn_19_6_0_;
    wire \ADC_VDC.genclk.n20759 ;
    wire \ADC_VDC.genclk.n20760 ;
    wire \ADC_VDC.genclk.n20761 ;
    wire \ADC_VDC.genclk.n20762 ;
    wire \ADC_VDC.genclk.n20763 ;
    wire \ADC_VDC.genclk.n20764 ;
    wire \ADC_VDC.genclk.n20765 ;
    wire \INVADC_VDC.genclk.t0on_i8C_net ;
    wire bfn_19_7_0_;
    wire n20819;
    wire n20820;
    wire n20821;
    wire n20822;
    wire n20823;
    wire n20824;
    wire n20825;
    wire INVdds0_mclkcnt_i7_3792__i0C_net;
    wire n10;
    wire dds0_mclkcnt_6;
    wire DDS_MCLK;
    wire INVdds0_mclk_297C_net;
    wire n6888_cascade_;
    wire n21865;
    wire n21981;
    wire n22027;
    wire n22018;
    wire dds0_mclkcnt_3;
    wire dds0_mclkcnt_5;
    wire dds0_mclkcnt_1;
    wire dds0_mclkcnt_4;
    wire dds0_mclkcnt_7;
    wire dds0_mclkcnt_0;
    wire n12_adj_1685_cascade_;
    wire dds0_mclkcnt_2;
    wire n21857;
    wire \INVcomm_spi.data_valid_85C_net ;
    wire \comm_spi.bit_cnt_3 ;
    wire \comm_spi.n18536 ;
    wire \comm_spi.iclk ;
    wire n22330;
    wire n22329;
    wire n15261;
    wire n22321_cascade_;
    wire n14851;
    wire n22352;
    wire comm_index_2;
    wire n21956;
    wire n21862;
    wire comm_index_0;
    wire n21862_cascade_;
    wire n30_adj_1720;
    wire n21968;
    wire n22_adj_1725_cascade_;
    wire n12677_cascade_;
    wire n21895;
    wire buf_data_vac_8;
    wire comm_rx_buf_0;
    wire comm_buf_4_0;
    wire buf_data_vac_15;
    wire comm_buf_4_7;
    wire comm_rx_buf_6;
    wire buf_data_vac_14;
    wire comm_buf_4_6;
    wire comm_rx_buf_5;
    wire buf_data_vac_13;
    wire comm_buf_4_5;
    wire comm_rx_buf_4;
    wire buf_data_vac_12;
    wire comm_buf_4_4;
    wire buf_data_vac_11;
    wire comm_buf_4_3;
    wire comm_rx_buf_2;
    wire buf_data_vac_10;
    wire comm_buf_4_2;
    wire comm_rx_buf_1;
    wire buf_data_vac_9;
    wire comm_buf_4_1;
    wire n12892;
    wire n15510;
    wire data_idxvec_7;
    wire data_cntvec_7;
    wire buf_data_iac_15;
    wire n26_adj_1716_cascade_;
    wire n22263_cascade_;
    wire n22272;
    wire n23420_cascade_;
    wire n22271;
    wire n111_adj_1719;
    wire n23423_cascade_;
    wire comm_rx_buf_7;
    wire comm_buf_1_7_N_559_7_cascade_;
    wire comm_buf_1_7;
    wire n12761;
    wire n15489;
    wire n18955;
    wire n22356;
    wire buf_dds0_13;
    wire n23348;
    wire req_data_cnt_7;
    wire acadc_skipCount_7;
    wire n22262;
    wire buf_data_iac_14;
    wire n22391;
    wire n12509;
    wire n14_adj_1660;
    wire buf_dds1_13;
    wire comm_buf_1_5;
    wire data_index_5;
    wire n9324;
    wire n8_adj_1623;
    wire n8_adj_1623_cascade_;
    wire n7_adj_1622;
    wire data_index_9_N_236_5;
    wire n21966;
    wire trig_dds1;
    wire n21920;
    wire n22399_cascade_;
    wire n40_adj_1689;
    wire data_idxvec_11;
    wire data_cntvec_11;
    wire comm_buf_1_4;
    wire n14_adj_1611;
    wire n14_adj_1654;
    wire \INVADC_VDC.genclk.div_state_i1C_net ;
    wire \ADC_VDC.genclk.n6 ;
    wire \ADC_VDC.genclk.t0on_6 ;
    wire \ADC_VDC.genclk.t0on_1 ;
    wire \ADC_VDC.genclk.t0on_4 ;
    wire \ADC_VDC.genclk.t0on_0 ;
    wire \ADC_VDC.genclk.n22308_cascade_ ;
    wire \ADC_VDC.genclk.t0on_12 ;
    wire \ADC_VDC.genclk.t0on_2 ;
    wire \ADC_VDC.genclk.t0on_7 ;
    wire \ADC_VDC.genclk.t0on_10 ;
    wire \ADC_VDC.genclk.n27_adj_1483 ;
    wire \ADC_VDC.genclk.t0on_14 ;
    wire \ADC_VDC.genclk.t0on_9 ;
    wire \ADC_VDC.genclk.t0on_15 ;
    wire \ADC_VDC.genclk.t0on_11 ;
    wire \ADC_VDC.genclk.n28_adj_1481 ;
    wire \ADC_VDC.genclk.t0on_13 ;
    wire \ADC_VDC.genclk.t0on_3 ;
    wire \ADC_VDC.genclk.t0on_5 ;
    wire \ADC_VDC.genclk.t0on_8 ;
    wire \ADC_VDC.genclk.n26_adj_1482 ;
    wire \ADC_VDC.genclk.div_state_1__N_1480 ;
    wire comm_clear;
    wire buf_data_iac_18;
    wire n22170;
    wire n12035;
    wire n7_adj_1687;
    wire comm_state_3_N_484_3;
    wire n1373;
    wire n2_cascade_;
    wire n23342;
    wire n9837;
    wire n23345_cascade_;
    wire n8_adj_1659;
    wire n2562;
    wire n22339;
    wire n22340_cascade_;
    wire n14_adj_1593;
    wire n5;
    wire n9725_cascade_;
    wire n4;
    wire n22492;
    wire n6_adj_1657_cascade_;
    wire n26_adj_1597_cascade_;
    wire n18_adj_1595;
    wire n21908;
    wire ICE_SPI_CE0;
    wire comm_data_vld;
    wire n4_adj_1718;
    wire req_data_cnt_11;
    wire n112_adj_1777;
    wire comm_buf_0_7_N_543_5;
    wire comm_cmd_5;
    wire comm_cmd_4;
    wire n22365;
    wire n22364_cascade_;
    wire n48;
    wire n22370_cascade_;
    wire n7148;
    wire n22368;
    wire n9_adj_1507;
    wire n23387;
    wire n23351;
    wire n23495;
    wire buf_data_iac_19;
    wire n22642;
    wire n23_adj_1791;
    wire n23501;
    wire n23459_cascade_;
    wire n112_adj_1795;
    wire n30_adj_1793_cascade_;
    wire comm_cmd_6;
    wire data_idxvec_13;
    wire buf_data_iac_21;
    wire n28_adj_1775_cascade_;
    wire comm_cmd_3;
    wire n23492;
    wire n23_adj_1773;
    wire req_data_cnt_13;
    wire n25_adj_1774;
    wire comm_cmd_1;
    wire comm_cmd_2;
    wire n22316;
    wire n26_adj_1792;
    wire n23456;
    wire buf_data_iac_13;
    wire n22313;
    wire buf_data_iac_11;
    wire n22300;
    wire buf_data_iac_8;
    wire comm_cmd_0;
    wire n22649;
    wire \ADC_VDC.genclk.n26 ;
    wire \ADC_VDC.genclk.n22305_cascade_ ;
    wire \ADC_VDC.genclk.n27 ;
    wire \ADC_VDC.genclk.n22303 ;
    wire \ADC_VDC.genclk.div_state_1 ;
    wire \ADC_VDC.genclk.n22303_cascade_ ;
    wire \ADC_VDC.genclk.n22302 ;
    wire \ADC_VDC.genclk.div_state_0 ;
    wire \INVADC_VDC.genclk.div_state_i0C_net ;
    wire \ADC_VDC.genclk.n28 ;
    wire ICE_GPMI_0;
    wire comm_state_2;
    wire comm_state_3;
    wire n12966;
    wire comm_state_0;
    wire n12045;
    wire comm_rx_buf_3;
    wire comm_state_1;
    wire comm_buf_0_7_N_543_3;
    wire comm_buf_0_3;
    wire clk_32MHz;
    wire n12677;
    wire n15482;
    wire \ADC_VDC.genclk.t0off_0 ;
    wire bfn_23_5_0_;
    wire \ADC_VDC.genclk.t0off_1 ;
    wire \ADC_VDC.genclk.n20736 ;
    wire \ADC_VDC.genclk.t0off_2 ;
    wire \ADC_VDC.genclk.n20737 ;
    wire \ADC_VDC.genclk.t0off_3 ;
    wire \ADC_VDC.genclk.n20738 ;
    wire \ADC_VDC.genclk.t0off_4 ;
    wire \ADC_VDC.genclk.n20739 ;
    wire \ADC_VDC.genclk.t0off_5 ;
    wire \ADC_VDC.genclk.n20740 ;
    wire \ADC_VDC.genclk.t0off_6 ;
    wire \ADC_VDC.genclk.n20741 ;
    wire \ADC_VDC.genclk.t0off_7 ;
    wire \ADC_VDC.genclk.n20742 ;
    wire \ADC_VDC.genclk.n20743 ;
    wire \INVADC_VDC.genclk.t0off_i0C_net ;
    wire \ADC_VDC.genclk.t0off_8 ;
    wire bfn_23_6_0_;
    wire \ADC_VDC.genclk.t0off_9 ;
    wire \ADC_VDC.genclk.n20744 ;
    wire \ADC_VDC.genclk.t0off_10 ;
    wire \ADC_VDC.genclk.n20745 ;
    wire \ADC_VDC.genclk.t0off_11 ;
    wire \ADC_VDC.genclk.n20746 ;
    wire \ADC_VDC.genclk.t0off_12 ;
    wire \ADC_VDC.genclk.n20747 ;
    wire \ADC_VDC.genclk.t0off_13 ;
    wire \ADC_VDC.genclk.n20748 ;
    wire \ADC_VDC.genclk.t0off_14 ;
    wire \ADC_VDC.genclk.n20749 ;
    wire CONSTANT_ONE_NET;
    wire \ADC_VDC.genclk.n20750 ;
    wire \ADC_VDC.genclk.t0off_15 ;
    wire _gnd_net_;
    wire \INVADC_VDC.genclk.t0off_i8C_net ;
    wire \ADC_VDC.genclk.n12361 ;
    wire \ADC_VDC.genclk.n15418 ;

    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_main.zim_pll_inst .TEST_MODE=1'b0;
    defparam \pll_main.zim_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll_main.zim_pll_inst .FILTER_RANGE=3'b011;
    defparam \pll_main.zim_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_main.zim_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_main.zim_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll_main.zim_pll_inst .DIVR=4'b0000;
    defparam \pll_main.zim_pll_inst .DIVQ=3'b101;
    defparam \pll_main.zim_pll_inst .DIVF=7'b0011111;
    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll_main.zim_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(),
            .REFERENCECLK(N__21256),
            .RESETB(N__64855),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(DDS_MCLK1),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(clk_32MHz),
            .SCLK(GNDG0));
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged2_physical (
            .RDATA({dangling_wire_0,dangling_wire_1,buf_data_iac_19,dangling_wire_2,dangling_wire_3,dangling_wire_4,buf_data_vac_19,dangling_wire_5,dangling_wire_6,dangling_wire_7,buf_data_iac_18,dangling_wire_8,dangling_wire_9,dangling_wire_10,buf_data_vac_18,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__44452,N__42274,N__44878,N__45073,N__56338,N__43771,N__39061,N__41731,N__40135,N__53098}),
            .WADDR({dangling_wire_13,N__29899,N__30007,N__30115,N__30214,N__29152,N__29260,N__29365,N__29473,N__29584,N__29686}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__28003,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__27841,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__30610,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__31495,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__61922),
            .RE(N__64829),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .WE(N__34523));
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged7_physical (
            .RDATA({dangling_wire_42,dangling_wire_43,buf_data_iac_9,dangling_wire_44,dangling_wire_45,dangling_wire_46,buf_data_vac_9,dangling_wire_47,dangling_wire_48,dangling_wire_49,buf_data_iac_8,dangling_wire_50,dangling_wire_51,dangling_wire_52,buf_data_vac_8,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__44412,N__42231,N__44835,N__45030,N__56289,N__43725,N__39018,N__41685,N__40092,N__53055}),
            .WADDR({dangling_wire_55,N__29865,N__29970,N__30078,N__30180,N__29115,N__29223,N__29328,N__29439,N__29553,N__29649}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__52720,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__23878,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__46956,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__25300,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__62013),
            .RE(N__64873),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .WE(N__34522));
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged1_physical (
            .RDATA({dangling_wire_84,dangling_wire_85,buf_data_iac_21,dangling_wire_86,dangling_wire_87,dangling_wire_88,buf_data_vac_21,dangling_wire_89,dangling_wire_90,dangling_wire_91,buf_data_iac_20,dangling_wire_92,dangling_wire_93,dangling_wire_94,buf_data_vac_20,dangling_wire_95}),
            .RADDR({dangling_wire_96,N__44470,N__42292,N__44896,N__45091,N__56356,N__43789,N__39079,N__41749,N__40153,N__53116}),
            .WADDR({dangling_wire_97,N__29917,N__30025,N__30133,N__30232,N__29170,N__29278,N__29383,N__29491,N__29602,N__29704}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({dangling_wire_114,dangling_wire_115,N__38623,dangling_wire_116,dangling_wire_117,dangling_wire_118,N__31210,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__37171,dangling_wire_122,dangling_wire_123,dangling_wire_124,N__25459,dangling_wire_125}),
            .RCLKE(),
            .RCLK(N__61852),
            .RE(N__64824),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .WE(N__34536));
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged6_physical (
            .RDATA({dangling_wire_126,dangling_wire_127,buf_data_iac_11,dangling_wire_128,dangling_wire_129,dangling_wire_130,buf_data_vac_11,dangling_wire_131,dangling_wire_132,dangling_wire_133,buf_data_iac_10,dangling_wire_134,dangling_wire_135,dangling_wire_136,buf_data_vac_10,dangling_wire_137}),
            .RADDR({dangling_wire_138,N__44424,N__42243,N__44847,N__45042,N__56301,N__43737,N__39030,N__41697,N__40104,N__53067}),
            .WADDR({dangling_wire_139,N__29875,N__29982,N__30090,N__30190,N__29127,N__29235,N__29340,N__29449,N__29560,N__29661}),
            .MASK({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155}),
            .WDATA({dangling_wire_156,dangling_wire_157,N__44229,dangling_wire_158,dangling_wire_159,dangling_wire_160,N__41230,dangling_wire_161,dangling_wire_162,dangling_wire_163,N__42076,dangling_wire_164,dangling_wire_165,dangling_wire_166,N__25087,dangling_wire_167}),
            .RCLKE(),
            .RCLK(N__62010),
            .RE(N__64869),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .WE(N__34499));
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged0_physical (
            .RDATA({dangling_wire_168,dangling_wire_169,buf_data_iac_23,dangling_wire_170,dangling_wire_171,dangling_wire_172,buf_data_vac_23,dangling_wire_173,dangling_wire_174,dangling_wire_175,buf_data_iac_22,dangling_wire_176,dangling_wire_177,dangling_wire_178,buf_data_vac_22,dangling_wire_179}),
            .RADDR({dangling_wire_180,N__44476,N__42298,N__44902,N__45097,N__56362,N__43795,N__39085,N__41755,N__40159,N__53122}),
            .WADDR({dangling_wire_181,N__29923,N__30031,N__30139,N__30238,N__29176,N__29284,N__29389,N__29497,N__29608,N__29710}),
            .MASK({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .WDATA({dangling_wire_198,dangling_wire_199,N__25402,dangling_wire_200,dangling_wire_201,dangling_wire_202,N__23254,dangling_wire_203,dangling_wire_204,dangling_wire_205,N__31690,dangling_wire_206,dangling_wire_207,dangling_wire_208,N__23104,dangling_wire_209}),
            .RCLKE(),
            .RCLK(N__61837),
            .RE(N__64856),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .WE(N__34540));
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged5_physical (
            .RDATA({dangling_wire_210,dangling_wire_211,buf_data_iac_13,dangling_wire_212,dangling_wire_213,dangling_wire_214,buf_data_vac_13,dangling_wire_215,dangling_wire_216,dangling_wire_217,buf_data_iac_12,dangling_wire_218,dangling_wire_219,dangling_wire_220,buf_data_vac_12,dangling_wire_221}),
            .RADDR({dangling_wire_222,N__44434,N__42255,N__44859,N__45054,N__56313,N__43749,N__39042,N__41709,N__40116,N__53079}),
            .WADDR({dangling_wire_223,N__29881,N__29989,N__30097,N__30196,N__29134,N__29242,N__29347,N__29455,N__29566,N__29668}),
            .MASK({dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .WDATA({dangling_wire_240,dangling_wire_241,N__52341,dangling_wire_242,dangling_wire_243,dangling_wire_244,N__38050,dangling_wire_245,dangling_wire_246,dangling_wire_247,N__36985,dangling_wire_248,dangling_wire_249,dangling_wire_250,N__30928,dangling_wire_251}),
            .RCLKE(),
            .RCLK(N__62003),
            .RE(N__64868),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .WE(N__34498));
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged9_physical (
            .RDATA({dangling_wire_252,dangling_wire_253,buf_data_iac_5,dangling_wire_254,dangling_wire_255,dangling_wire_256,buf_data_vac_5,dangling_wire_257,dangling_wire_258,dangling_wire_259,buf_data_iac_4,dangling_wire_260,dangling_wire_261,dangling_wire_262,buf_data_vac_4,dangling_wire_263}),
            .RADDR({dangling_wire_264,N__44421,N__42246,N__44850,N__45045,N__56316,N__43746,N__39033,N__41706,N__40107,N__53070}),
            .WADDR({dangling_wire_265,N__29862,N__29973,N__30081,N__30177,N__29118,N__29226,N__29331,N__29436,N__29544,N__29652}),
            .MASK({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281}),
            .WDATA({dangling_wire_282,dangling_wire_283,N__22165,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__22930,dangling_wire_287,dangling_wire_288,dangling_wire_289,N__21961,dangling_wire_290,dangling_wire_291,dangling_wire_292,N__21562,dangling_wire_293}),
            .RCLKE(),
            .RCLK(N__61881),
            .RE(N__64617),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .WE(N__34518));
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged4_physical (
            .RDATA({dangling_wire_294,dangling_wire_295,buf_data_iac_15,dangling_wire_296,dangling_wire_297,dangling_wire_298,buf_data_vac_15,dangling_wire_299,dangling_wire_300,dangling_wire_301,buf_data_iac_14,dangling_wire_302,dangling_wire_303,dangling_wire_304,buf_data_vac_14,dangling_wire_305}),
            .RADDR({dangling_wire_306,N__44440,N__42262,N__44866,N__45061,N__56325,N__43759,N__39049,N__41719,N__40123,N__53086}),
            .WADDR({dangling_wire_307,N__29887,N__29995,N__30103,N__30202,N__29140,N__29248,N__29353,N__29461,N__29572,N__29674}),
            .MASK({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323}),
            .WDATA({dangling_wire_324,dangling_wire_325,N__46924,dangling_wire_326,dangling_wire_327,dangling_wire_328,N__24232,dangling_wire_329,dangling_wire_330,dangling_wire_331,N__41310,dangling_wire_332,dangling_wire_333,dangling_wire_334,N__28675,dangling_wire_335}),
            .RCLKE(),
            .RCLK(N__61988),
            .RE(N__64858),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .WE(N__34503));
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged8_physical (
            .RDATA({dangling_wire_336,dangling_wire_337,buf_data_iac_7,dangling_wire_338,dangling_wire_339,dangling_wire_340,buf_data_vac_7,dangling_wire_341,dangling_wire_342,dangling_wire_343,buf_data_iac_6,dangling_wire_344,dangling_wire_345,dangling_wire_346,buf_data_vac_6,dangling_wire_347}),
            .RADDR({dangling_wire_348,N__44433,N__42258,N__44862,N__45057,N__56328,N__43758,N__39045,N__41718,N__40119,N__53082}),
            .WADDR({dangling_wire_349,N__29874,N__29985,N__30093,N__30189,N__29130,N__29238,N__29343,N__29448,N__29556,N__29664}),
            .MASK({dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .WDATA({dangling_wire_366,dangling_wire_367,N__22048,dangling_wire_368,dangling_wire_369,dangling_wire_370,N__21988,dangling_wire_371,dangling_wire_372,dangling_wire_373,N__22069,dangling_wire_374,dangling_wire_375,dangling_wire_376,N__21865,dangling_wire_377}),
            .RCLKE(),
            .RCLK(N__61859),
            .RE(N__64616),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .WE(N__34534));
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged10_physical (
            .RDATA({dangling_wire_378,dangling_wire_379,buf_data_iac_3,dangling_wire_380,dangling_wire_381,dangling_wire_382,buf_data_vac_3,dangling_wire_383,dangling_wire_384,dangling_wire_385,buf_data_iac_2,dangling_wire_386,dangling_wire_387,dangling_wire_388,buf_data_vac_2,dangling_wire_389}),
            .RADDR({dangling_wire_390,N__44464,N__42286,N__44890,N__45085,N__56350,N__43783,N__39073,N__41743,N__40147,N__53110}),
            .WADDR({dangling_wire_391,N__29911,N__30019,N__30127,N__30226,N__29164,N__29272,N__29377,N__29485,N__29596,N__29698}),
            .MASK({dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407}),
            .WDATA({dangling_wire_408,dangling_wire_409,N__33700,dangling_wire_410,dangling_wire_411,dangling_wire_412,N__33655,dangling_wire_413,dangling_wire_414,dangling_wire_415,N__36067,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__35458,dangling_wire_419}),
            .RCLKE(),
            .RCLK(N__61867),
            .RE(N__64823),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .WE(N__34535));
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged3_physical (
            .RDATA({dangling_wire_420,dangling_wire_421,buf_data_iac_17,dangling_wire_422,dangling_wire_423,dangling_wire_424,buf_data_vac_17,dangling_wire_425,dangling_wire_426,dangling_wire_427,buf_data_iac_16,dangling_wire_428,dangling_wire_429,dangling_wire_430,buf_data_vac_16,dangling_wire_431}),
            .RADDR({dangling_wire_432,N__44446,N__42268,N__44872,N__45067,N__56332,N__43765,N__39055,N__41725,N__40129,N__53092}),
            .WADDR({dangling_wire_433,N__29893,N__30001,N__30109,N__30208,N__29146,N__29254,N__29359,N__29467,N__29578,N__29680}),
            .MASK({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449}),
            .WDATA({dangling_wire_450,dangling_wire_451,N__30271,dangling_wire_452,dangling_wire_453,dangling_wire_454,N__48613,dangling_wire_455,dangling_wire_456,dangling_wire_457,N__34390,dangling_wire_458,dangling_wire_459,dangling_wire_460,N__43516,dangling_wire_461}),
            .RCLKE(),
            .RCLK(N__61959),
            .RE(N__64857),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .WE(N__34504));
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged11_physical (
            .RDATA({dangling_wire_462,dangling_wire_463,buf_data_iac_1,dangling_wire_464,dangling_wire_465,dangling_wire_466,buf_data_vac_1,dangling_wire_467,dangling_wire_468,dangling_wire_469,buf_data_iac_0,dangling_wire_470,dangling_wire_471,dangling_wire_472,buf_data_vac_0,dangling_wire_473}),
            .RADDR({dangling_wire_474,N__44458,N__42280,N__44884,N__45079,N__56344,N__43777,N__39067,N__41737,N__40141,N__53104}),
            .WADDR({dangling_wire_475,N__29905,N__30013,N__30121,N__30220,N__29158,N__29266,N__29371,N__29479,N__29590,N__29692}),
            .MASK({dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .WDATA({dangling_wire_492,dangling_wire_493,N__36094,dangling_wire_494,dangling_wire_495,dangling_wire_496,N__33610,dangling_wire_497,dangling_wire_498,dangling_wire_499,N__38098,dangling_wire_500,dangling_wire_501,dangling_wire_502,N__37882,dangling_wire_503}),
            .RCLKE(),
            .RCLK(N__61892),
            .RE(N__64828),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .WE(N__34524));
    IO_PAD ipInertedIOPad_VAC_DRDY_iopad (
            .OE(N__65921),
            .DIN(N__65920),
            .DOUT(N__65919),
            .PACKAGEPIN(VAC_DRDY));
    defparam ipInertedIOPad_VAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_DRDY_preio (
            .PADOEN(N__65921),
            .PADOUT(N__65920),
            .PADIN(N__65919),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT1_iopad (
            .OE(N__65912),
            .DIN(N__65911),
            .DOUT(N__65910),
            .PACKAGEPIN(IAC_FLT1));
    defparam ipInertedIOPad_IAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT1_preio (
            .PADOEN(N__65912),
            .PADOUT(N__65911),
            .PADIN(N__65910),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29809),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK_iopad (
            .OE(N__65903),
            .DIN(N__65902),
            .DOUT(N__65901),
            .PACKAGEPIN(DDS_SCK));
    defparam ipInertedIOPad_DDS_SCK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK_preio (
            .PADOEN(N__65903),
            .PADOUT(N__65902),
            .PADIN(N__65901),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__47614),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_166_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_166_iopad (
            .OE(N__65894),
            .DIN(N__65893),
            .DOUT(N__65892),
            .PACKAGEPIN(ICE_IOR_166));
    defparam ipInertedIOPad_ICE_IOR_166_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_166_preio (
            .PADOEN(N__65894),
            .PADOUT(N__65893),
            .PADIN(N__65892),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_119_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_119_iopad (
            .OE(N__65885),
            .DIN(N__65884),
            .DOUT(N__65883),
            .PACKAGEPIN(ICE_IOR_119));
    defparam ipInertedIOPad_ICE_IOR_119_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_119_preio (
            .PADOEN(N__65885),
            .PADOUT(N__65884),
            .PADIN(N__65883),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI_iopad (
            .OE(N__65876),
            .DIN(N__65875),
            .DOUT(N__65874),
            .PACKAGEPIN(DDS_MOSI));
    defparam ipInertedIOPad_DDS_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI_preio (
            .PADOEN(N__65876),
            .PADOUT(N__65875),
            .PADIN(N__65874),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__40024),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MISO_iopad (
            .OE(N__65867),
            .DIN(N__65866),
            .DOUT(N__65865),
            .PACKAGEPIN(VAC_MISO));
    defparam ipInertedIOPad_VAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_MISO_preio (
            .PADOEN(N__65867),
            .PADOUT(N__65866),
            .PADIN(N__65865),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI1_iopad (
            .OE(N__65858),
            .DIN(N__65857),
            .DOUT(N__65856),
            .PACKAGEPIN(DDS_MOSI1));
    defparam ipInertedIOPad_DDS_MOSI1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI1_preio (
            .PADOEN(N__65858),
            .PADOUT(N__65857),
            .PADIN(N__65856),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24289),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_146_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_146_iopad (
            .OE(N__65849),
            .DIN(N__65848),
            .DOUT(N__65847),
            .PACKAGEPIN(ICE_IOR_146));
    defparam ipInertedIOPad_ICE_IOR_146_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_146_preio (
            .PADOEN(N__65849),
            .PADOUT(N__65848),
            .PADIN(N__65847),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_CLK_iopad (
            .OE(N__65840),
            .DIN(N__65839),
            .DOUT(N__65838),
            .PACKAGEPIN(VDC_CLK));
    defparam ipInertedIOPad_VDC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_CLK_preio (
            .PADOEN(N__65840),
            .PADOUT(N__65839),
            .PADIN(N__65838),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__42760),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_222_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_222_iopad (
            .OE(N__65831),
            .DIN(N__65830),
            .DOUT(N__65829),
            .PACKAGEPIN(ICE_IOT_222));
    defparam ipInertedIOPad_ICE_IOT_222_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_222_preio (
            .PADOEN(N__65831),
            .PADOUT(N__65830),
            .PADIN(N__65829),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CS_iopad (
            .OE(N__65822),
            .DIN(N__65821),
            .DOUT(N__65820),
            .PACKAGEPIN(IAC_CS));
    defparam ipInertedIOPad_IAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CS_preio (
            .PADOEN(N__65822),
            .PADOUT(N__65821),
            .PADIN(N__65820),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25771),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_18B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_18B_iopad (
            .OE(N__65813),
            .DIN(N__65812),
            .DOUT(N__65811),
            .PACKAGEPIN(ICE_IOL_18B));
    defparam ipInertedIOPad_ICE_IOL_18B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_18B_preio (
            .PADOEN(N__65813),
            .PADOUT(N__65812),
            .PADIN(N__65811),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13A_iopad (
            .OE(N__65804),
            .DIN(N__65803),
            .DOUT(N__65802),
            .PACKAGEPIN(ICE_IOL_13A));
    defparam ipInertedIOPad_ICE_IOL_13A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13A_preio (
            .PADOEN(N__65804),
            .PADOUT(N__65803),
            .PADIN(N__65802),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_81_iopad (
            .OE(N__65795),
            .DIN(N__65794),
            .DOUT(N__65793),
            .PACKAGEPIN(ICE_IOB_81));
    defparam ipInertedIOPad_ICE_IOB_81_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_81_preio (
            .PADOEN(N__65795),
            .PADOUT(N__65794),
            .PADIN(N__65793),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR1_iopad (
            .OE(N__65786),
            .DIN(N__65785),
            .DOUT(N__65784),
            .PACKAGEPIN(VAC_OSR1));
    defparam ipInertedIOPad_VAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR1_preio (
            .PADOEN(N__65786),
            .PADOUT(N__65785),
            .PADIN(N__65784),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__38668),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MOSI_iopad (
            .OE(N__65777),
            .DIN(N__65776),
            .DOUT(N__65775),
            .PACKAGEPIN(IAC_MOSI));
    defparam ipInertedIOPad_IAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_MOSI_preio (
            .PADOEN(N__65777),
            .PADOUT(N__65776),
            .PADIN(N__65775),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS1_iopad (
            .OE(N__65768),
            .DIN(N__65767),
            .DOUT(N__65766),
            .PACKAGEPIN(DDS_CS1));
    defparam ipInertedIOPad_DDS_CS1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS1_preio (
            .PADOEN(N__65768),
            .PADOUT(N__65767),
            .PADIN(N__65766),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21658),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4B_iopad (
            .OE(N__65759),
            .DIN(N__65758),
            .DOUT(N__65757),
            .PACKAGEPIN(ICE_IOL_4B));
    defparam ipInertedIOPad_ICE_IOL_4B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4B_preio (
            .PADOEN(N__65759),
            .PADOUT(N__65758),
            .PADIN(N__65757),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_94_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_94_iopad (
            .OE(N__65750),
            .DIN(N__65749),
            .DOUT(N__65748),
            .PACKAGEPIN(ICE_IOB_94));
    defparam ipInertedIOPad_ICE_IOB_94_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_94_preio (
            .PADOEN(N__65750),
            .PADOUT(N__65749),
            .PADIN(N__65748),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CS_iopad (
            .OE(N__65741),
            .DIN(N__65740),
            .DOUT(N__65739),
            .PACKAGEPIN(VAC_CS));
    defparam ipInertedIOPad_VAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CS_preio (
            .PADOEN(N__65741),
            .PADOUT(N__65740),
            .PADIN(N__65739),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21352),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CLK_iopad (
            .OE(N__65732),
            .DIN(N__65731),
            .DOUT(N__65730),
            .PACKAGEPIN(VAC_CLK));
    defparam ipInertedIOPad_VAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CLK_preio (
            .PADOEN(N__65732),
            .PADOUT(N__65731),
            .PADIN(N__65730),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26026),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_CE0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_CE0_iopad (
            .OE(N__65723),
            .DIN(N__65722),
            .DOUT(N__65721),
            .PACKAGEPIN(ICE_SPI_CE0));
    defparam ipInertedIOPad_ICE_SPI_CE0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_CE0_preio (
            .PADOEN(N__65723),
            .PADOUT(N__65722),
            .PADIN(N__65721),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_CE0),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_167_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_167_iopad (
            .OE(N__65714),
            .DIN(N__65713),
            .DOUT(N__65712),
            .PACKAGEPIN(ICE_IOR_167));
    defparam ipInertedIOPad_ICE_IOR_167_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_167_preio (
            .PADOEN(N__65714),
            .PADOUT(N__65713),
            .PADIN(N__65712),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_118_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_118_iopad (
            .OE(N__65705),
            .DIN(N__65704),
            .DOUT(N__65703),
            .PACKAGEPIN(ICE_IOR_118));
    defparam ipInertedIOPad_ICE_IOR_118_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_118_preio (
            .PADOEN(N__65705),
            .PADOUT(N__65704),
            .PADIN(N__65703),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_SDO_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_SDO_iopad (
            .OE(N__65696),
            .DIN(N__65695),
            .DOUT(N__65694),
            .PACKAGEPIN(RTD_SDO));
    defparam ipInertedIOPad_RTD_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_SDO_preio (
            .PADOEN(N__65696),
            .PADOUT(N__65695),
            .PADIN(N__65694),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_SDO),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR0_iopad (
            .OE(N__65687),
            .DIN(N__65686),
            .DOUT(N__65685),
            .PACKAGEPIN(IAC_OSR0));
    defparam ipInertedIOPad_IAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR0_preio (
            .PADOEN(N__65687),
            .PADOUT(N__65686),
            .PADIN(N__65685),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__37087),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SCLK_iopad (
            .OE(N__65678),
            .DIN(N__65677),
            .DOUT(N__65676),
            .PACKAGEPIN(VDC_SCLK));
    defparam ipInertedIOPad_VDC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_SCLK_preio (
            .PADOEN(N__65678),
            .PADOUT(N__65677),
            .PADIN(N__65676),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24877),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT1_iopad (
            .OE(N__65669),
            .DIN(N__65668),
            .DOUT(N__65667),
            .PACKAGEPIN(VAC_FLT1));
    defparam ipInertedIOPad_VAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT1_preio (
            .PADOEN(N__65669),
            .PADOUT(N__65668),
            .PADIN(N__65667),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31618),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_MOSI_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_MOSI_iopad (
            .OE(N__65660),
            .DIN(N__65659),
            .DOUT(N__65658),
            .PACKAGEPIN(ICE_SPI_MOSI));
    defparam ipInertedIOPad_ICE_SPI_MOSI_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_MOSI_preio (
            .PADOEN(N__65660),
            .PADOUT(N__65659),
            .PADIN(N__65658),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_MOSI),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_165_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_165_iopad (
            .OE(N__65651),
            .DIN(N__65650),
            .DOUT(N__65649),
            .PACKAGEPIN(ICE_IOR_165));
    defparam ipInertedIOPad_ICE_IOR_165_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_165_preio (
            .PADOEN(N__65651),
            .PADOUT(N__65650),
            .PADIN(N__65649),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_147_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_147_iopad (
            .OE(N__65642),
            .DIN(N__65641),
            .DOUT(N__65640),
            .PACKAGEPIN(ICE_IOR_147));
    defparam ipInertedIOPad_ICE_IOR_147_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_147_preio (
            .PADOEN(N__65642),
            .PADOUT(N__65641),
            .PADIN(N__65640),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_14A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_14A_iopad (
            .OE(N__65633),
            .DIN(N__65632),
            .DOUT(N__65631),
            .PACKAGEPIN(ICE_IOL_14A));
    defparam ipInertedIOPad_ICE_IOL_14A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_14A_preio (
            .PADOEN(N__65633),
            .PADOUT(N__65632),
            .PADIN(N__65631),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13B_iopad (
            .OE(N__65624),
            .DIN(N__65623),
            .DOUT(N__65622),
            .PACKAGEPIN(ICE_IOL_13B));
    defparam ipInertedIOPad_ICE_IOL_13B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13B_preio (
            .PADOEN(N__65624),
            .PADOUT(N__65623),
            .PADIN(N__65622),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_91_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_91_iopad (
            .OE(N__65615),
            .DIN(N__65614),
            .DOUT(N__65613),
            .PACKAGEPIN(ICE_IOB_91));
    defparam ipInertedIOPad_ICE_IOB_91_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_91_preio (
            .PADOEN(N__65615),
            .PADOUT(N__65614),
            .PADIN(N__65613),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_0_iopad (
            .OE(N__65606),
            .DIN(N__65605),
            .DOUT(N__65604),
            .PACKAGEPIN(ICE_GPMO_0));
    defparam ipInertedIOPad_ICE_GPMO_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_0_preio (
            .PADOEN(N__65606),
            .PADOUT(N__65605),
            .PADIN(N__65604),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_RNG_0_iopad (
            .OE(N__65597),
            .DIN(N__65596),
            .DOUT(N__65595),
            .PACKAGEPIN(DDS_RNG_0));
    defparam ipInertedIOPad_DDS_RNG_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_RNG_0_preio (
            .PADOEN(N__65597),
            .PADOUT(N__65596),
            .PADIN(N__65595),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__49897),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_RNG0_iopad (
            .OE(N__65588),
            .DIN(N__65587),
            .DOUT(N__65586),
            .PACKAGEPIN(VDC_RNG0));
    defparam ipInertedIOPad_VDC_RNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_RNG0_preio (
            .PADOEN(N__65588),
            .PADOUT(N__65587),
            .PADIN(N__65586),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__39892),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_SCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_SCLK_iopad (
            .OE(N__65579),
            .DIN(N__65578),
            .DOUT(N__65577),
            .PACKAGEPIN(ICE_SPI_SCLK));
    defparam ipInertedIOPad_ICE_SPI_SCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_SCLK_preio (
            .PADOEN(N__65579),
            .PADOUT(N__65578),
            .PADIN(N__65577),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_SCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_152_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_152_iopad (
            .OE(N__65570),
            .DIN(N__65569),
            .DOUT(N__65568),
            .PACKAGEPIN(ICE_IOR_152));
    defparam ipInertedIOPad_ICE_IOR_152_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_152_preio (
            .PADOEN(N__65570),
            .PADOUT(N__65569),
            .PADIN(N__65568),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12A_iopad (
            .OE(N__65561),
            .DIN(N__65560),
            .DOUT(N__65559),
            .PACKAGEPIN(ICE_IOL_12A));
    defparam ipInertedIOPad_ICE_IOL_12A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12A_preio (
            .PADOEN(N__65561),
            .PADOUT(N__65560),
            .PADIN(N__65559),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_DRDY_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_DRDY_iopad (
            .OE(N__65552),
            .DIN(N__65551),
            .DOUT(N__65550),
            .PACKAGEPIN(RTD_DRDY));
    defparam ipInertedIOPad_RTD_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_DRDY_preio (
            .PADOEN(N__65552),
            .PADOUT(N__65551),
            .PADIN(N__65550),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_SPI_MISO_iopad (
            .OE(N__65543),
            .DIN(N__65542),
            .DOUT(N__65541),
            .PACKAGEPIN(ICE_SPI_MISO));
    defparam ipInertedIOPad_ICE_SPI_MISO_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_SPI_MISO_preio (
            .PADOEN(N__65543),
            .PADOUT(N__65542),
            .PADIN(N__65541),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__35257),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_177_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_177_iopad (
            .OE(N__65534),
            .DIN(N__65533),
            .DOUT(N__65532),
            .PACKAGEPIN(ICE_IOT_177));
    defparam ipInertedIOPad_ICE_IOT_177_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_177_preio (
            .PADOEN(N__65534),
            .PADOUT(N__65533),
            .PADIN(N__65532),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_141_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_141_iopad (
            .OE(N__65525),
            .DIN(N__65524),
            .DOUT(N__65523),
            .PACKAGEPIN(ICE_IOR_141));
    defparam ipInertedIOPad_ICE_IOR_141_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_141_preio (
            .PADOEN(N__65525),
            .PADOUT(N__65524),
            .PADIN(N__65523),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_80_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_80_iopad (
            .OE(N__65516),
            .DIN(N__65515),
            .DOUT(N__65514),
            .PACKAGEPIN(ICE_IOB_80));
    defparam ipInertedIOPad_ICE_IOB_80_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_80_preio (
            .PADOEN(N__65516),
            .PADOUT(N__65515),
            .PADIN(N__65514),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_102_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_102_iopad (
            .OE(N__65507),
            .DIN(N__65506),
            .DOUT(N__65505),
            .PACKAGEPIN(ICE_IOB_102));
    defparam ipInertedIOPad_ICE_IOB_102_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_102_preio (
            .PADOEN(N__65507),
            .PADOUT(N__65506),
            .PADIN(N__65505),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_2_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_2_iopad (
            .OE(N__65498),
            .DIN(N__65497),
            .DOUT(N__65496),
            .PACKAGEPIN(ICE_GPMO_2));
    defparam ipInertedIOPad_ICE_GPMO_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_2_preio (
            .PADOEN(N__65498),
            .PADOUT(N__65497),
            .PADIN(N__65496),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_2),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_GPMI_0_iopad (
            .OE(N__65489),
            .DIN(N__65488),
            .DOUT(N__65487),
            .PACKAGEPIN(ICE_GPMI_0));
    defparam ipInertedIOPad_ICE_GPMI_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_GPMI_0_preio (
            .PADOEN(N__65489),
            .PADOUT(N__65488),
            .PADIN(N__65487),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__64132),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MISO_iopad (
            .OE(N__65480),
            .DIN(N__65479),
            .DOUT(N__65478),
            .PACKAGEPIN(IAC_MISO));
    defparam ipInertedIOPad_IAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_MISO_preio (
            .PADOEN(N__65480),
            .PADOUT(N__65479),
            .PADIN(N__65478),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR0_iopad (
            .OE(N__65471),
            .DIN(N__65470),
            .DOUT(N__65469),
            .PACKAGEPIN(VAC_OSR0));
    defparam ipInertedIOPad_VAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR0_preio (
            .PADOEN(N__65471),
            .PADOUT(N__65470),
            .PADIN(N__65469),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__38803),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MOSI_iopad (
            .OE(N__65462),
            .DIN(N__65461),
            .DOUT(N__65460),
            .PACKAGEPIN(VAC_MOSI));
    defparam ipInertedIOPad_VAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_MOSI_preio (
            .PADOEN(N__65462),
            .PADOUT(N__65461),
            .PADIN(N__65460),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TEST_LED_iopad (
            .OE(N__65453),
            .DIN(N__65452),
            .DOUT(N__65451),
            .PACKAGEPIN(TEST_LED));
    defparam ipInertedIOPad_TEST_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_TEST_LED_preio (
            .PADOEN(N__65453),
            .PADOUT(N__65452),
            .PADIN(N__65451),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__42808),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_148_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_148_iopad (
            .OE(N__65444),
            .DIN(N__65443),
            .DOUT(N__65442),
            .PACKAGEPIN(ICE_IOR_148));
    defparam ipInertedIOPad_ICE_IOR_148_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_148_preio (
            .PADOEN(N__65444),
            .PADOUT(N__65443),
            .PADIN(N__65442),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_STAT_COMM_iopad (
            .OE(N__65435),
            .DIN(N__65434),
            .DOUT(N__65433),
            .PACKAGEPIN(STAT_COMM));
    defparam ipInertedIOPad_STAT_COMM_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_STAT_COMM_preio (
            .PADOEN(N__65435),
            .PADOUT(N__65434),
            .PADIN(N__65433),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21241),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SYSCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SYSCLK_iopad (
            .OE(N__65426),
            .DIN(N__65425),
            .DOUT(N__65424),
            .PACKAGEPIN(ICE_SYSCLK));
    defparam ipInertedIOPad_ICE_SYSCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SYSCLK_preio (
            .PADOEN(N__65426),
            .PADOUT(N__65425),
            .PADIN(N__65424),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SYSCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_161_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_161_iopad (
            .OE(N__65417),
            .DIN(N__65416),
            .DOUT(N__65415),
            .PACKAGEPIN(ICE_IOR_161));
    defparam ipInertedIOPad_ICE_IOR_161_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_161_preio (
            .PADOEN(N__65417),
            .PADOUT(N__65416),
            .PADIN(N__65415),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_95_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_95_iopad (
            .OE(N__65408),
            .DIN(N__65407),
            .DOUT(N__65406),
            .PACKAGEPIN(ICE_IOB_95));
    defparam ipInertedIOPad_ICE_IOB_95_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_95_preio (
            .PADOEN(N__65408),
            .PADOUT(N__65407),
            .PADIN(N__65406),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_82_iopad (
            .OE(N__65399),
            .DIN(N__65398),
            .DOUT(N__65397),
            .PACKAGEPIN(ICE_IOB_82));
    defparam ipInertedIOPad_ICE_IOB_82_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_82_preio (
            .PADOEN(N__65399),
            .PADOUT(N__65398),
            .PADIN(N__65397),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_104_iopad (
            .OE(N__65390),
            .DIN(N__65389),
            .DOUT(N__65388),
            .PACKAGEPIN(ICE_IOB_104));
    defparam ipInertedIOPad_ICE_IOB_104_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_104_preio (
            .PADOEN(N__65390),
            .PADOUT(N__65389),
            .PADIN(N__65388),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CLK_iopad (
            .OE(N__65381),
            .DIN(N__65380),
            .DOUT(N__65379),
            .PACKAGEPIN(IAC_CLK));
    defparam ipInertedIOPad_IAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CLK_preio (
            .PADOEN(N__65381),
            .PADOUT(N__65380),
            .PADIN(N__65379),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26025),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS_iopad (
            .OE(N__65372),
            .DIN(N__65371),
            .DOUT(N__65370),
            .PACKAGEPIN(DDS_CS));
    defparam ipInertedIOPad_DDS_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS_preio (
            .PADOEN(N__65372),
            .PADOUT(N__65371),
            .PADIN(N__65370),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__50263),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG0_iopad (
            .OE(N__65363),
            .DIN(N__65362),
            .DOUT(N__65361),
            .PACKAGEPIN(SELIRNG0));
    defparam ipInertedIOPad_SELIRNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG0_preio (
            .PADOEN(N__65363),
            .PADOUT(N__65362),
            .PADIN(N__65361),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__39943),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SDI_iopad (
            .OE(N__65354),
            .DIN(N__65353),
            .DOUT(N__65352),
            .PACKAGEPIN(RTD_SDI));
    defparam ipInertedIOPad_RTD_SDI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SDI_preio (
            .PADOEN(N__65354),
            .PADOUT(N__65353),
            .PADIN(N__65352),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21280),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_221_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_221_iopad (
            .OE(N__65345),
            .DIN(N__65344),
            .DOUT(N__65343),
            .PACKAGEPIN(ICE_IOT_221));
    defparam ipInertedIOPad_ICE_IOT_221_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_221_preio (
            .PADOEN(N__65345),
            .PADOUT(N__65344),
            .PADIN(N__65343),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_197_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_197_iopad (
            .OE(N__65336),
            .DIN(N__65335),
            .DOUT(N__65334),
            .PACKAGEPIN(ICE_IOT_197));
    defparam ipInertedIOPad_ICE_IOT_197_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_197_preio (
            .PADOEN(N__65336),
            .PADOUT(N__65335),
            .PADIN(N__65334),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK_iopad (
            .OE(N__65327),
            .DIN(N__65326),
            .DOUT(N__65325),
            .PACKAGEPIN(DDS_MCLK));
    defparam ipInertedIOPad_DDS_MCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK_preio (
            .PADOEN(N__65327),
            .PADOUT(N__65326),
            .PADIN(N__65325),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__53380),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SCLK_iopad (
            .OE(N__65318),
            .DIN(N__65317),
            .DOUT(N__65316),
            .PACKAGEPIN(RTD_SCLK));
    defparam ipInertedIOPad_RTD_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SCLK_preio (
            .PADOEN(N__65318),
            .PADOUT(N__65317),
            .PADIN(N__65316),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21304),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_CS_iopad (
            .OE(N__65309),
            .DIN(N__65308),
            .DOUT(N__65307),
            .PACKAGEPIN(RTD_CS));
    defparam ipInertedIOPad_RTD_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_CS_preio (
            .PADOEN(N__65309),
            .PADOUT(N__65308),
            .PADIN(N__65307),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22243),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_137_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_137_iopad (
            .OE(N__65300),
            .DIN(N__65299),
            .DOUT(N__65298),
            .PACKAGEPIN(ICE_IOR_137));
    defparam ipInertedIOPad_ICE_IOR_137_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_137_preio (
            .PADOEN(N__65300),
            .PADOUT(N__65299),
            .PADIN(N__65298),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR1_iopad (
            .OE(N__65291),
            .DIN(N__65290),
            .DOUT(N__65289),
            .PACKAGEPIN(IAC_OSR1));
    defparam ipInertedIOPad_IAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR1_preio (
            .PADOEN(N__65291),
            .PADOUT(N__65290),
            .PADIN(N__65289),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__37054),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT0_iopad (
            .OE(N__65282),
            .DIN(N__65281),
            .DOUT(N__65280),
            .PACKAGEPIN(VAC_FLT0));
    defparam ipInertedIOPad_VAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT0_preio (
            .PADOEN(N__65282),
            .PADOUT(N__65281),
            .PADIN(N__65280),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31654),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_144_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_144_iopad (
            .OE(N__65273),
            .DIN(N__65272),
            .DOUT(N__65271),
            .PACKAGEPIN(ICE_IOR_144));
    defparam ipInertedIOPad_ICE_IOR_144_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_144_preio (
            .PADOEN(N__65273),
            .PADOUT(N__65272),
            .PADIN(N__65271),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_128_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_128_iopad (
            .OE(N__65264),
            .DIN(N__65263),
            .DOUT(N__65262),
            .PACKAGEPIN(ICE_IOR_128));
    defparam ipInertedIOPad_ICE_IOR_128_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_128_preio (
            .PADOEN(N__65264),
            .PADOUT(N__65263),
            .PADIN(N__65262),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_1_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_1_iopad (
            .OE(N__65255),
            .DIN(N__65254),
            .DOUT(N__65253),
            .PACKAGEPIN(ICE_GPMO_1));
    defparam ipInertedIOPad_ICE_GPMO_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_1_preio (
            .PADOEN(N__65255),
            .PADOUT(N__65254),
            .PADIN(N__65253),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_SCLK_iopad (
            .OE(N__65246),
            .DIN(N__65245),
            .DOUT(N__65244),
            .PACKAGEPIN(IAC_SCLK));
    defparam ipInertedIOPad_IAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_SCLK_preio (
            .PADOEN(N__65246),
            .PADOUT(N__65245),
            .PADIN(N__65244),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27889),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_EIS_SYNCCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_EIS_SYNCCLK_iopad (
            .OE(N__65237),
            .DIN(N__65236),
            .DOUT(N__65235),
            .PACKAGEPIN(EIS_SYNCCLK));
    defparam ipInertedIOPad_EIS_SYNCCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_EIS_SYNCCLK_preio (
            .PADOEN(N__65237),
            .PADOUT(N__65236),
            .PADIN(N__65235),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(EIS_SYNCCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_139_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_139_iopad (
            .OE(N__65228),
            .DIN(N__65227),
            .DOUT(N__65226),
            .PACKAGEPIN(ICE_IOR_139));
    defparam ipInertedIOPad_ICE_IOR_139_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_139_preio (
            .PADOEN(N__65228),
            .PADOUT(N__65227),
            .PADIN(N__65226),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4A_iopad (
            .OE(N__65219),
            .DIN(N__65218),
            .DOUT(N__65217),
            .PACKAGEPIN(ICE_IOL_4A));
    defparam ipInertedIOPad_ICE_IOL_4A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4A_preio (
            .PADOEN(N__65219),
            .PADOUT(N__65218),
            .PADIN(N__65217),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_SCLK_iopad (
            .OE(N__65210),
            .DIN(N__65209),
            .DOUT(N__65208),
            .PACKAGEPIN(VAC_SCLK));
    defparam ipInertedIOPad_VAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_SCLK_preio (
            .PADOEN(N__65210),
            .PADOUT(N__65209),
            .PADIN(N__65208),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21382),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_THERMOSTAT_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_THERMOSTAT_iopad (
            .OE(N__65201),
            .DIN(N__65200),
            .DOUT(N__65199),
            .PACKAGEPIN(THERMOSTAT));
    defparam ipInertedIOPad_THERMOSTAT_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_THERMOSTAT_preio (
            .PADOEN(N__65201),
            .PADOUT(N__65200),
            .PADIN(N__65199),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(THERMOSTAT),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_164_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_164_iopad (
            .OE(N__65192),
            .DIN(N__65191),
            .DOUT(N__65190),
            .PACKAGEPIN(ICE_IOR_164));
    defparam ipInertedIOPad_ICE_IOR_164_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_164_preio (
            .PADOEN(N__65192),
            .PADOUT(N__65191),
            .PADIN(N__65190),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_103_iopad (
            .OE(N__65183),
            .DIN(N__65182),
            .DOUT(N__65181),
            .PACKAGEPIN(ICE_IOB_103));
    defparam ipInertedIOPad_ICE_IOB_103_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_103_preio (
            .PADOEN(N__65183),
            .PADOUT(N__65182),
            .PADIN(N__65181),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AMPV_POW_iopad (
            .OE(N__65174),
            .DIN(N__65173),
            .DOUT(N__65172),
            .PACKAGEPIN(AMPV_POW));
    defparam ipInertedIOPad_AMPV_POW_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AMPV_POW_preio (
            .PADOEN(N__65174),
            .PADOUT(N__65173),
            .PADIN(N__65172),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36514),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SDO_iopad (
            .OE(N__65165),
            .DIN(N__65164),
            .DOUT(N__65163),
            .PACKAGEPIN(VDC_SDO));
    defparam ipInertedIOPad_VDC_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDC_SDO_preio (
            .PADOEN(N__65165),
            .PADOUT(N__65164),
            .PADIN(N__65163),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VDC_SDO),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_174_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_174_iopad (
            .OE(N__65156),
            .DIN(N__65155),
            .DOUT(N__65154),
            .PACKAGEPIN(ICE_IOT_174));
    defparam ipInertedIOPad_ICE_IOT_174_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_174_preio (
            .PADOEN(N__65156),
            .PADOUT(N__65155),
            .PADIN(N__65154),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_140_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_140_iopad (
            .OE(N__65147),
            .DIN(N__65146),
            .DOUT(N__65145),
            .PACKAGEPIN(ICE_IOR_140));
    defparam ipInertedIOPad_ICE_IOR_140_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_140_preio (
            .PADOEN(N__65147),
            .PADOUT(N__65146),
            .PADIN(N__65145),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_96_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_96_iopad (
            .OE(N__65138),
            .DIN(N__65137),
            .DOUT(N__65136),
            .PACKAGEPIN(ICE_IOB_96));
    defparam ipInertedIOPad_ICE_IOB_96_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_96_preio (
            .PADOEN(N__65138),
            .PADOUT(N__65137),
            .PADIN(N__65136),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_CONT_SD_iopad (
            .OE(N__65129),
            .DIN(N__65128),
            .DOUT(N__65127),
            .PACKAGEPIN(CONT_SD));
    defparam ipInertedIOPad_CONT_SD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_CONT_SD_preio (
            .PADOEN(N__65129),
            .PADOUT(N__65128),
            .PADIN(N__65127),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__52606),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AC_ADC_SYNC_iopad (
            .OE(N__65120),
            .DIN(N__65119),
            .DOUT(N__65118),
            .PACKAGEPIN(AC_ADC_SYNC));
    defparam ipInertedIOPad_AC_ADC_SYNC_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AC_ADC_SYNC_preio (
            .PADOEN(N__65120),
            .PADOUT(N__65119),
            .PADIN(N__65118),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23071),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG1_iopad (
            .OE(N__65111),
            .DIN(N__65110),
            .DOUT(N__65109),
            .PACKAGEPIN(SELIRNG1));
    defparam ipInertedIOPad_SELIRNG1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG1_preio (
            .PADOEN(N__65111),
            .PADOUT(N__65110),
            .PADIN(N__65109),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__52780),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12B_iopad (
            .OE(N__65102),
            .DIN(N__65101),
            .DOUT(N__65100),
            .PACKAGEPIN(ICE_IOL_12B));
    defparam ipInertedIOPad_ICE_IOL_12B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12B_preio (
            .PADOEN(N__65102),
            .PADOUT(N__65101),
            .PADIN(N__65100),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_160_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_160_iopad (
            .OE(N__65093),
            .DIN(N__65092),
            .DOUT(N__65091),
            .PACKAGEPIN(ICE_IOR_160));
    defparam ipInertedIOPad_ICE_IOR_160_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_160_preio (
            .PADOEN(N__65093),
            .PADOUT(N__65092),
            .PADIN(N__65091),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_136_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_136_iopad (
            .OE(N__65084),
            .DIN(N__65083),
            .DOUT(N__65082),
            .PACKAGEPIN(ICE_IOR_136));
    defparam ipInertedIOPad_ICE_IOR_136_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_136_preio (
            .PADOEN(N__65084),
            .PADOUT(N__65083),
            .PADIN(N__65082),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK1_iopad (
            .OE(N__65075),
            .DIN(N__65074),
            .DOUT(N__65073),
            .PACKAGEPIN(DDS_MCLK1));
    defparam ipInertedIOPad_DDS_MCLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK1_preio (
            .PADOEN(N__65075),
            .PADOUT(N__65074),
            .PADIN(N__65073),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24829),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_198_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_198_iopad (
            .OE(N__65066),
            .DIN(N__65065),
            .DOUT(N__65064),
            .PACKAGEPIN(ICE_IOT_198));
    defparam ipInertedIOPad_ICE_IOT_198_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_198_preio (
            .PADOEN(N__65066),
            .PADOUT(N__65065),
            .PADIN(N__65064),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_173_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_173_iopad (
            .OE(N__65057),
            .DIN(N__65056),
            .DOUT(N__65055),
            .PACKAGEPIN(ICE_IOT_173));
    defparam ipInertedIOPad_ICE_IOT_173_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_173_preio (
            .PADOEN(N__65057),
            .PADOUT(N__65056),
            .PADIN(N__65055),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_DRDY_iopad (
            .OE(N__65048),
            .DIN(N__65047),
            .DOUT(N__65046),
            .PACKAGEPIN(IAC_DRDY));
    defparam ipInertedIOPad_IAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_DRDY_preio (
            .PADOEN(N__65048),
            .PADOUT(N__65047),
            .PADIN(N__65046),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_DRDY),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_178_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_178_iopad (
            .OE(N__65039),
            .DIN(N__65038),
            .DOUT(N__65037),
            .PACKAGEPIN(ICE_IOT_178));
    defparam ipInertedIOPad_ICE_IOT_178_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_178_preio (
            .PADOEN(N__65039),
            .PADOUT(N__65038),
            .PADIN(N__65037),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_138_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_138_iopad (
            .OE(N__65030),
            .DIN(N__65029),
            .DOUT(N__65028),
            .PACKAGEPIN(ICE_IOR_138));
    defparam ipInertedIOPad_ICE_IOR_138_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_138_preio (
            .PADOEN(N__65030),
            .PADOUT(N__65029),
            .PADIN(N__65028),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_120_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_120_iopad (
            .OE(N__65021),
            .DIN(N__65020),
            .DOUT(N__65019),
            .PACKAGEPIN(ICE_IOR_120));
    defparam ipInertedIOPad_ICE_IOR_120_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_120_preio (
            .PADOEN(N__65021),
            .PADOUT(N__65020),
            .PADIN(N__65019),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT0_iopad (
            .OE(N__65012),
            .DIN(N__65011),
            .DOUT(N__65010),
            .PACKAGEPIN(IAC_FLT0));
    defparam ipInertedIOPad_IAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT0_preio (
            .PADOEN(N__65012),
            .PADOUT(N__65011),
            .PADIN(N__65010),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30574),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK1_iopad (
            .OE(N__65003),
            .DIN(N__65002),
            .DOUT(N__65001),
            .PACKAGEPIN(DDS_SCK1));
    defparam ipInertedIOPad_DDS_SCK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK1_preio (
            .PADOEN(N__65003),
            .PADOUT(N__65002),
            .PADIN(N__65001),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21331),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    CascadeMux I__16328 (
            .O(N__64984),
            .I(N__64981));
    InMux I__16327 (
            .O(N__64981),
            .I(N__64977));
    InMux I__16326 (
            .O(N__64980),
            .I(N__64974));
    LocalMux I__16325 (
            .O(N__64977),
            .I(N__64971));
    LocalMux I__16324 (
            .O(N__64974),
            .I(\ADC_VDC.genclk.t0off_8 ));
    Odrv4 I__16323 (
            .O(N__64971),
            .I(\ADC_VDC.genclk.t0off_8 ));
    InMux I__16322 (
            .O(N__64966),
            .I(bfn_23_6_0_));
    InMux I__16321 (
            .O(N__64963),
            .I(N__64959));
    InMux I__16320 (
            .O(N__64962),
            .I(N__64956));
    LocalMux I__16319 (
            .O(N__64959),
            .I(\ADC_VDC.genclk.t0off_9 ));
    LocalMux I__16318 (
            .O(N__64956),
            .I(\ADC_VDC.genclk.t0off_9 ));
    InMux I__16317 (
            .O(N__64951),
            .I(\ADC_VDC.genclk.n20744 ));
    InMux I__16316 (
            .O(N__64948),
            .I(N__64944));
    InMux I__16315 (
            .O(N__64947),
            .I(N__64941));
    LocalMux I__16314 (
            .O(N__64944),
            .I(\ADC_VDC.genclk.t0off_10 ));
    LocalMux I__16313 (
            .O(N__64941),
            .I(\ADC_VDC.genclk.t0off_10 ));
    InMux I__16312 (
            .O(N__64936),
            .I(\ADC_VDC.genclk.n20745 ));
    InMux I__16311 (
            .O(N__64933),
            .I(N__64929));
    InMux I__16310 (
            .O(N__64932),
            .I(N__64926));
    LocalMux I__16309 (
            .O(N__64929),
            .I(\ADC_VDC.genclk.t0off_11 ));
    LocalMux I__16308 (
            .O(N__64926),
            .I(\ADC_VDC.genclk.t0off_11 ));
    InMux I__16307 (
            .O(N__64921),
            .I(\ADC_VDC.genclk.n20746 ));
    InMux I__16306 (
            .O(N__64918),
            .I(N__64914));
    InMux I__16305 (
            .O(N__64917),
            .I(N__64911));
    LocalMux I__16304 (
            .O(N__64914),
            .I(\ADC_VDC.genclk.t0off_12 ));
    LocalMux I__16303 (
            .O(N__64911),
            .I(\ADC_VDC.genclk.t0off_12 ));
    InMux I__16302 (
            .O(N__64906),
            .I(\ADC_VDC.genclk.n20747 ));
    InMux I__16301 (
            .O(N__64903),
            .I(N__64899));
    InMux I__16300 (
            .O(N__64902),
            .I(N__64896));
    LocalMux I__16299 (
            .O(N__64899),
            .I(\ADC_VDC.genclk.t0off_13 ));
    LocalMux I__16298 (
            .O(N__64896),
            .I(\ADC_VDC.genclk.t0off_13 ));
    InMux I__16297 (
            .O(N__64891),
            .I(\ADC_VDC.genclk.n20748 ));
    InMux I__16296 (
            .O(N__64888),
            .I(N__64884));
    InMux I__16295 (
            .O(N__64887),
            .I(N__64881));
    LocalMux I__16294 (
            .O(N__64884),
            .I(\ADC_VDC.genclk.t0off_14 ));
    LocalMux I__16293 (
            .O(N__64881),
            .I(\ADC_VDC.genclk.t0off_14 ));
    InMux I__16292 (
            .O(N__64876),
            .I(\ADC_VDC.genclk.n20749 ));
    SRMux I__16291 (
            .O(N__64873),
            .I(N__64870));
    LocalMux I__16290 (
            .O(N__64870),
            .I(N__64865));
    SRMux I__16289 (
            .O(N__64869),
            .I(N__64862));
    SRMux I__16288 (
            .O(N__64868),
            .I(N__64859));
    Span4Mux_v I__16287 (
            .O(N__64865),
            .I(N__64841));
    LocalMux I__16286 (
            .O(N__64862),
            .I(N__64836));
    LocalMux I__16285 (
            .O(N__64859),
            .I(N__64836));
    SRMux I__16284 (
            .O(N__64858),
            .I(N__64833));
    SRMux I__16283 (
            .O(N__64857),
            .I(N__64830));
    SRMux I__16282 (
            .O(N__64856),
            .I(N__64825));
    IoInMux I__16281 (
            .O(N__64855),
            .I(N__64820));
    CascadeMux I__16280 (
            .O(N__64854),
            .I(N__64816));
    CascadeMux I__16279 (
            .O(N__64853),
            .I(N__64812));
    CascadeMux I__16278 (
            .O(N__64852),
            .I(N__64808));
    CascadeMux I__16277 (
            .O(N__64851),
            .I(N__64804));
    CascadeMux I__16276 (
            .O(N__64850),
            .I(N__64800));
    CascadeMux I__16275 (
            .O(N__64849),
            .I(N__64796));
    CascadeMux I__16274 (
            .O(N__64848),
            .I(N__64792));
    CascadeMux I__16273 (
            .O(N__64847),
            .I(N__64789));
    CascadeMux I__16272 (
            .O(N__64846),
            .I(N__64785));
    CascadeMux I__16271 (
            .O(N__64845),
            .I(N__64781));
    CascadeMux I__16270 (
            .O(N__64844),
            .I(N__64777));
    Span4Mux_v I__16269 (
            .O(N__64841),
            .I(N__64774));
    Span4Mux_v I__16268 (
            .O(N__64836),
            .I(N__64767));
    LocalMux I__16267 (
            .O(N__64833),
            .I(N__64767));
    LocalMux I__16266 (
            .O(N__64830),
            .I(N__64767));
    SRMux I__16265 (
            .O(N__64829),
            .I(N__64764));
    SRMux I__16264 (
            .O(N__64828),
            .I(N__64761));
    LocalMux I__16263 (
            .O(N__64825),
            .I(N__64758));
    SRMux I__16262 (
            .O(N__64824),
            .I(N__64755));
    SRMux I__16261 (
            .O(N__64823),
            .I(N__64752));
    LocalMux I__16260 (
            .O(N__64820),
            .I(N__64749));
    InMux I__16259 (
            .O(N__64819),
            .I(N__64734));
    InMux I__16258 (
            .O(N__64816),
            .I(N__64734));
    InMux I__16257 (
            .O(N__64815),
            .I(N__64734));
    InMux I__16256 (
            .O(N__64812),
            .I(N__64734));
    InMux I__16255 (
            .O(N__64811),
            .I(N__64734));
    InMux I__16254 (
            .O(N__64808),
            .I(N__64734));
    InMux I__16253 (
            .O(N__64807),
            .I(N__64734));
    InMux I__16252 (
            .O(N__64804),
            .I(N__64712));
    InMux I__16251 (
            .O(N__64803),
            .I(N__64712));
    InMux I__16250 (
            .O(N__64800),
            .I(N__64712));
    InMux I__16249 (
            .O(N__64799),
            .I(N__64712));
    InMux I__16248 (
            .O(N__64796),
            .I(N__64712));
    InMux I__16247 (
            .O(N__64795),
            .I(N__64712));
    InMux I__16246 (
            .O(N__64792),
            .I(N__64712));
    InMux I__16245 (
            .O(N__64789),
            .I(N__64697));
    InMux I__16244 (
            .O(N__64788),
            .I(N__64697));
    InMux I__16243 (
            .O(N__64785),
            .I(N__64697));
    InMux I__16242 (
            .O(N__64784),
            .I(N__64697));
    InMux I__16241 (
            .O(N__64781),
            .I(N__64697));
    InMux I__16240 (
            .O(N__64780),
            .I(N__64697));
    InMux I__16239 (
            .O(N__64777),
            .I(N__64697));
    Span4Mux_v I__16238 (
            .O(N__64774),
            .I(N__64684));
    Span4Mux_v I__16237 (
            .O(N__64767),
            .I(N__64684));
    LocalMux I__16236 (
            .O(N__64764),
            .I(N__64684));
    LocalMux I__16235 (
            .O(N__64761),
            .I(N__64684));
    Span4Mux_v I__16234 (
            .O(N__64758),
            .I(N__64677));
    LocalMux I__16233 (
            .O(N__64755),
            .I(N__64677));
    LocalMux I__16232 (
            .O(N__64752),
            .I(N__64677));
    Span4Mux_s3_v I__16231 (
            .O(N__64749),
            .I(N__64673));
    LocalMux I__16230 (
            .O(N__64734),
            .I(N__64670));
    CascadeMux I__16229 (
            .O(N__64733),
            .I(N__64667));
    CascadeMux I__16228 (
            .O(N__64732),
            .I(N__64663));
    CascadeMux I__16227 (
            .O(N__64731),
            .I(N__64660));
    CascadeMux I__16226 (
            .O(N__64730),
            .I(N__64657));
    CascadeMux I__16225 (
            .O(N__64729),
            .I(N__64654));
    CascadeMux I__16224 (
            .O(N__64728),
            .I(N__64651));
    CascadeMux I__16223 (
            .O(N__64727),
            .I(N__64648));
    LocalMux I__16222 (
            .O(N__64712),
            .I(N__64645));
    LocalMux I__16221 (
            .O(N__64697),
            .I(N__64642));
    CascadeMux I__16220 (
            .O(N__64696),
            .I(N__64638));
    CascadeMux I__16219 (
            .O(N__64695),
            .I(N__64634));
    CascadeMux I__16218 (
            .O(N__64694),
            .I(N__64630));
    CascadeMux I__16217 (
            .O(N__64693),
            .I(N__64626));
    Span4Mux_v I__16216 (
            .O(N__64684),
            .I(N__64621));
    Span4Mux_v I__16215 (
            .O(N__64677),
            .I(N__64621));
    InMux I__16214 (
            .O(N__64676),
            .I(N__64618));
    Span4Mux_v I__16213 (
            .O(N__64673),
            .I(N__64613));
    Span4Mux_h I__16212 (
            .O(N__64670),
            .I(N__64610));
    InMux I__16211 (
            .O(N__64667),
            .I(N__64601));
    InMux I__16210 (
            .O(N__64666),
            .I(N__64601));
    InMux I__16209 (
            .O(N__64663),
            .I(N__64601));
    InMux I__16208 (
            .O(N__64660),
            .I(N__64601));
    InMux I__16207 (
            .O(N__64657),
            .I(N__64592));
    InMux I__16206 (
            .O(N__64654),
            .I(N__64592));
    InMux I__16205 (
            .O(N__64651),
            .I(N__64592));
    InMux I__16204 (
            .O(N__64648),
            .I(N__64592));
    Span4Mux_v I__16203 (
            .O(N__64645),
            .I(N__64587));
    Span4Mux_v I__16202 (
            .O(N__64642),
            .I(N__64587));
    InMux I__16201 (
            .O(N__64641),
            .I(N__64570));
    InMux I__16200 (
            .O(N__64638),
            .I(N__64570));
    InMux I__16199 (
            .O(N__64637),
            .I(N__64570));
    InMux I__16198 (
            .O(N__64634),
            .I(N__64570));
    InMux I__16197 (
            .O(N__64633),
            .I(N__64570));
    InMux I__16196 (
            .O(N__64630),
            .I(N__64570));
    InMux I__16195 (
            .O(N__64629),
            .I(N__64570));
    InMux I__16194 (
            .O(N__64626),
            .I(N__64570));
    Span4Mux_h I__16193 (
            .O(N__64621),
            .I(N__64567));
    LocalMux I__16192 (
            .O(N__64618),
            .I(N__64564));
    SRMux I__16191 (
            .O(N__64617),
            .I(N__64561));
    SRMux I__16190 (
            .O(N__64616),
            .I(N__64558));
    Span4Mux_v I__16189 (
            .O(N__64613),
            .I(N__64554));
    Sp12to4 I__16188 (
            .O(N__64610),
            .I(N__64551));
    LocalMux I__16187 (
            .O(N__64601),
            .I(N__64542));
    LocalMux I__16186 (
            .O(N__64592),
            .I(N__64542));
    Sp12to4 I__16185 (
            .O(N__64587),
            .I(N__64542));
    LocalMux I__16184 (
            .O(N__64570),
            .I(N__64542));
    Span4Mux_h I__16183 (
            .O(N__64567),
            .I(N__64537));
    Span4Mux_v I__16182 (
            .O(N__64564),
            .I(N__64537));
    LocalMux I__16181 (
            .O(N__64561),
            .I(N__64534));
    LocalMux I__16180 (
            .O(N__64558),
            .I(N__64531));
    InMux I__16179 (
            .O(N__64557),
            .I(N__64528));
    Sp12to4 I__16178 (
            .O(N__64554),
            .I(N__64521));
    Span12Mux_v I__16177 (
            .O(N__64551),
            .I(N__64521));
    Span12Mux_h I__16176 (
            .O(N__64542),
            .I(N__64521));
    Span4Mux_h I__16175 (
            .O(N__64537),
            .I(N__64518));
    Span4Mux_v I__16174 (
            .O(N__64534),
            .I(N__64513));
    Span4Mux_v I__16173 (
            .O(N__64531),
            .I(N__64513));
    LocalMux I__16172 (
            .O(N__64528),
            .I(N__64510));
    Odrv12 I__16171 (
            .O(N__64521),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__16170 (
            .O(N__64518),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__16169 (
            .O(N__64513),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__16168 (
            .O(N__64510),
            .I(CONSTANT_ONE_NET));
    InMux I__16167 (
            .O(N__64501),
            .I(\ADC_VDC.genclk.n20750 ));
    CascadeMux I__16166 (
            .O(N__64498),
            .I(N__64494));
    InMux I__16165 (
            .O(N__64497),
            .I(N__64491));
    InMux I__16164 (
            .O(N__64494),
            .I(N__64488));
    LocalMux I__16163 (
            .O(N__64491),
            .I(\ADC_VDC.genclk.t0off_15 ));
    LocalMux I__16162 (
            .O(N__64488),
            .I(\ADC_VDC.genclk.t0off_15 ));
    CEMux I__16161 (
            .O(N__64483),
            .I(N__64480));
    LocalMux I__16160 (
            .O(N__64480),
            .I(N__64476));
    CEMux I__16159 (
            .O(N__64479),
            .I(N__64473));
    Span4Mux_v I__16158 (
            .O(N__64476),
            .I(N__64470));
    LocalMux I__16157 (
            .O(N__64473),
            .I(N__64467));
    Span4Mux_h I__16156 (
            .O(N__64470),
            .I(N__64462));
    Span4Mux_h I__16155 (
            .O(N__64467),
            .I(N__64462));
    Odrv4 I__16154 (
            .O(N__64462),
            .I(\ADC_VDC.genclk.n12361 ));
    SRMux I__16153 (
            .O(N__64459),
            .I(N__64454));
    SRMux I__16152 (
            .O(N__64458),
            .I(N__64451));
    SRMux I__16151 (
            .O(N__64457),
            .I(N__64448));
    LocalMux I__16150 (
            .O(N__64454),
            .I(N__64444));
    LocalMux I__16149 (
            .O(N__64451),
            .I(N__64441));
    LocalMux I__16148 (
            .O(N__64448),
            .I(N__64438));
    SRMux I__16147 (
            .O(N__64447),
            .I(N__64435));
    Span4Mux_h I__16146 (
            .O(N__64444),
            .I(N__64432));
    Span4Mux_h I__16145 (
            .O(N__64441),
            .I(N__64427));
    Span4Mux_h I__16144 (
            .O(N__64438),
            .I(N__64427));
    LocalMux I__16143 (
            .O(N__64435),
            .I(N__64424));
    Odrv4 I__16142 (
            .O(N__64432),
            .I(\ADC_VDC.genclk.n15418 ));
    Odrv4 I__16141 (
            .O(N__64427),
            .I(\ADC_VDC.genclk.n15418 ));
    Odrv4 I__16140 (
            .O(N__64424),
            .I(\ADC_VDC.genclk.n15418 ));
    SRMux I__16139 (
            .O(N__64417),
            .I(N__64413));
    SRMux I__16138 (
            .O(N__64416),
            .I(N__64410));
    LocalMux I__16137 (
            .O(N__64413),
            .I(N__64407));
    LocalMux I__16136 (
            .O(N__64410),
            .I(N__64404));
    Span4Mux_h I__16135 (
            .O(N__64407),
            .I(N__64401));
    Span4Mux_h I__16134 (
            .O(N__64404),
            .I(N__64398));
    Odrv4 I__16133 (
            .O(N__64401),
            .I(n15482));
    Odrv4 I__16132 (
            .O(N__64398),
            .I(n15482));
    InMux I__16131 (
            .O(N__64393),
            .I(N__64389));
    InMux I__16130 (
            .O(N__64392),
            .I(N__64386));
    LocalMux I__16129 (
            .O(N__64389),
            .I(\ADC_VDC.genclk.t0off_0 ));
    LocalMux I__16128 (
            .O(N__64386),
            .I(\ADC_VDC.genclk.t0off_0 ));
    InMux I__16127 (
            .O(N__64381),
            .I(bfn_23_5_0_));
    InMux I__16126 (
            .O(N__64378),
            .I(N__64374));
    InMux I__16125 (
            .O(N__64377),
            .I(N__64371));
    LocalMux I__16124 (
            .O(N__64374),
            .I(\ADC_VDC.genclk.t0off_1 ));
    LocalMux I__16123 (
            .O(N__64371),
            .I(\ADC_VDC.genclk.t0off_1 ));
    InMux I__16122 (
            .O(N__64366),
            .I(\ADC_VDC.genclk.n20736 ));
    CascadeMux I__16121 (
            .O(N__64363),
            .I(N__64360));
    InMux I__16120 (
            .O(N__64360),
            .I(N__64356));
    InMux I__16119 (
            .O(N__64359),
            .I(N__64353));
    LocalMux I__16118 (
            .O(N__64356),
            .I(N__64348));
    LocalMux I__16117 (
            .O(N__64353),
            .I(N__64348));
    Odrv4 I__16116 (
            .O(N__64348),
            .I(\ADC_VDC.genclk.t0off_2 ));
    InMux I__16115 (
            .O(N__64345),
            .I(\ADC_VDC.genclk.n20737 ));
    InMux I__16114 (
            .O(N__64342),
            .I(N__64338));
    InMux I__16113 (
            .O(N__64341),
            .I(N__64335));
    LocalMux I__16112 (
            .O(N__64338),
            .I(\ADC_VDC.genclk.t0off_3 ));
    LocalMux I__16111 (
            .O(N__64335),
            .I(\ADC_VDC.genclk.t0off_3 ));
    InMux I__16110 (
            .O(N__64330),
            .I(\ADC_VDC.genclk.n20738 ));
    CascadeMux I__16109 (
            .O(N__64327),
            .I(N__64323));
    CascadeMux I__16108 (
            .O(N__64326),
            .I(N__64320));
    InMux I__16107 (
            .O(N__64323),
            .I(N__64317));
    InMux I__16106 (
            .O(N__64320),
            .I(N__64314));
    LocalMux I__16105 (
            .O(N__64317),
            .I(N__64311));
    LocalMux I__16104 (
            .O(N__64314),
            .I(\ADC_VDC.genclk.t0off_4 ));
    Odrv4 I__16103 (
            .O(N__64311),
            .I(\ADC_VDC.genclk.t0off_4 ));
    InMux I__16102 (
            .O(N__64306),
            .I(\ADC_VDC.genclk.n20739 ));
    InMux I__16101 (
            .O(N__64303),
            .I(N__64299));
    InMux I__16100 (
            .O(N__64302),
            .I(N__64296));
    LocalMux I__16099 (
            .O(N__64299),
            .I(\ADC_VDC.genclk.t0off_5 ));
    LocalMux I__16098 (
            .O(N__64296),
            .I(\ADC_VDC.genclk.t0off_5 ));
    InMux I__16097 (
            .O(N__64291),
            .I(\ADC_VDC.genclk.n20740 ));
    CascadeMux I__16096 (
            .O(N__64288),
            .I(N__64285));
    InMux I__16095 (
            .O(N__64285),
            .I(N__64281));
    InMux I__16094 (
            .O(N__64284),
            .I(N__64278));
    LocalMux I__16093 (
            .O(N__64281),
            .I(\ADC_VDC.genclk.t0off_6 ));
    LocalMux I__16092 (
            .O(N__64278),
            .I(\ADC_VDC.genclk.t0off_6 ));
    InMux I__16091 (
            .O(N__64273),
            .I(\ADC_VDC.genclk.n20741 ));
    CascadeMux I__16090 (
            .O(N__64270),
            .I(N__64266));
    InMux I__16089 (
            .O(N__64269),
            .I(N__64263));
    InMux I__16088 (
            .O(N__64266),
            .I(N__64260));
    LocalMux I__16087 (
            .O(N__64263),
            .I(\ADC_VDC.genclk.t0off_7 ));
    LocalMux I__16086 (
            .O(N__64260),
            .I(\ADC_VDC.genclk.t0off_7 ));
    InMux I__16085 (
            .O(N__64255),
            .I(\ADC_VDC.genclk.n20742 ));
    InMux I__16084 (
            .O(N__64252),
            .I(N__64249));
    LocalMux I__16083 (
            .O(N__64249),
            .I(\ADC_VDC.genclk.n26 ));
    CascadeMux I__16082 (
            .O(N__64246),
            .I(\ADC_VDC.genclk.n22305_cascade_ ));
    InMux I__16081 (
            .O(N__64243),
            .I(N__64240));
    LocalMux I__16080 (
            .O(N__64240),
            .I(\ADC_VDC.genclk.n27 ));
    InMux I__16079 (
            .O(N__64237),
            .I(N__64234));
    LocalMux I__16078 (
            .O(N__64234),
            .I(N__64231));
    Odrv4 I__16077 (
            .O(N__64231),
            .I(\ADC_VDC.genclk.n22303 ));
    InMux I__16076 (
            .O(N__64228),
            .I(N__64224));
    InMux I__16075 (
            .O(N__64227),
            .I(N__64221));
    LocalMux I__16074 (
            .O(N__64224),
            .I(N__64211));
    LocalMux I__16073 (
            .O(N__64221),
            .I(N__64211));
    InMux I__16072 (
            .O(N__64220),
            .I(N__64206));
    InMux I__16071 (
            .O(N__64219),
            .I(N__64206));
    InMux I__16070 (
            .O(N__64218),
            .I(N__64203));
    InMux I__16069 (
            .O(N__64217),
            .I(N__64198));
    InMux I__16068 (
            .O(N__64216),
            .I(N__64198));
    Odrv12 I__16067 (
            .O(N__64211),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__16066 (
            .O(N__64206),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__16065 (
            .O(N__64203),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__16064 (
            .O(N__64198),
            .I(\ADC_VDC.genclk.div_state_1 ));
    CascadeMux I__16063 (
            .O(N__64189),
            .I(\ADC_VDC.genclk.n22303_cascade_ ));
    InMux I__16062 (
            .O(N__64186),
            .I(N__64183));
    LocalMux I__16061 (
            .O(N__64183),
            .I(N__64180));
    Span4Mux_v I__16060 (
            .O(N__64180),
            .I(N__64176));
    InMux I__16059 (
            .O(N__64179),
            .I(N__64173));
    Odrv4 I__16058 (
            .O(N__64176),
            .I(\ADC_VDC.genclk.n22302 ));
    LocalMux I__16057 (
            .O(N__64173),
            .I(\ADC_VDC.genclk.n22302 ));
    CascadeMux I__16056 (
            .O(N__64168),
            .I(N__64164));
    InMux I__16055 (
            .O(N__64167),
            .I(N__64154));
    InMux I__16054 (
            .O(N__64164),
            .I(N__64154));
    InMux I__16053 (
            .O(N__64163),
            .I(N__64154));
    InMux I__16052 (
            .O(N__64162),
            .I(N__64151));
    InMux I__16051 (
            .O(N__64161),
            .I(N__64148));
    LocalMux I__16050 (
            .O(N__64154),
            .I(N__64143));
    LocalMux I__16049 (
            .O(N__64151),
            .I(N__64143));
    LocalMux I__16048 (
            .O(N__64148),
            .I(\ADC_VDC.genclk.div_state_0 ));
    Odrv4 I__16047 (
            .O(N__64143),
            .I(\ADC_VDC.genclk.div_state_0 ));
    InMux I__16046 (
            .O(N__64138),
            .I(N__64135));
    LocalMux I__16045 (
            .O(N__64135),
            .I(\ADC_VDC.genclk.n28 ));
    IoInMux I__16044 (
            .O(N__64132),
            .I(N__64129));
    LocalMux I__16043 (
            .O(N__64129),
            .I(N__64126));
    IoSpan4Mux I__16042 (
            .O(N__64126),
            .I(N__64123));
    IoSpan4Mux I__16041 (
            .O(N__64123),
            .I(N__64120));
    IoSpan4Mux I__16040 (
            .O(N__64120),
            .I(N__64117));
    Span4Mux_s3_h I__16039 (
            .O(N__64117),
            .I(N__64114));
    Odrv4 I__16038 (
            .O(N__64114),
            .I(ICE_GPMI_0));
    InMux I__16037 (
            .O(N__64111),
            .I(N__64102));
    InMux I__16036 (
            .O(N__64110),
            .I(N__64102));
    InMux I__16035 (
            .O(N__64109),
            .I(N__64102));
    LocalMux I__16034 (
            .O(N__64102),
            .I(N__64098));
    CascadeMux I__16033 (
            .O(N__64101),
            .I(N__64092));
    Span4Mux_v I__16032 (
            .O(N__64098),
            .I(N__64085));
    InMux I__16031 (
            .O(N__64097),
            .I(N__64080));
    InMux I__16030 (
            .O(N__64096),
            .I(N__64080));
    InMux I__16029 (
            .O(N__64095),
            .I(N__64067));
    InMux I__16028 (
            .O(N__64092),
            .I(N__64067));
    InMux I__16027 (
            .O(N__64091),
            .I(N__64067));
    InMux I__16026 (
            .O(N__64090),
            .I(N__64067));
    InMux I__16025 (
            .O(N__64089),
            .I(N__64062));
    InMux I__16024 (
            .O(N__64088),
            .I(N__64059));
    Span4Mux_h I__16023 (
            .O(N__64085),
            .I(N__64054));
    LocalMux I__16022 (
            .O(N__64080),
            .I(N__64054));
    InMux I__16021 (
            .O(N__64079),
            .I(N__64051));
    InMux I__16020 (
            .O(N__64078),
            .I(N__64041));
    InMux I__16019 (
            .O(N__64077),
            .I(N__64041));
    InMux I__16018 (
            .O(N__64076),
            .I(N__64041));
    LocalMux I__16017 (
            .O(N__64067),
            .I(N__64038));
    CascadeMux I__16016 (
            .O(N__64066),
            .I(N__64035));
    InMux I__16015 (
            .O(N__64065),
            .I(N__64026));
    LocalMux I__16014 (
            .O(N__64062),
            .I(N__64017));
    LocalMux I__16013 (
            .O(N__64059),
            .I(N__64017));
    Span4Mux_v I__16012 (
            .O(N__64054),
            .I(N__64012));
    LocalMux I__16011 (
            .O(N__64051),
            .I(N__64012));
    CascadeMux I__16010 (
            .O(N__64050),
            .I(N__64008));
    InMux I__16009 (
            .O(N__64049),
            .I(N__64001));
    InMux I__16008 (
            .O(N__64048),
            .I(N__64001));
    LocalMux I__16007 (
            .O(N__64041),
            .I(N__63998));
    Span4Mux_v I__16006 (
            .O(N__64038),
            .I(N__63995));
    InMux I__16005 (
            .O(N__64035),
            .I(N__63980));
    InMux I__16004 (
            .O(N__64034),
            .I(N__63980));
    InMux I__16003 (
            .O(N__64033),
            .I(N__63973));
    InMux I__16002 (
            .O(N__64032),
            .I(N__63973));
    InMux I__16001 (
            .O(N__64031),
            .I(N__63973));
    InMux I__16000 (
            .O(N__64030),
            .I(N__63970));
    CascadeMux I__15999 (
            .O(N__64029),
            .I(N__63967));
    LocalMux I__15998 (
            .O(N__64026),
            .I(N__63963));
    InMux I__15997 (
            .O(N__64025),
            .I(N__63960));
    InMux I__15996 (
            .O(N__64024),
            .I(N__63956));
    InMux I__15995 (
            .O(N__64023),
            .I(N__63951));
    InMux I__15994 (
            .O(N__64022),
            .I(N__63951));
    Span4Mux_v I__15993 (
            .O(N__64017),
            .I(N__63946));
    Span4Mux_v I__15992 (
            .O(N__64012),
            .I(N__63946));
    InMux I__15991 (
            .O(N__64011),
            .I(N__63941));
    InMux I__15990 (
            .O(N__64008),
            .I(N__63941));
    InMux I__15989 (
            .O(N__64007),
            .I(N__63936));
    InMux I__15988 (
            .O(N__64006),
            .I(N__63936));
    LocalMux I__15987 (
            .O(N__64001),
            .I(N__63931));
    Span4Mux_h I__15986 (
            .O(N__63998),
            .I(N__63931));
    Span4Mux_h I__15985 (
            .O(N__63995),
            .I(N__63928));
    InMux I__15984 (
            .O(N__63994),
            .I(N__63923));
    InMux I__15983 (
            .O(N__63993),
            .I(N__63923));
    InMux I__15982 (
            .O(N__63992),
            .I(N__63920));
    InMux I__15981 (
            .O(N__63991),
            .I(N__63911));
    InMux I__15980 (
            .O(N__63990),
            .I(N__63911));
    InMux I__15979 (
            .O(N__63989),
            .I(N__63911));
    InMux I__15978 (
            .O(N__63988),
            .I(N__63911));
    CascadeMux I__15977 (
            .O(N__63987),
            .I(N__63905));
    CascadeMux I__15976 (
            .O(N__63986),
            .I(N__63902));
    InMux I__15975 (
            .O(N__63985),
            .I(N__63899));
    LocalMux I__15974 (
            .O(N__63980),
            .I(N__63896));
    LocalMux I__15973 (
            .O(N__63973),
            .I(N__63893));
    LocalMux I__15972 (
            .O(N__63970),
            .I(N__63890));
    InMux I__15971 (
            .O(N__63967),
            .I(N__63885));
    InMux I__15970 (
            .O(N__63966),
            .I(N__63882));
    Span4Mux_h I__15969 (
            .O(N__63963),
            .I(N__63879));
    LocalMux I__15968 (
            .O(N__63960),
            .I(N__63876));
    InMux I__15967 (
            .O(N__63959),
            .I(N__63873));
    LocalMux I__15966 (
            .O(N__63956),
            .I(N__63868));
    LocalMux I__15965 (
            .O(N__63951),
            .I(N__63868));
    Span4Mux_h I__15964 (
            .O(N__63946),
            .I(N__63865));
    LocalMux I__15963 (
            .O(N__63941),
            .I(N__63860));
    LocalMux I__15962 (
            .O(N__63936),
            .I(N__63860));
    Span4Mux_v I__15961 (
            .O(N__63931),
            .I(N__63853));
    Span4Mux_v I__15960 (
            .O(N__63928),
            .I(N__63853));
    LocalMux I__15959 (
            .O(N__63923),
            .I(N__63853));
    LocalMux I__15958 (
            .O(N__63920),
            .I(N__63848));
    LocalMux I__15957 (
            .O(N__63911),
            .I(N__63848));
    InMux I__15956 (
            .O(N__63910),
            .I(N__63845));
    InMux I__15955 (
            .O(N__63909),
            .I(N__63836));
    InMux I__15954 (
            .O(N__63908),
            .I(N__63836));
    InMux I__15953 (
            .O(N__63905),
            .I(N__63836));
    InMux I__15952 (
            .O(N__63902),
            .I(N__63836));
    LocalMux I__15951 (
            .O(N__63899),
            .I(N__63827));
    Span4Mux_v I__15950 (
            .O(N__63896),
            .I(N__63827));
    Span4Mux_v I__15949 (
            .O(N__63893),
            .I(N__63827));
    Span4Mux_v I__15948 (
            .O(N__63890),
            .I(N__63827));
    InMux I__15947 (
            .O(N__63889),
            .I(N__63822));
    InMux I__15946 (
            .O(N__63888),
            .I(N__63822));
    LocalMux I__15945 (
            .O(N__63885),
            .I(N__63815));
    LocalMux I__15944 (
            .O(N__63882),
            .I(N__63815));
    Span4Mux_h I__15943 (
            .O(N__63879),
            .I(N__63815));
    Span4Mux_v I__15942 (
            .O(N__63876),
            .I(N__63802));
    LocalMux I__15941 (
            .O(N__63873),
            .I(N__63802));
    Span4Mux_h I__15940 (
            .O(N__63868),
            .I(N__63802));
    Span4Mux_h I__15939 (
            .O(N__63865),
            .I(N__63802));
    Span4Mux_v I__15938 (
            .O(N__63860),
            .I(N__63802));
    Span4Mux_v I__15937 (
            .O(N__63853),
            .I(N__63802));
    Span12Mux_v I__15936 (
            .O(N__63848),
            .I(N__63799));
    LocalMux I__15935 (
            .O(N__63845),
            .I(comm_state_2));
    LocalMux I__15934 (
            .O(N__63836),
            .I(comm_state_2));
    Odrv4 I__15933 (
            .O(N__63827),
            .I(comm_state_2));
    LocalMux I__15932 (
            .O(N__63822),
            .I(comm_state_2));
    Odrv4 I__15931 (
            .O(N__63815),
            .I(comm_state_2));
    Odrv4 I__15930 (
            .O(N__63802),
            .I(comm_state_2));
    Odrv12 I__15929 (
            .O(N__63799),
            .I(comm_state_2));
    CascadeMux I__15928 (
            .O(N__63784),
            .I(N__63774));
    InMux I__15927 (
            .O(N__63783),
            .I(N__63771));
    CascadeMux I__15926 (
            .O(N__63782),
            .I(N__63757));
    CascadeMux I__15925 (
            .O(N__63781),
            .I(N__63753));
    CascadeMux I__15924 (
            .O(N__63780),
            .I(N__63749));
    CascadeMux I__15923 (
            .O(N__63779),
            .I(N__63745));
    InMux I__15922 (
            .O(N__63778),
            .I(N__63732));
    InMux I__15921 (
            .O(N__63777),
            .I(N__63727));
    InMux I__15920 (
            .O(N__63774),
            .I(N__63727));
    LocalMux I__15919 (
            .O(N__63771),
            .I(N__63719));
    CascadeMux I__15918 (
            .O(N__63770),
            .I(N__63714));
    CascadeMux I__15917 (
            .O(N__63769),
            .I(N__63711));
    CascadeMux I__15916 (
            .O(N__63768),
            .I(N__63708));
    CascadeMux I__15915 (
            .O(N__63767),
            .I(N__63705));
    CascadeMux I__15914 (
            .O(N__63766),
            .I(N__63702));
    CascadeMux I__15913 (
            .O(N__63765),
            .I(N__63699));
    CascadeMux I__15912 (
            .O(N__63764),
            .I(N__63696));
    CascadeMux I__15911 (
            .O(N__63763),
            .I(N__63693));
    CascadeMux I__15910 (
            .O(N__63762),
            .I(N__63690));
    InMux I__15909 (
            .O(N__63761),
            .I(N__63687));
    InMux I__15908 (
            .O(N__63760),
            .I(N__63670));
    InMux I__15907 (
            .O(N__63757),
            .I(N__63670));
    InMux I__15906 (
            .O(N__63756),
            .I(N__63670));
    InMux I__15905 (
            .O(N__63753),
            .I(N__63670));
    InMux I__15904 (
            .O(N__63752),
            .I(N__63670));
    InMux I__15903 (
            .O(N__63749),
            .I(N__63670));
    InMux I__15902 (
            .O(N__63748),
            .I(N__63670));
    InMux I__15901 (
            .O(N__63745),
            .I(N__63670));
    InMux I__15900 (
            .O(N__63744),
            .I(N__63667));
    InMux I__15899 (
            .O(N__63743),
            .I(N__63656));
    InMux I__15898 (
            .O(N__63742),
            .I(N__63656));
    InMux I__15897 (
            .O(N__63741),
            .I(N__63656));
    InMux I__15896 (
            .O(N__63740),
            .I(N__63656));
    InMux I__15895 (
            .O(N__63739),
            .I(N__63656));
    InMux I__15894 (
            .O(N__63738),
            .I(N__63651));
    CascadeMux I__15893 (
            .O(N__63737),
            .I(N__63645));
    InMux I__15892 (
            .O(N__63736),
            .I(N__63637));
    InMux I__15891 (
            .O(N__63735),
            .I(N__63637));
    LocalMux I__15890 (
            .O(N__63732),
            .I(N__63634));
    LocalMux I__15889 (
            .O(N__63727),
            .I(N__63631));
    InMux I__15888 (
            .O(N__63726),
            .I(N__63628));
    InMux I__15887 (
            .O(N__63725),
            .I(N__63625));
    InMux I__15886 (
            .O(N__63724),
            .I(N__63622));
    CascadeMux I__15885 (
            .O(N__63723),
            .I(N__63619));
    InMux I__15884 (
            .O(N__63722),
            .I(N__63614));
    Span4Mux_v I__15883 (
            .O(N__63719),
            .I(N__63598));
    InMux I__15882 (
            .O(N__63718),
            .I(N__63589));
    InMux I__15881 (
            .O(N__63717),
            .I(N__63589));
    InMux I__15880 (
            .O(N__63714),
            .I(N__63580));
    InMux I__15879 (
            .O(N__63711),
            .I(N__63580));
    InMux I__15878 (
            .O(N__63708),
            .I(N__63580));
    InMux I__15877 (
            .O(N__63705),
            .I(N__63580));
    InMux I__15876 (
            .O(N__63702),
            .I(N__63571));
    InMux I__15875 (
            .O(N__63699),
            .I(N__63571));
    InMux I__15874 (
            .O(N__63696),
            .I(N__63571));
    InMux I__15873 (
            .O(N__63693),
            .I(N__63571));
    InMux I__15872 (
            .O(N__63690),
            .I(N__63568));
    LocalMux I__15871 (
            .O(N__63687),
            .I(N__63559));
    LocalMux I__15870 (
            .O(N__63670),
            .I(N__63559));
    LocalMux I__15869 (
            .O(N__63667),
            .I(N__63559));
    LocalMux I__15868 (
            .O(N__63656),
            .I(N__63559));
    InMux I__15867 (
            .O(N__63655),
            .I(N__63554));
    InMux I__15866 (
            .O(N__63654),
            .I(N__63554));
    LocalMux I__15865 (
            .O(N__63651),
            .I(N__63551));
    InMux I__15864 (
            .O(N__63650),
            .I(N__63548));
    InMux I__15863 (
            .O(N__63649),
            .I(N__63545));
    InMux I__15862 (
            .O(N__63648),
            .I(N__63542));
    InMux I__15861 (
            .O(N__63645),
            .I(N__63536));
    InMux I__15860 (
            .O(N__63644),
            .I(N__63529));
    InMux I__15859 (
            .O(N__63643),
            .I(N__63529));
    InMux I__15858 (
            .O(N__63642),
            .I(N__63529));
    LocalMux I__15857 (
            .O(N__63637),
            .I(N__63514));
    Span4Mux_h I__15856 (
            .O(N__63634),
            .I(N__63514));
    Span4Mux_v I__15855 (
            .O(N__63631),
            .I(N__63514));
    LocalMux I__15854 (
            .O(N__63628),
            .I(N__63514));
    LocalMux I__15853 (
            .O(N__63625),
            .I(N__63514));
    LocalMux I__15852 (
            .O(N__63622),
            .I(N__63511));
    InMux I__15851 (
            .O(N__63619),
            .I(N__63506));
    InMux I__15850 (
            .O(N__63618),
            .I(N__63506));
    SRMux I__15849 (
            .O(N__63617),
            .I(N__63501));
    LocalMux I__15848 (
            .O(N__63614),
            .I(N__63498));
    InMux I__15847 (
            .O(N__63613),
            .I(N__63495));
    InMux I__15846 (
            .O(N__63612),
            .I(N__63479));
    InMux I__15845 (
            .O(N__63611),
            .I(N__63474));
    InMux I__15844 (
            .O(N__63610),
            .I(N__63474));
    InMux I__15843 (
            .O(N__63609),
            .I(N__63469));
    InMux I__15842 (
            .O(N__63608),
            .I(N__63469));
    InMux I__15841 (
            .O(N__63607),
            .I(N__63466));
    InMux I__15840 (
            .O(N__63606),
            .I(N__63457));
    InMux I__15839 (
            .O(N__63605),
            .I(N__63457));
    InMux I__15838 (
            .O(N__63604),
            .I(N__63457));
    InMux I__15837 (
            .O(N__63603),
            .I(N__63457));
    InMux I__15836 (
            .O(N__63602),
            .I(N__63454));
    InMux I__15835 (
            .O(N__63601),
            .I(N__63451));
    Span4Mux_h I__15834 (
            .O(N__63598),
            .I(N__63448));
    InMux I__15833 (
            .O(N__63597),
            .I(N__63445));
    InMux I__15832 (
            .O(N__63596),
            .I(N__63438));
    InMux I__15831 (
            .O(N__63595),
            .I(N__63438));
    InMux I__15830 (
            .O(N__63594),
            .I(N__63438));
    LocalMux I__15829 (
            .O(N__63589),
            .I(N__63421));
    LocalMux I__15828 (
            .O(N__63580),
            .I(N__63421));
    LocalMux I__15827 (
            .O(N__63571),
            .I(N__63421));
    LocalMux I__15826 (
            .O(N__63568),
            .I(N__63421));
    Span4Mux_v I__15825 (
            .O(N__63559),
            .I(N__63421));
    LocalMux I__15824 (
            .O(N__63554),
            .I(N__63421));
    Span4Mux_v I__15823 (
            .O(N__63551),
            .I(N__63421));
    LocalMux I__15822 (
            .O(N__63548),
            .I(N__63421));
    LocalMux I__15821 (
            .O(N__63545),
            .I(N__63418));
    LocalMux I__15820 (
            .O(N__63542),
            .I(N__63415));
    InMux I__15819 (
            .O(N__63541),
            .I(N__63412));
    InMux I__15818 (
            .O(N__63540),
            .I(N__63407));
    InMux I__15817 (
            .O(N__63539),
            .I(N__63407));
    LocalMux I__15816 (
            .O(N__63536),
            .I(N__63402));
    LocalMux I__15815 (
            .O(N__63529),
            .I(N__63402));
    InMux I__15814 (
            .O(N__63528),
            .I(N__63397));
    InMux I__15813 (
            .O(N__63527),
            .I(N__63397));
    InMux I__15812 (
            .O(N__63526),
            .I(N__63394));
    InMux I__15811 (
            .O(N__63525),
            .I(N__63390));
    Span4Mux_v I__15810 (
            .O(N__63514),
            .I(N__63383));
    Span4Mux_v I__15809 (
            .O(N__63511),
            .I(N__63383));
    LocalMux I__15808 (
            .O(N__63506),
            .I(N__63383));
    InMux I__15807 (
            .O(N__63505),
            .I(N__63373));
    InMux I__15806 (
            .O(N__63504),
            .I(N__63373));
    LocalMux I__15805 (
            .O(N__63501),
            .I(N__63366));
    Span4Mux_h I__15804 (
            .O(N__63498),
            .I(N__63366));
    LocalMux I__15803 (
            .O(N__63495),
            .I(N__63366));
    InMux I__15802 (
            .O(N__63494),
            .I(N__63359));
    InMux I__15801 (
            .O(N__63493),
            .I(N__63359));
    InMux I__15800 (
            .O(N__63492),
            .I(N__63359));
    InMux I__15799 (
            .O(N__63491),
            .I(N__63354));
    InMux I__15798 (
            .O(N__63490),
            .I(N__63349));
    InMux I__15797 (
            .O(N__63489),
            .I(N__63349));
    InMux I__15796 (
            .O(N__63488),
            .I(N__63346));
    InMux I__15795 (
            .O(N__63487),
            .I(N__63341));
    InMux I__15794 (
            .O(N__63486),
            .I(N__63341));
    InMux I__15793 (
            .O(N__63485),
            .I(N__63338));
    InMux I__15792 (
            .O(N__63484),
            .I(N__63331));
    InMux I__15791 (
            .O(N__63483),
            .I(N__63331));
    InMux I__15790 (
            .O(N__63482),
            .I(N__63331));
    LocalMux I__15789 (
            .O(N__63479),
            .I(N__63320));
    LocalMux I__15788 (
            .O(N__63474),
            .I(N__63320));
    LocalMux I__15787 (
            .O(N__63469),
            .I(N__63320));
    LocalMux I__15786 (
            .O(N__63466),
            .I(N__63320));
    LocalMux I__15785 (
            .O(N__63457),
            .I(N__63320));
    LocalMux I__15784 (
            .O(N__63454),
            .I(N__63317));
    LocalMux I__15783 (
            .O(N__63451),
            .I(N__63314));
    Span4Mux_h I__15782 (
            .O(N__63448),
            .I(N__63305));
    LocalMux I__15781 (
            .O(N__63445),
            .I(N__63305));
    LocalMux I__15780 (
            .O(N__63438),
            .I(N__63305));
    Span4Mux_v I__15779 (
            .O(N__63421),
            .I(N__63305));
    Span4Mux_v I__15778 (
            .O(N__63418),
            .I(N__63300));
    Span4Mux_v I__15777 (
            .O(N__63415),
            .I(N__63300));
    LocalMux I__15776 (
            .O(N__63412),
            .I(N__63291));
    LocalMux I__15775 (
            .O(N__63407),
            .I(N__63291));
    Span4Mux_v I__15774 (
            .O(N__63402),
            .I(N__63291));
    LocalMux I__15773 (
            .O(N__63397),
            .I(N__63291));
    LocalMux I__15772 (
            .O(N__63394),
            .I(N__63288));
    InMux I__15771 (
            .O(N__63393),
            .I(N__63285));
    LocalMux I__15770 (
            .O(N__63390),
            .I(N__63282));
    Span4Mux_h I__15769 (
            .O(N__63383),
            .I(N__63279));
    InMux I__15768 (
            .O(N__63382),
            .I(N__63270));
    InMux I__15767 (
            .O(N__63381),
            .I(N__63270));
    InMux I__15766 (
            .O(N__63380),
            .I(N__63270));
    InMux I__15765 (
            .O(N__63379),
            .I(N__63270));
    InMux I__15764 (
            .O(N__63378),
            .I(N__63267));
    LocalMux I__15763 (
            .O(N__63373),
            .I(N__63260));
    Span4Mux_h I__15762 (
            .O(N__63366),
            .I(N__63260));
    LocalMux I__15761 (
            .O(N__63359),
            .I(N__63260));
    InMux I__15760 (
            .O(N__63358),
            .I(N__63255));
    InMux I__15759 (
            .O(N__63357),
            .I(N__63255));
    LocalMux I__15758 (
            .O(N__63354),
            .I(N__63240));
    LocalMux I__15757 (
            .O(N__63349),
            .I(N__63240));
    LocalMux I__15756 (
            .O(N__63346),
            .I(N__63240));
    LocalMux I__15755 (
            .O(N__63341),
            .I(N__63240));
    LocalMux I__15754 (
            .O(N__63338),
            .I(N__63240));
    LocalMux I__15753 (
            .O(N__63331),
            .I(N__63240));
    Span12Mux_v I__15752 (
            .O(N__63320),
            .I(N__63240));
    Span4Mux_v I__15751 (
            .O(N__63317),
            .I(N__63229));
    Span4Mux_v I__15750 (
            .O(N__63314),
            .I(N__63229));
    Span4Mux_v I__15749 (
            .O(N__63305),
            .I(N__63229));
    Span4Mux_h I__15748 (
            .O(N__63300),
            .I(N__63229));
    Span4Mux_v I__15747 (
            .O(N__63291),
            .I(N__63229));
    Span12Mux_h I__15746 (
            .O(N__63288),
            .I(N__63218));
    LocalMux I__15745 (
            .O(N__63285),
            .I(N__63218));
    Span12Mux_s9_v I__15744 (
            .O(N__63282),
            .I(N__63218));
    Sp12to4 I__15743 (
            .O(N__63279),
            .I(N__63218));
    LocalMux I__15742 (
            .O(N__63270),
            .I(N__63218));
    LocalMux I__15741 (
            .O(N__63267),
            .I(comm_state_3));
    Odrv4 I__15740 (
            .O(N__63260),
            .I(comm_state_3));
    LocalMux I__15739 (
            .O(N__63255),
            .I(comm_state_3));
    Odrv12 I__15738 (
            .O(N__63240),
            .I(comm_state_3));
    Odrv4 I__15737 (
            .O(N__63229),
            .I(comm_state_3));
    Odrv12 I__15736 (
            .O(N__63218),
            .I(comm_state_3));
    CascadeMux I__15735 (
            .O(N__63205),
            .I(N__63201));
    InMux I__15734 (
            .O(N__63204),
            .I(N__63197));
    InMux I__15733 (
            .O(N__63201),
            .I(N__63191));
    CascadeMux I__15732 (
            .O(N__63200),
            .I(N__63185));
    LocalMux I__15731 (
            .O(N__63197),
            .I(N__63182));
    InMux I__15730 (
            .O(N__63196),
            .I(N__63177));
    InMux I__15729 (
            .O(N__63195),
            .I(N__63177));
    InMux I__15728 (
            .O(N__63194),
            .I(N__63174));
    LocalMux I__15727 (
            .O(N__63191),
            .I(N__63170));
    InMux I__15726 (
            .O(N__63190),
            .I(N__63167));
    CascadeMux I__15725 (
            .O(N__63189),
            .I(N__63164));
    InMux I__15724 (
            .O(N__63188),
            .I(N__63157));
    InMux I__15723 (
            .O(N__63185),
            .I(N__63157));
    Span4Mux_v I__15722 (
            .O(N__63182),
            .I(N__63152));
    LocalMux I__15721 (
            .O(N__63177),
            .I(N__63152));
    LocalMux I__15720 (
            .O(N__63174),
            .I(N__63149));
    InMux I__15719 (
            .O(N__63173),
            .I(N__63146));
    Span4Mux_v I__15718 (
            .O(N__63170),
            .I(N__63140));
    LocalMux I__15717 (
            .O(N__63167),
            .I(N__63140));
    InMux I__15716 (
            .O(N__63164),
            .I(N__63133));
    InMux I__15715 (
            .O(N__63163),
            .I(N__63133));
    InMux I__15714 (
            .O(N__63162),
            .I(N__63133));
    LocalMux I__15713 (
            .O(N__63157),
            .I(N__63128));
    Span4Mux_v I__15712 (
            .O(N__63152),
            .I(N__63128));
    Span4Mux_h I__15711 (
            .O(N__63149),
            .I(N__63125));
    LocalMux I__15710 (
            .O(N__63146),
            .I(N__63122));
    InMux I__15709 (
            .O(N__63145),
            .I(N__63119));
    Span4Mux_h I__15708 (
            .O(N__63140),
            .I(N__63114));
    LocalMux I__15707 (
            .O(N__63133),
            .I(N__63114));
    Span4Mux_v I__15706 (
            .O(N__63128),
            .I(N__63111));
    Span4Mux_v I__15705 (
            .O(N__63125),
            .I(N__63105));
    Span4Mux_v I__15704 (
            .O(N__63122),
            .I(N__63105));
    LocalMux I__15703 (
            .O(N__63119),
            .I(N__63100));
    Span4Mux_h I__15702 (
            .O(N__63114),
            .I(N__63100));
    Sp12to4 I__15701 (
            .O(N__63111),
            .I(N__63097));
    InMux I__15700 (
            .O(N__63110),
            .I(N__63094));
    Odrv4 I__15699 (
            .O(N__63105),
            .I(n12966));
    Odrv4 I__15698 (
            .O(N__63100),
            .I(n12966));
    Odrv12 I__15697 (
            .O(N__63097),
            .I(n12966));
    LocalMux I__15696 (
            .O(N__63094),
            .I(n12966));
    CascadeMux I__15695 (
            .O(N__63085),
            .I(N__63067));
    InMux I__15694 (
            .O(N__63084),
            .I(N__63061));
    InMux I__15693 (
            .O(N__63083),
            .I(N__63061));
    InMux I__15692 (
            .O(N__63082),
            .I(N__63052));
    InMux I__15691 (
            .O(N__63081),
            .I(N__63042));
    InMux I__15690 (
            .O(N__63080),
            .I(N__63039));
    InMux I__15689 (
            .O(N__63079),
            .I(N__63034));
    InMux I__15688 (
            .O(N__63078),
            .I(N__63034));
    InMux I__15687 (
            .O(N__63077),
            .I(N__63031));
    InMux I__15686 (
            .O(N__63076),
            .I(N__63024));
    CascadeMux I__15685 (
            .O(N__63075),
            .I(N__63021));
    InMux I__15684 (
            .O(N__63074),
            .I(N__63018));
    InMux I__15683 (
            .O(N__63073),
            .I(N__63015));
    InMux I__15682 (
            .O(N__63072),
            .I(N__63012));
    InMux I__15681 (
            .O(N__63071),
            .I(N__63003));
    InMux I__15680 (
            .O(N__63070),
            .I(N__63003));
    InMux I__15679 (
            .O(N__63067),
            .I(N__63003));
    InMux I__15678 (
            .O(N__63066),
            .I(N__63003));
    LocalMux I__15677 (
            .O(N__63061),
            .I(N__63000));
    InMux I__15676 (
            .O(N__63060),
            .I(N__62991));
    InMux I__15675 (
            .O(N__63059),
            .I(N__62991));
    InMux I__15674 (
            .O(N__63058),
            .I(N__62991));
    InMux I__15673 (
            .O(N__63057),
            .I(N__62991));
    InMux I__15672 (
            .O(N__63056),
            .I(N__62986));
    InMux I__15671 (
            .O(N__63055),
            .I(N__62986));
    LocalMux I__15670 (
            .O(N__63052),
            .I(N__62983));
    InMux I__15669 (
            .O(N__63051),
            .I(N__62980));
    InMux I__15668 (
            .O(N__63050),
            .I(N__62973));
    InMux I__15667 (
            .O(N__63049),
            .I(N__62973));
    InMux I__15666 (
            .O(N__63048),
            .I(N__62973));
    InMux I__15665 (
            .O(N__63047),
            .I(N__62970));
    InMux I__15664 (
            .O(N__63046),
            .I(N__62964));
    InMux I__15663 (
            .O(N__63045),
            .I(N__62964));
    LocalMux I__15662 (
            .O(N__63042),
            .I(N__62957));
    LocalMux I__15661 (
            .O(N__63039),
            .I(N__62957));
    LocalMux I__15660 (
            .O(N__63034),
            .I(N__62957));
    LocalMux I__15659 (
            .O(N__63031),
            .I(N__62954));
    InMux I__15658 (
            .O(N__63030),
            .I(N__62949));
    InMux I__15657 (
            .O(N__63029),
            .I(N__62949));
    InMux I__15656 (
            .O(N__63028),
            .I(N__62944));
    InMux I__15655 (
            .O(N__63027),
            .I(N__62944));
    LocalMux I__15654 (
            .O(N__63024),
            .I(N__62940));
    InMux I__15653 (
            .O(N__63021),
            .I(N__62937));
    LocalMux I__15652 (
            .O(N__63018),
            .I(N__62927));
    LocalMux I__15651 (
            .O(N__63015),
            .I(N__62924));
    LocalMux I__15650 (
            .O(N__63012),
            .I(N__62913));
    LocalMux I__15649 (
            .O(N__63003),
            .I(N__62913));
    Span4Mux_v I__15648 (
            .O(N__63000),
            .I(N__62913));
    LocalMux I__15647 (
            .O(N__62991),
            .I(N__62913));
    LocalMux I__15646 (
            .O(N__62986),
            .I(N__62913));
    Span4Mux_v I__15645 (
            .O(N__62983),
            .I(N__62908));
    LocalMux I__15644 (
            .O(N__62980),
            .I(N__62908));
    LocalMux I__15643 (
            .O(N__62973),
            .I(N__62902));
    LocalMux I__15642 (
            .O(N__62970),
            .I(N__62899));
    InMux I__15641 (
            .O(N__62969),
            .I(N__62896));
    LocalMux I__15640 (
            .O(N__62964),
            .I(N__62891));
    Span4Mux_v I__15639 (
            .O(N__62957),
            .I(N__62891));
    Span4Mux_h I__15638 (
            .O(N__62954),
            .I(N__62884));
    LocalMux I__15637 (
            .O(N__62949),
            .I(N__62884));
    LocalMux I__15636 (
            .O(N__62944),
            .I(N__62884));
    InMux I__15635 (
            .O(N__62943),
            .I(N__62881));
    Span4Mux_h I__15634 (
            .O(N__62940),
            .I(N__62878));
    LocalMux I__15633 (
            .O(N__62937),
            .I(N__62875));
    InMux I__15632 (
            .O(N__62936),
            .I(N__62872));
    InMux I__15631 (
            .O(N__62935),
            .I(N__62863));
    InMux I__15630 (
            .O(N__62934),
            .I(N__62863));
    InMux I__15629 (
            .O(N__62933),
            .I(N__62863));
    InMux I__15628 (
            .O(N__62932),
            .I(N__62863));
    InMux I__15627 (
            .O(N__62931),
            .I(N__62858));
    InMux I__15626 (
            .O(N__62930),
            .I(N__62858));
    Span4Mux_h I__15625 (
            .O(N__62927),
            .I(N__62849));
    Span4Mux_v I__15624 (
            .O(N__62924),
            .I(N__62849));
    Span4Mux_v I__15623 (
            .O(N__62913),
            .I(N__62849));
    Span4Mux_v I__15622 (
            .O(N__62908),
            .I(N__62849));
    InMux I__15621 (
            .O(N__62907),
            .I(N__62844));
    InMux I__15620 (
            .O(N__62906),
            .I(N__62844));
    InMux I__15619 (
            .O(N__62905),
            .I(N__62841));
    Sp12to4 I__15618 (
            .O(N__62902),
            .I(N__62836));
    Span12Mux_h I__15617 (
            .O(N__62899),
            .I(N__62836));
    LocalMux I__15616 (
            .O(N__62896),
            .I(N__62831));
    Span4Mux_h I__15615 (
            .O(N__62891),
            .I(N__62831));
    Span4Mux_h I__15614 (
            .O(N__62884),
            .I(N__62822));
    LocalMux I__15613 (
            .O(N__62881),
            .I(N__62822));
    Span4Mux_h I__15612 (
            .O(N__62878),
            .I(N__62822));
    Span4Mux_h I__15611 (
            .O(N__62875),
            .I(N__62822));
    LocalMux I__15610 (
            .O(N__62872),
            .I(comm_state_0));
    LocalMux I__15609 (
            .O(N__62863),
            .I(comm_state_0));
    LocalMux I__15608 (
            .O(N__62858),
            .I(comm_state_0));
    Odrv4 I__15607 (
            .O(N__62849),
            .I(comm_state_0));
    LocalMux I__15606 (
            .O(N__62844),
            .I(comm_state_0));
    LocalMux I__15605 (
            .O(N__62841),
            .I(comm_state_0));
    Odrv12 I__15604 (
            .O(N__62836),
            .I(comm_state_0));
    Odrv4 I__15603 (
            .O(N__62831),
            .I(comm_state_0));
    Odrv4 I__15602 (
            .O(N__62822),
            .I(comm_state_0));
    CEMux I__15601 (
            .O(N__62803),
            .I(N__62800));
    LocalMux I__15600 (
            .O(N__62800),
            .I(N__62797));
    Odrv4 I__15599 (
            .O(N__62797),
            .I(n12045));
    CascadeMux I__15598 (
            .O(N__62794),
            .I(N__62791));
    InMux I__15597 (
            .O(N__62791),
            .I(N__62785));
    InMux I__15596 (
            .O(N__62790),
            .I(N__62781));
    InMux I__15595 (
            .O(N__62789),
            .I(N__62776));
    InMux I__15594 (
            .O(N__62788),
            .I(N__62772));
    LocalMux I__15593 (
            .O(N__62785),
            .I(N__62769));
    InMux I__15592 (
            .O(N__62784),
            .I(N__62766));
    LocalMux I__15591 (
            .O(N__62781),
            .I(N__62763));
    InMux I__15590 (
            .O(N__62780),
            .I(N__62760));
    CascadeMux I__15589 (
            .O(N__62779),
            .I(N__62757));
    LocalMux I__15588 (
            .O(N__62776),
            .I(N__62754));
    CascadeMux I__15587 (
            .O(N__62775),
            .I(N__62751));
    LocalMux I__15586 (
            .O(N__62772),
            .I(N__62748));
    Span4Mux_v I__15585 (
            .O(N__62769),
            .I(N__62743));
    LocalMux I__15584 (
            .O(N__62766),
            .I(N__62743));
    Span4Mux_v I__15583 (
            .O(N__62763),
            .I(N__62740));
    LocalMux I__15582 (
            .O(N__62760),
            .I(N__62737));
    InMux I__15581 (
            .O(N__62757),
            .I(N__62734));
    Span4Mux_h I__15580 (
            .O(N__62754),
            .I(N__62731));
    InMux I__15579 (
            .O(N__62751),
            .I(N__62728));
    Span4Mux_h I__15578 (
            .O(N__62748),
            .I(N__62724));
    Span4Mux_v I__15577 (
            .O(N__62743),
            .I(N__62721));
    Span4Mux_h I__15576 (
            .O(N__62740),
            .I(N__62716));
    Span4Mux_v I__15575 (
            .O(N__62737),
            .I(N__62716));
    LocalMux I__15574 (
            .O(N__62734),
            .I(N__62713));
    Span4Mux_h I__15573 (
            .O(N__62731),
            .I(N__62708));
    LocalMux I__15572 (
            .O(N__62728),
            .I(N__62708));
    InMux I__15571 (
            .O(N__62727),
            .I(N__62705));
    Odrv4 I__15570 (
            .O(N__62724),
            .I(comm_rx_buf_3));
    Odrv4 I__15569 (
            .O(N__62721),
            .I(comm_rx_buf_3));
    Odrv4 I__15568 (
            .O(N__62716),
            .I(comm_rx_buf_3));
    Odrv12 I__15567 (
            .O(N__62713),
            .I(comm_rx_buf_3));
    Odrv4 I__15566 (
            .O(N__62708),
            .I(comm_rx_buf_3));
    LocalMux I__15565 (
            .O(N__62705),
            .I(comm_rx_buf_3));
    InMux I__15564 (
            .O(N__62692),
            .I(N__62686));
    CascadeMux I__15563 (
            .O(N__62691),
            .I(N__62682));
    CascadeMux I__15562 (
            .O(N__62690),
            .I(N__62679));
    InMux I__15561 (
            .O(N__62689),
            .I(N__62667));
    LocalMux I__15560 (
            .O(N__62686),
            .I(N__62664));
    CascadeMux I__15559 (
            .O(N__62685),
            .I(N__62649));
    InMux I__15558 (
            .O(N__62682),
            .I(N__62638));
    InMux I__15557 (
            .O(N__62679),
            .I(N__62638));
    InMux I__15556 (
            .O(N__62678),
            .I(N__62638));
    CascadeMux I__15555 (
            .O(N__62677),
            .I(N__62634));
    CascadeMux I__15554 (
            .O(N__62676),
            .I(N__62612));
    InMux I__15553 (
            .O(N__62675),
            .I(N__62588));
    InMux I__15552 (
            .O(N__62674),
            .I(N__62588));
    InMux I__15551 (
            .O(N__62673),
            .I(N__62588));
    InMux I__15550 (
            .O(N__62672),
            .I(N__62585));
    InMux I__15549 (
            .O(N__62671),
            .I(N__62582));
    InMux I__15548 (
            .O(N__62670),
            .I(N__62579));
    LocalMux I__15547 (
            .O(N__62667),
            .I(N__62576));
    Span4Mux_v I__15546 (
            .O(N__62664),
            .I(N__62573));
    InMux I__15545 (
            .O(N__62663),
            .I(N__62561));
    InMux I__15544 (
            .O(N__62662),
            .I(N__62548));
    InMux I__15543 (
            .O(N__62661),
            .I(N__62548));
    InMux I__15542 (
            .O(N__62660),
            .I(N__62548));
    InMux I__15541 (
            .O(N__62659),
            .I(N__62548));
    InMux I__15540 (
            .O(N__62658),
            .I(N__62548));
    InMux I__15539 (
            .O(N__62657),
            .I(N__62548));
    InMux I__15538 (
            .O(N__62656),
            .I(N__62531));
    InMux I__15537 (
            .O(N__62655),
            .I(N__62531));
    InMux I__15536 (
            .O(N__62654),
            .I(N__62531));
    InMux I__15535 (
            .O(N__62653),
            .I(N__62531));
    InMux I__15534 (
            .O(N__62652),
            .I(N__62531));
    InMux I__15533 (
            .O(N__62649),
            .I(N__62531));
    InMux I__15532 (
            .O(N__62648),
            .I(N__62531));
    InMux I__15531 (
            .O(N__62647),
            .I(N__62531));
    InMux I__15530 (
            .O(N__62646),
            .I(N__62516));
    InMux I__15529 (
            .O(N__62645),
            .I(N__62516));
    LocalMux I__15528 (
            .O(N__62638),
            .I(N__62513));
    InMux I__15527 (
            .O(N__62637),
            .I(N__62510));
    InMux I__15526 (
            .O(N__62634),
            .I(N__62507));
    CascadeMux I__15525 (
            .O(N__62633),
            .I(N__62504));
    InMux I__15524 (
            .O(N__62632),
            .I(N__62487));
    InMux I__15523 (
            .O(N__62631),
            .I(N__62487));
    InMux I__15522 (
            .O(N__62630),
            .I(N__62487));
    InMux I__15521 (
            .O(N__62629),
            .I(N__62487));
    InMux I__15520 (
            .O(N__62628),
            .I(N__62487));
    InMux I__15519 (
            .O(N__62627),
            .I(N__62487));
    InMux I__15518 (
            .O(N__62626),
            .I(N__62487));
    InMux I__15517 (
            .O(N__62625),
            .I(N__62487));
    InMux I__15516 (
            .O(N__62624),
            .I(N__62482));
    InMux I__15515 (
            .O(N__62623),
            .I(N__62463));
    InMux I__15514 (
            .O(N__62622),
            .I(N__62463));
    InMux I__15513 (
            .O(N__62621),
            .I(N__62463));
    InMux I__15512 (
            .O(N__62620),
            .I(N__62463));
    InMux I__15511 (
            .O(N__62619),
            .I(N__62463));
    InMux I__15510 (
            .O(N__62618),
            .I(N__62463));
    InMux I__15509 (
            .O(N__62617),
            .I(N__62463));
    InMux I__15508 (
            .O(N__62616),
            .I(N__62463));
    InMux I__15507 (
            .O(N__62615),
            .I(N__62460));
    InMux I__15506 (
            .O(N__62612),
            .I(N__62451));
    InMux I__15505 (
            .O(N__62611),
            .I(N__62451));
    InMux I__15504 (
            .O(N__62610),
            .I(N__62451));
    InMux I__15503 (
            .O(N__62609),
            .I(N__62451));
    CascadeMux I__15502 (
            .O(N__62608),
            .I(N__62446));
    InMux I__15501 (
            .O(N__62607),
            .I(N__62443));
    InMux I__15500 (
            .O(N__62606),
            .I(N__62440));
    InMux I__15499 (
            .O(N__62605),
            .I(N__62435));
    InMux I__15498 (
            .O(N__62604),
            .I(N__62435));
    InMux I__15497 (
            .O(N__62603),
            .I(N__62432));
    InMux I__15496 (
            .O(N__62602),
            .I(N__62429));
    CascadeMux I__15495 (
            .O(N__62601),
            .I(N__62423));
    InMux I__15494 (
            .O(N__62600),
            .I(N__62418));
    InMux I__15493 (
            .O(N__62599),
            .I(N__62411));
    InMux I__15492 (
            .O(N__62598),
            .I(N__62411));
    InMux I__15491 (
            .O(N__62597),
            .I(N__62411));
    InMux I__15490 (
            .O(N__62596),
            .I(N__62406));
    InMux I__15489 (
            .O(N__62595),
            .I(N__62406));
    LocalMux I__15488 (
            .O(N__62588),
            .I(N__62403));
    LocalMux I__15487 (
            .O(N__62585),
            .I(N__62392));
    LocalMux I__15486 (
            .O(N__62582),
            .I(N__62392));
    LocalMux I__15485 (
            .O(N__62579),
            .I(N__62392));
    Span4Mux_h I__15484 (
            .O(N__62576),
            .I(N__62392));
    Span4Mux_h I__15483 (
            .O(N__62573),
            .I(N__62392));
    InMux I__15482 (
            .O(N__62572),
            .I(N__62385));
    InMux I__15481 (
            .O(N__62571),
            .I(N__62385));
    InMux I__15480 (
            .O(N__62570),
            .I(N__62385));
    InMux I__15479 (
            .O(N__62569),
            .I(N__62380));
    InMux I__15478 (
            .O(N__62568),
            .I(N__62380));
    InMux I__15477 (
            .O(N__62567),
            .I(N__62373));
    InMux I__15476 (
            .O(N__62566),
            .I(N__62373));
    InMux I__15475 (
            .O(N__62565),
            .I(N__62373));
    InMux I__15474 (
            .O(N__62564),
            .I(N__62370));
    LocalMux I__15473 (
            .O(N__62561),
            .I(N__62361));
    LocalMux I__15472 (
            .O(N__62548),
            .I(N__62361));
    LocalMux I__15471 (
            .O(N__62531),
            .I(N__62361));
    InMux I__15470 (
            .O(N__62530),
            .I(N__62358));
    InMux I__15469 (
            .O(N__62529),
            .I(N__62355));
    InMux I__15468 (
            .O(N__62528),
            .I(N__62338));
    InMux I__15467 (
            .O(N__62527),
            .I(N__62338));
    InMux I__15466 (
            .O(N__62526),
            .I(N__62338));
    InMux I__15465 (
            .O(N__62525),
            .I(N__62338));
    InMux I__15464 (
            .O(N__62524),
            .I(N__62338));
    InMux I__15463 (
            .O(N__62523),
            .I(N__62338));
    InMux I__15462 (
            .O(N__62522),
            .I(N__62338));
    InMux I__15461 (
            .O(N__62521),
            .I(N__62338));
    LocalMux I__15460 (
            .O(N__62516),
            .I(N__62335));
    Span4Mux_v I__15459 (
            .O(N__62513),
            .I(N__62332));
    LocalMux I__15458 (
            .O(N__62510),
            .I(N__62327));
    LocalMux I__15457 (
            .O(N__62507),
            .I(N__62327));
    InMux I__15456 (
            .O(N__62504),
            .I(N__62324));
    LocalMux I__15455 (
            .O(N__62487),
            .I(N__62321));
    InMux I__15454 (
            .O(N__62486),
            .I(N__62316));
    InMux I__15453 (
            .O(N__62485),
            .I(N__62316));
    LocalMux I__15452 (
            .O(N__62482),
            .I(N__62313));
    InMux I__15451 (
            .O(N__62481),
            .I(N__62308));
    InMux I__15450 (
            .O(N__62480),
            .I(N__62308));
    LocalMux I__15449 (
            .O(N__62463),
            .I(N__62301));
    LocalMux I__15448 (
            .O(N__62460),
            .I(N__62301));
    LocalMux I__15447 (
            .O(N__62451),
            .I(N__62301));
    InMux I__15446 (
            .O(N__62450),
            .I(N__62298));
    InMux I__15445 (
            .O(N__62449),
            .I(N__62285));
    InMux I__15444 (
            .O(N__62446),
            .I(N__62285));
    LocalMux I__15443 (
            .O(N__62443),
            .I(N__62276));
    LocalMux I__15442 (
            .O(N__62440),
            .I(N__62276));
    LocalMux I__15441 (
            .O(N__62435),
            .I(N__62276));
    LocalMux I__15440 (
            .O(N__62432),
            .I(N__62276));
    LocalMux I__15439 (
            .O(N__62429),
            .I(N__62273));
    InMux I__15438 (
            .O(N__62428),
            .I(N__62260));
    InMux I__15437 (
            .O(N__62427),
            .I(N__62260));
    InMux I__15436 (
            .O(N__62426),
            .I(N__62260));
    InMux I__15435 (
            .O(N__62423),
            .I(N__62260));
    InMux I__15434 (
            .O(N__62422),
            .I(N__62260));
    InMux I__15433 (
            .O(N__62421),
            .I(N__62260));
    LocalMux I__15432 (
            .O(N__62418),
            .I(N__62243));
    LocalMux I__15431 (
            .O(N__62411),
            .I(N__62243));
    LocalMux I__15430 (
            .O(N__62406),
            .I(N__62243));
    Span4Mux_h I__15429 (
            .O(N__62403),
            .I(N__62243));
    Span4Mux_v I__15428 (
            .O(N__62392),
            .I(N__62243));
    LocalMux I__15427 (
            .O(N__62385),
            .I(N__62243));
    LocalMux I__15426 (
            .O(N__62380),
            .I(N__62243));
    LocalMux I__15425 (
            .O(N__62373),
            .I(N__62243));
    LocalMux I__15424 (
            .O(N__62370),
            .I(N__62237));
    InMux I__15423 (
            .O(N__62369),
            .I(N__62232));
    InMux I__15422 (
            .O(N__62368),
            .I(N__62232));
    Span4Mux_h I__15421 (
            .O(N__62361),
            .I(N__62227));
    LocalMux I__15420 (
            .O(N__62358),
            .I(N__62227));
    LocalMux I__15419 (
            .O(N__62355),
            .I(N__62218));
    LocalMux I__15418 (
            .O(N__62338),
            .I(N__62218));
    Span4Mux_v I__15417 (
            .O(N__62335),
            .I(N__62218));
    Span4Mux_h I__15416 (
            .O(N__62332),
            .I(N__62218));
    Span4Mux_h I__15415 (
            .O(N__62327),
            .I(N__62215));
    LocalMux I__15414 (
            .O(N__62324),
            .I(N__62212));
    Span4Mux_v I__15413 (
            .O(N__62321),
            .I(N__62205));
    LocalMux I__15412 (
            .O(N__62316),
            .I(N__62205));
    Span4Mux_h I__15411 (
            .O(N__62313),
            .I(N__62205));
    LocalMux I__15410 (
            .O(N__62308),
            .I(N__62200));
    Span4Mux_h I__15409 (
            .O(N__62301),
            .I(N__62200));
    LocalMux I__15408 (
            .O(N__62298),
            .I(N__62197));
    InMux I__15407 (
            .O(N__62297),
            .I(N__62192));
    InMux I__15406 (
            .O(N__62296),
            .I(N__62192));
    InMux I__15405 (
            .O(N__62295),
            .I(N__62187));
    InMux I__15404 (
            .O(N__62294),
            .I(N__62187));
    InMux I__15403 (
            .O(N__62293),
            .I(N__62184));
    InMux I__15402 (
            .O(N__62292),
            .I(N__62179));
    InMux I__15401 (
            .O(N__62291),
            .I(N__62179));
    InMux I__15400 (
            .O(N__62290),
            .I(N__62176));
    LocalMux I__15399 (
            .O(N__62285),
            .I(N__62171));
    Span12Mux_v I__15398 (
            .O(N__62276),
            .I(N__62171));
    Span4Mux_v I__15397 (
            .O(N__62273),
            .I(N__62164));
    LocalMux I__15396 (
            .O(N__62260),
            .I(N__62164));
    Span4Mux_v I__15395 (
            .O(N__62243),
            .I(N__62164));
    InMux I__15394 (
            .O(N__62242),
            .I(N__62157));
    InMux I__15393 (
            .O(N__62241),
            .I(N__62157));
    InMux I__15392 (
            .O(N__62240),
            .I(N__62157));
    Span4Mux_v I__15391 (
            .O(N__62237),
            .I(N__62154));
    LocalMux I__15390 (
            .O(N__62232),
            .I(N__62145));
    Span4Mux_h I__15389 (
            .O(N__62227),
            .I(N__62145));
    Span4Mux_v I__15388 (
            .O(N__62218),
            .I(N__62145));
    Span4Mux_h I__15387 (
            .O(N__62215),
            .I(N__62145));
    Span4Mux_h I__15386 (
            .O(N__62212),
            .I(N__62138));
    Span4Mux_h I__15385 (
            .O(N__62205),
            .I(N__62138));
    Span4Mux_h I__15384 (
            .O(N__62200),
            .I(N__62138));
    Odrv4 I__15383 (
            .O(N__62197),
            .I(comm_state_1));
    LocalMux I__15382 (
            .O(N__62192),
            .I(comm_state_1));
    LocalMux I__15381 (
            .O(N__62187),
            .I(comm_state_1));
    LocalMux I__15380 (
            .O(N__62184),
            .I(comm_state_1));
    LocalMux I__15379 (
            .O(N__62179),
            .I(comm_state_1));
    LocalMux I__15378 (
            .O(N__62176),
            .I(comm_state_1));
    Odrv12 I__15377 (
            .O(N__62171),
            .I(comm_state_1));
    Odrv4 I__15376 (
            .O(N__62164),
            .I(comm_state_1));
    LocalMux I__15375 (
            .O(N__62157),
            .I(comm_state_1));
    Odrv4 I__15374 (
            .O(N__62154),
            .I(comm_state_1));
    Odrv4 I__15373 (
            .O(N__62145),
            .I(comm_state_1));
    Odrv4 I__15372 (
            .O(N__62138),
            .I(comm_state_1));
    InMux I__15371 (
            .O(N__62113),
            .I(N__62110));
    LocalMux I__15370 (
            .O(N__62110),
            .I(N__62107));
    Span4Mux_h I__15369 (
            .O(N__62107),
            .I(N__62104));
    Odrv4 I__15368 (
            .O(N__62104),
            .I(comm_buf_0_7_N_543_3));
    CascadeMux I__15367 (
            .O(N__62101),
            .I(N__62097));
    CascadeMux I__15366 (
            .O(N__62100),
            .I(N__62094));
    InMux I__15365 (
            .O(N__62097),
            .I(N__62087));
    InMux I__15364 (
            .O(N__62094),
            .I(N__62087));
    InMux I__15363 (
            .O(N__62093),
            .I(N__62083));
    CascadeMux I__15362 (
            .O(N__62092),
            .I(N__62080));
    LocalMux I__15361 (
            .O(N__62087),
            .I(N__62076));
    InMux I__15360 (
            .O(N__62086),
            .I(N__62073));
    LocalMux I__15359 (
            .O(N__62083),
            .I(N__62070));
    InMux I__15358 (
            .O(N__62080),
            .I(N__62065));
    InMux I__15357 (
            .O(N__62079),
            .I(N__62065));
    Span4Mux_h I__15356 (
            .O(N__62076),
            .I(N__62060));
    LocalMux I__15355 (
            .O(N__62073),
            .I(N__62060));
    Span4Mux_v I__15354 (
            .O(N__62070),
            .I(N__62057));
    LocalMux I__15353 (
            .O(N__62065),
            .I(N__62053));
    Span4Mux_h I__15352 (
            .O(N__62060),
            .I(N__62050));
    Span4Mux_h I__15351 (
            .O(N__62057),
            .I(N__62047));
    InMux I__15350 (
            .O(N__62056),
            .I(N__62044));
    Span4Mux_v I__15349 (
            .O(N__62053),
            .I(N__62041));
    Span4Mux_h I__15348 (
            .O(N__62050),
            .I(N__62038));
    Span4Mux_h I__15347 (
            .O(N__62047),
            .I(N__62033));
    LocalMux I__15346 (
            .O(N__62044),
            .I(N__62033));
    Span4Mux_h I__15345 (
            .O(N__62041),
            .I(N__62030));
    Span4Mux_h I__15344 (
            .O(N__62038),
            .I(N__62025));
    Span4Mux_h I__15343 (
            .O(N__62033),
            .I(N__62025));
    Sp12to4 I__15342 (
            .O(N__62030),
            .I(N__62022));
    Span4Mux_v I__15341 (
            .O(N__62025),
            .I(N__62019));
    Odrv12 I__15340 (
            .O(N__62022),
            .I(comm_buf_0_3));
    Odrv4 I__15339 (
            .O(N__62019),
            .I(comm_buf_0_3));
    ClkMux I__15338 (
            .O(N__62014),
            .I(N__61441));
    ClkMux I__15337 (
            .O(N__62013),
            .I(N__61441));
    ClkMux I__15336 (
            .O(N__62012),
            .I(N__61441));
    ClkMux I__15335 (
            .O(N__62011),
            .I(N__61441));
    ClkMux I__15334 (
            .O(N__62010),
            .I(N__61441));
    ClkMux I__15333 (
            .O(N__62009),
            .I(N__61441));
    ClkMux I__15332 (
            .O(N__62008),
            .I(N__61441));
    ClkMux I__15331 (
            .O(N__62007),
            .I(N__61441));
    ClkMux I__15330 (
            .O(N__62006),
            .I(N__61441));
    ClkMux I__15329 (
            .O(N__62005),
            .I(N__61441));
    ClkMux I__15328 (
            .O(N__62004),
            .I(N__61441));
    ClkMux I__15327 (
            .O(N__62003),
            .I(N__61441));
    ClkMux I__15326 (
            .O(N__62002),
            .I(N__61441));
    ClkMux I__15325 (
            .O(N__62001),
            .I(N__61441));
    ClkMux I__15324 (
            .O(N__62000),
            .I(N__61441));
    ClkMux I__15323 (
            .O(N__61999),
            .I(N__61441));
    ClkMux I__15322 (
            .O(N__61998),
            .I(N__61441));
    ClkMux I__15321 (
            .O(N__61997),
            .I(N__61441));
    ClkMux I__15320 (
            .O(N__61996),
            .I(N__61441));
    ClkMux I__15319 (
            .O(N__61995),
            .I(N__61441));
    ClkMux I__15318 (
            .O(N__61994),
            .I(N__61441));
    ClkMux I__15317 (
            .O(N__61993),
            .I(N__61441));
    ClkMux I__15316 (
            .O(N__61992),
            .I(N__61441));
    ClkMux I__15315 (
            .O(N__61991),
            .I(N__61441));
    ClkMux I__15314 (
            .O(N__61990),
            .I(N__61441));
    ClkMux I__15313 (
            .O(N__61989),
            .I(N__61441));
    ClkMux I__15312 (
            .O(N__61988),
            .I(N__61441));
    ClkMux I__15311 (
            .O(N__61987),
            .I(N__61441));
    ClkMux I__15310 (
            .O(N__61986),
            .I(N__61441));
    ClkMux I__15309 (
            .O(N__61985),
            .I(N__61441));
    ClkMux I__15308 (
            .O(N__61984),
            .I(N__61441));
    ClkMux I__15307 (
            .O(N__61983),
            .I(N__61441));
    ClkMux I__15306 (
            .O(N__61982),
            .I(N__61441));
    ClkMux I__15305 (
            .O(N__61981),
            .I(N__61441));
    ClkMux I__15304 (
            .O(N__61980),
            .I(N__61441));
    ClkMux I__15303 (
            .O(N__61979),
            .I(N__61441));
    ClkMux I__15302 (
            .O(N__61978),
            .I(N__61441));
    ClkMux I__15301 (
            .O(N__61977),
            .I(N__61441));
    ClkMux I__15300 (
            .O(N__61976),
            .I(N__61441));
    ClkMux I__15299 (
            .O(N__61975),
            .I(N__61441));
    ClkMux I__15298 (
            .O(N__61974),
            .I(N__61441));
    ClkMux I__15297 (
            .O(N__61973),
            .I(N__61441));
    ClkMux I__15296 (
            .O(N__61972),
            .I(N__61441));
    ClkMux I__15295 (
            .O(N__61971),
            .I(N__61441));
    ClkMux I__15294 (
            .O(N__61970),
            .I(N__61441));
    ClkMux I__15293 (
            .O(N__61969),
            .I(N__61441));
    ClkMux I__15292 (
            .O(N__61968),
            .I(N__61441));
    ClkMux I__15291 (
            .O(N__61967),
            .I(N__61441));
    ClkMux I__15290 (
            .O(N__61966),
            .I(N__61441));
    ClkMux I__15289 (
            .O(N__61965),
            .I(N__61441));
    ClkMux I__15288 (
            .O(N__61964),
            .I(N__61441));
    ClkMux I__15287 (
            .O(N__61963),
            .I(N__61441));
    ClkMux I__15286 (
            .O(N__61962),
            .I(N__61441));
    ClkMux I__15285 (
            .O(N__61961),
            .I(N__61441));
    ClkMux I__15284 (
            .O(N__61960),
            .I(N__61441));
    ClkMux I__15283 (
            .O(N__61959),
            .I(N__61441));
    ClkMux I__15282 (
            .O(N__61958),
            .I(N__61441));
    ClkMux I__15281 (
            .O(N__61957),
            .I(N__61441));
    ClkMux I__15280 (
            .O(N__61956),
            .I(N__61441));
    ClkMux I__15279 (
            .O(N__61955),
            .I(N__61441));
    ClkMux I__15278 (
            .O(N__61954),
            .I(N__61441));
    ClkMux I__15277 (
            .O(N__61953),
            .I(N__61441));
    ClkMux I__15276 (
            .O(N__61952),
            .I(N__61441));
    ClkMux I__15275 (
            .O(N__61951),
            .I(N__61441));
    ClkMux I__15274 (
            .O(N__61950),
            .I(N__61441));
    ClkMux I__15273 (
            .O(N__61949),
            .I(N__61441));
    ClkMux I__15272 (
            .O(N__61948),
            .I(N__61441));
    ClkMux I__15271 (
            .O(N__61947),
            .I(N__61441));
    ClkMux I__15270 (
            .O(N__61946),
            .I(N__61441));
    ClkMux I__15269 (
            .O(N__61945),
            .I(N__61441));
    ClkMux I__15268 (
            .O(N__61944),
            .I(N__61441));
    ClkMux I__15267 (
            .O(N__61943),
            .I(N__61441));
    ClkMux I__15266 (
            .O(N__61942),
            .I(N__61441));
    ClkMux I__15265 (
            .O(N__61941),
            .I(N__61441));
    ClkMux I__15264 (
            .O(N__61940),
            .I(N__61441));
    ClkMux I__15263 (
            .O(N__61939),
            .I(N__61441));
    ClkMux I__15262 (
            .O(N__61938),
            .I(N__61441));
    ClkMux I__15261 (
            .O(N__61937),
            .I(N__61441));
    ClkMux I__15260 (
            .O(N__61936),
            .I(N__61441));
    ClkMux I__15259 (
            .O(N__61935),
            .I(N__61441));
    ClkMux I__15258 (
            .O(N__61934),
            .I(N__61441));
    ClkMux I__15257 (
            .O(N__61933),
            .I(N__61441));
    ClkMux I__15256 (
            .O(N__61932),
            .I(N__61441));
    ClkMux I__15255 (
            .O(N__61931),
            .I(N__61441));
    ClkMux I__15254 (
            .O(N__61930),
            .I(N__61441));
    ClkMux I__15253 (
            .O(N__61929),
            .I(N__61441));
    ClkMux I__15252 (
            .O(N__61928),
            .I(N__61441));
    ClkMux I__15251 (
            .O(N__61927),
            .I(N__61441));
    ClkMux I__15250 (
            .O(N__61926),
            .I(N__61441));
    ClkMux I__15249 (
            .O(N__61925),
            .I(N__61441));
    ClkMux I__15248 (
            .O(N__61924),
            .I(N__61441));
    ClkMux I__15247 (
            .O(N__61923),
            .I(N__61441));
    ClkMux I__15246 (
            .O(N__61922),
            .I(N__61441));
    ClkMux I__15245 (
            .O(N__61921),
            .I(N__61441));
    ClkMux I__15244 (
            .O(N__61920),
            .I(N__61441));
    ClkMux I__15243 (
            .O(N__61919),
            .I(N__61441));
    ClkMux I__15242 (
            .O(N__61918),
            .I(N__61441));
    ClkMux I__15241 (
            .O(N__61917),
            .I(N__61441));
    ClkMux I__15240 (
            .O(N__61916),
            .I(N__61441));
    ClkMux I__15239 (
            .O(N__61915),
            .I(N__61441));
    ClkMux I__15238 (
            .O(N__61914),
            .I(N__61441));
    ClkMux I__15237 (
            .O(N__61913),
            .I(N__61441));
    ClkMux I__15236 (
            .O(N__61912),
            .I(N__61441));
    ClkMux I__15235 (
            .O(N__61911),
            .I(N__61441));
    ClkMux I__15234 (
            .O(N__61910),
            .I(N__61441));
    ClkMux I__15233 (
            .O(N__61909),
            .I(N__61441));
    ClkMux I__15232 (
            .O(N__61908),
            .I(N__61441));
    ClkMux I__15231 (
            .O(N__61907),
            .I(N__61441));
    ClkMux I__15230 (
            .O(N__61906),
            .I(N__61441));
    ClkMux I__15229 (
            .O(N__61905),
            .I(N__61441));
    ClkMux I__15228 (
            .O(N__61904),
            .I(N__61441));
    ClkMux I__15227 (
            .O(N__61903),
            .I(N__61441));
    ClkMux I__15226 (
            .O(N__61902),
            .I(N__61441));
    ClkMux I__15225 (
            .O(N__61901),
            .I(N__61441));
    ClkMux I__15224 (
            .O(N__61900),
            .I(N__61441));
    ClkMux I__15223 (
            .O(N__61899),
            .I(N__61441));
    ClkMux I__15222 (
            .O(N__61898),
            .I(N__61441));
    ClkMux I__15221 (
            .O(N__61897),
            .I(N__61441));
    ClkMux I__15220 (
            .O(N__61896),
            .I(N__61441));
    ClkMux I__15219 (
            .O(N__61895),
            .I(N__61441));
    ClkMux I__15218 (
            .O(N__61894),
            .I(N__61441));
    ClkMux I__15217 (
            .O(N__61893),
            .I(N__61441));
    ClkMux I__15216 (
            .O(N__61892),
            .I(N__61441));
    ClkMux I__15215 (
            .O(N__61891),
            .I(N__61441));
    ClkMux I__15214 (
            .O(N__61890),
            .I(N__61441));
    ClkMux I__15213 (
            .O(N__61889),
            .I(N__61441));
    ClkMux I__15212 (
            .O(N__61888),
            .I(N__61441));
    ClkMux I__15211 (
            .O(N__61887),
            .I(N__61441));
    ClkMux I__15210 (
            .O(N__61886),
            .I(N__61441));
    ClkMux I__15209 (
            .O(N__61885),
            .I(N__61441));
    ClkMux I__15208 (
            .O(N__61884),
            .I(N__61441));
    ClkMux I__15207 (
            .O(N__61883),
            .I(N__61441));
    ClkMux I__15206 (
            .O(N__61882),
            .I(N__61441));
    ClkMux I__15205 (
            .O(N__61881),
            .I(N__61441));
    ClkMux I__15204 (
            .O(N__61880),
            .I(N__61441));
    ClkMux I__15203 (
            .O(N__61879),
            .I(N__61441));
    ClkMux I__15202 (
            .O(N__61878),
            .I(N__61441));
    ClkMux I__15201 (
            .O(N__61877),
            .I(N__61441));
    ClkMux I__15200 (
            .O(N__61876),
            .I(N__61441));
    ClkMux I__15199 (
            .O(N__61875),
            .I(N__61441));
    ClkMux I__15198 (
            .O(N__61874),
            .I(N__61441));
    ClkMux I__15197 (
            .O(N__61873),
            .I(N__61441));
    ClkMux I__15196 (
            .O(N__61872),
            .I(N__61441));
    ClkMux I__15195 (
            .O(N__61871),
            .I(N__61441));
    ClkMux I__15194 (
            .O(N__61870),
            .I(N__61441));
    ClkMux I__15193 (
            .O(N__61869),
            .I(N__61441));
    ClkMux I__15192 (
            .O(N__61868),
            .I(N__61441));
    ClkMux I__15191 (
            .O(N__61867),
            .I(N__61441));
    ClkMux I__15190 (
            .O(N__61866),
            .I(N__61441));
    ClkMux I__15189 (
            .O(N__61865),
            .I(N__61441));
    ClkMux I__15188 (
            .O(N__61864),
            .I(N__61441));
    ClkMux I__15187 (
            .O(N__61863),
            .I(N__61441));
    ClkMux I__15186 (
            .O(N__61862),
            .I(N__61441));
    ClkMux I__15185 (
            .O(N__61861),
            .I(N__61441));
    ClkMux I__15184 (
            .O(N__61860),
            .I(N__61441));
    ClkMux I__15183 (
            .O(N__61859),
            .I(N__61441));
    ClkMux I__15182 (
            .O(N__61858),
            .I(N__61441));
    ClkMux I__15181 (
            .O(N__61857),
            .I(N__61441));
    ClkMux I__15180 (
            .O(N__61856),
            .I(N__61441));
    ClkMux I__15179 (
            .O(N__61855),
            .I(N__61441));
    ClkMux I__15178 (
            .O(N__61854),
            .I(N__61441));
    ClkMux I__15177 (
            .O(N__61853),
            .I(N__61441));
    ClkMux I__15176 (
            .O(N__61852),
            .I(N__61441));
    ClkMux I__15175 (
            .O(N__61851),
            .I(N__61441));
    ClkMux I__15174 (
            .O(N__61850),
            .I(N__61441));
    ClkMux I__15173 (
            .O(N__61849),
            .I(N__61441));
    ClkMux I__15172 (
            .O(N__61848),
            .I(N__61441));
    ClkMux I__15171 (
            .O(N__61847),
            .I(N__61441));
    ClkMux I__15170 (
            .O(N__61846),
            .I(N__61441));
    ClkMux I__15169 (
            .O(N__61845),
            .I(N__61441));
    ClkMux I__15168 (
            .O(N__61844),
            .I(N__61441));
    ClkMux I__15167 (
            .O(N__61843),
            .I(N__61441));
    ClkMux I__15166 (
            .O(N__61842),
            .I(N__61441));
    ClkMux I__15165 (
            .O(N__61841),
            .I(N__61441));
    ClkMux I__15164 (
            .O(N__61840),
            .I(N__61441));
    ClkMux I__15163 (
            .O(N__61839),
            .I(N__61441));
    ClkMux I__15162 (
            .O(N__61838),
            .I(N__61441));
    ClkMux I__15161 (
            .O(N__61837),
            .I(N__61441));
    ClkMux I__15160 (
            .O(N__61836),
            .I(N__61441));
    ClkMux I__15159 (
            .O(N__61835),
            .I(N__61441));
    ClkMux I__15158 (
            .O(N__61834),
            .I(N__61441));
    ClkMux I__15157 (
            .O(N__61833),
            .I(N__61441));
    ClkMux I__15156 (
            .O(N__61832),
            .I(N__61441));
    ClkMux I__15155 (
            .O(N__61831),
            .I(N__61441));
    ClkMux I__15154 (
            .O(N__61830),
            .I(N__61441));
    ClkMux I__15153 (
            .O(N__61829),
            .I(N__61441));
    ClkMux I__15152 (
            .O(N__61828),
            .I(N__61441));
    ClkMux I__15151 (
            .O(N__61827),
            .I(N__61441));
    ClkMux I__15150 (
            .O(N__61826),
            .I(N__61441));
    ClkMux I__15149 (
            .O(N__61825),
            .I(N__61441));
    ClkMux I__15148 (
            .O(N__61824),
            .I(N__61441));
    GlobalMux I__15147 (
            .O(N__61441),
            .I(clk_32MHz));
    CEMux I__15146 (
            .O(N__61438),
            .I(N__61434));
    CEMux I__15145 (
            .O(N__61437),
            .I(N__61431));
    LocalMux I__15144 (
            .O(N__61434),
            .I(N__61428));
    LocalMux I__15143 (
            .O(N__61431),
            .I(N__61425));
    Span4Mux_h I__15142 (
            .O(N__61428),
            .I(N__61420));
    Span4Mux_h I__15141 (
            .O(N__61425),
            .I(N__61420));
    Odrv4 I__15140 (
            .O(N__61420),
            .I(n12677));
    CascadeMux I__15139 (
            .O(N__61417),
            .I(n30_adj_1793_cascade_));
    CascadeMux I__15138 (
            .O(N__61414),
            .I(N__61402));
    CascadeMux I__15137 (
            .O(N__61413),
            .I(N__61391));
    InMux I__15136 (
            .O(N__61412),
            .I(N__61387));
    InMux I__15135 (
            .O(N__61411),
            .I(N__61384));
    InMux I__15134 (
            .O(N__61410),
            .I(N__61376));
    InMux I__15133 (
            .O(N__61409),
            .I(N__61370));
    InMux I__15132 (
            .O(N__61408),
            .I(N__61367));
    InMux I__15131 (
            .O(N__61407),
            .I(N__61364));
    InMux I__15130 (
            .O(N__61406),
            .I(N__61359));
    InMux I__15129 (
            .O(N__61405),
            .I(N__61356));
    InMux I__15128 (
            .O(N__61402),
            .I(N__61353));
    InMux I__15127 (
            .O(N__61401),
            .I(N__61349));
    InMux I__15126 (
            .O(N__61400),
            .I(N__61344));
    InMux I__15125 (
            .O(N__61399),
            .I(N__61339));
    InMux I__15124 (
            .O(N__61398),
            .I(N__61339));
    InMux I__15123 (
            .O(N__61397),
            .I(N__61336));
    InMux I__15122 (
            .O(N__61396),
            .I(N__61333));
    InMux I__15121 (
            .O(N__61395),
            .I(N__61330));
    InMux I__15120 (
            .O(N__61394),
            .I(N__61327));
    InMux I__15119 (
            .O(N__61391),
            .I(N__61322));
    InMux I__15118 (
            .O(N__61390),
            .I(N__61322));
    LocalMux I__15117 (
            .O(N__61387),
            .I(N__61319));
    LocalMux I__15116 (
            .O(N__61384),
            .I(N__61316));
    InMux I__15115 (
            .O(N__61383),
            .I(N__61313));
    InMux I__15114 (
            .O(N__61382),
            .I(N__61310));
    InMux I__15113 (
            .O(N__61381),
            .I(N__61307));
    InMux I__15112 (
            .O(N__61380),
            .I(N__61304));
    InMux I__15111 (
            .O(N__61379),
            .I(N__61301));
    LocalMux I__15110 (
            .O(N__61376),
            .I(N__61297));
    InMux I__15109 (
            .O(N__61375),
            .I(N__61292));
    InMux I__15108 (
            .O(N__61374),
            .I(N__61292));
    InMux I__15107 (
            .O(N__61373),
            .I(N__61288));
    LocalMux I__15106 (
            .O(N__61370),
            .I(N__61281));
    LocalMux I__15105 (
            .O(N__61367),
            .I(N__61281));
    LocalMux I__15104 (
            .O(N__61364),
            .I(N__61281));
    InMux I__15103 (
            .O(N__61363),
            .I(N__61276));
    InMux I__15102 (
            .O(N__61362),
            .I(N__61276));
    LocalMux I__15101 (
            .O(N__61359),
            .I(N__61269));
    LocalMux I__15100 (
            .O(N__61356),
            .I(N__61269));
    LocalMux I__15099 (
            .O(N__61353),
            .I(N__61269));
    InMux I__15098 (
            .O(N__61352),
            .I(N__61264));
    LocalMux I__15097 (
            .O(N__61349),
            .I(N__61261));
    InMux I__15096 (
            .O(N__61348),
            .I(N__61255));
    InMux I__15095 (
            .O(N__61347),
            .I(N__61255));
    LocalMux I__15094 (
            .O(N__61344),
            .I(N__61248));
    LocalMux I__15093 (
            .O(N__61339),
            .I(N__61248));
    LocalMux I__15092 (
            .O(N__61336),
            .I(N__61245));
    LocalMux I__15091 (
            .O(N__61333),
            .I(N__61242));
    LocalMux I__15090 (
            .O(N__61330),
            .I(N__61233));
    LocalMux I__15089 (
            .O(N__61327),
            .I(N__61233));
    LocalMux I__15088 (
            .O(N__61322),
            .I(N__61233));
    Span4Mux_v I__15087 (
            .O(N__61319),
            .I(N__61233));
    Span4Mux_h I__15086 (
            .O(N__61316),
            .I(N__61226));
    LocalMux I__15085 (
            .O(N__61313),
            .I(N__61226));
    LocalMux I__15084 (
            .O(N__61310),
            .I(N__61223));
    LocalMux I__15083 (
            .O(N__61307),
            .I(N__61218));
    LocalMux I__15082 (
            .O(N__61304),
            .I(N__61218));
    LocalMux I__15081 (
            .O(N__61301),
            .I(N__61215));
    InMux I__15080 (
            .O(N__61300),
            .I(N__61212));
    Span4Mux_v I__15079 (
            .O(N__61297),
            .I(N__61207));
    LocalMux I__15078 (
            .O(N__61292),
            .I(N__61207));
    InMux I__15077 (
            .O(N__61291),
            .I(N__61204));
    LocalMux I__15076 (
            .O(N__61288),
            .I(N__61201));
    Span4Mux_v I__15075 (
            .O(N__61281),
            .I(N__61194));
    LocalMux I__15074 (
            .O(N__61276),
            .I(N__61194));
    Span4Mux_h I__15073 (
            .O(N__61269),
            .I(N__61194));
    InMux I__15072 (
            .O(N__61268),
            .I(N__61189));
    InMux I__15071 (
            .O(N__61267),
            .I(N__61189));
    LocalMux I__15070 (
            .O(N__61264),
            .I(N__61184));
    Span4Mux_h I__15069 (
            .O(N__61261),
            .I(N__61184));
    CascadeMux I__15068 (
            .O(N__61260),
            .I(N__61179));
    LocalMux I__15067 (
            .O(N__61255),
            .I(N__61175));
    InMux I__15066 (
            .O(N__61254),
            .I(N__61172));
    InMux I__15065 (
            .O(N__61253),
            .I(N__61169));
    Span4Mux_v I__15064 (
            .O(N__61248),
            .I(N__61160));
    Span4Mux_v I__15063 (
            .O(N__61245),
            .I(N__61160));
    Span4Mux_v I__15062 (
            .O(N__61242),
            .I(N__61160));
    Span4Mux_h I__15061 (
            .O(N__61233),
            .I(N__61160));
    InMux I__15060 (
            .O(N__61232),
            .I(N__61157));
    InMux I__15059 (
            .O(N__61231),
            .I(N__61154));
    Span4Mux_v I__15058 (
            .O(N__61226),
            .I(N__61141));
    Span4Mux_v I__15057 (
            .O(N__61223),
            .I(N__61141));
    Span4Mux_v I__15056 (
            .O(N__61218),
            .I(N__61141));
    Span4Mux_h I__15055 (
            .O(N__61215),
            .I(N__61141));
    LocalMux I__15054 (
            .O(N__61212),
            .I(N__61141));
    Span4Mux_h I__15053 (
            .O(N__61207),
            .I(N__61141));
    LocalMux I__15052 (
            .O(N__61204),
            .I(N__61130));
    Span4Mux_v I__15051 (
            .O(N__61201),
            .I(N__61130));
    Span4Mux_h I__15050 (
            .O(N__61194),
            .I(N__61130));
    LocalMux I__15049 (
            .O(N__61189),
            .I(N__61130));
    Span4Mux_h I__15048 (
            .O(N__61184),
            .I(N__61130));
    InMux I__15047 (
            .O(N__61183),
            .I(N__61121));
    InMux I__15046 (
            .O(N__61182),
            .I(N__61121));
    InMux I__15045 (
            .O(N__61179),
            .I(N__61121));
    InMux I__15044 (
            .O(N__61178),
            .I(N__61121));
    Odrv12 I__15043 (
            .O(N__61175),
            .I(comm_cmd_6));
    LocalMux I__15042 (
            .O(N__61172),
            .I(comm_cmd_6));
    LocalMux I__15041 (
            .O(N__61169),
            .I(comm_cmd_6));
    Odrv4 I__15040 (
            .O(N__61160),
            .I(comm_cmd_6));
    LocalMux I__15039 (
            .O(N__61157),
            .I(comm_cmd_6));
    LocalMux I__15038 (
            .O(N__61154),
            .I(comm_cmd_6));
    Odrv4 I__15037 (
            .O(N__61141),
            .I(comm_cmd_6));
    Odrv4 I__15036 (
            .O(N__61130),
            .I(comm_cmd_6));
    LocalMux I__15035 (
            .O(N__61121),
            .I(comm_cmd_6));
    CascadeMux I__15034 (
            .O(N__61102),
            .I(N__61099));
    InMux I__15033 (
            .O(N__61099),
            .I(N__61096));
    LocalMux I__15032 (
            .O(N__61096),
            .I(N__61092));
    CascadeMux I__15031 (
            .O(N__61095),
            .I(N__61089));
    Span4Mux_v I__15030 (
            .O(N__61092),
            .I(N__61086));
    InMux I__15029 (
            .O(N__61089),
            .I(N__61083));
    Span4Mux_h I__15028 (
            .O(N__61086),
            .I(N__61080));
    LocalMux I__15027 (
            .O(N__61083),
            .I(data_idxvec_13));
    Odrv4 I__15026 (
            .O(N__61080),
            .I(data_idxvec_13));
    InMux I__15025 (
            .O(N__61075),
            .I(N__61072));
    LocalMux I__15024 (
            .O(N__61072),
            .I(N__61069));
    Span4Mux_v I__15023 (
            .O(N__61069),
            .I(N__61066));
    Span4Mux_v I__15022 (
            .O(N__61066),
            .I(N__61063));
    Odrv4 I__15021 (
            .O(N__61063),
            .I(buf_data_iac_21));
    CascadeMux I__15020 (
            .O(N__61060),
            .I(n28_adj_1775_cascade_));
    CascadeMux I__15019 (
            .O(N__61057),
            .I(N__61048));
    InMux I__15018 (
            .O(N__61056),
            .I(N__61045));
    InMux I__15017 (
            .O(N__61055),
            .I(N__61042));
    InMux I__15016 (
            .O(N__61054),
            .I(N__61037));
    InMux I__15015 (
            .O(N__61053),
            .I(N__61037));
    InMux I__15014 (
            .O(N__61052),
            .I(N__61029));
    InMux I__15013 (
            .O(N__61051),
            .I(N__61026));
    InMux I__15012 (
            .O(N__61048),
            .I(N__61014));
    LocalMux I__15011 (
            .O(N__61045),
            .I(N__61010));
    LocalMux I__15010 (
            .O(N__61042),
            .I(N__61007));
    LocalMux I__15009 (
            .O(N__61037),
            .I(N__61004));
    InMux I__15008 (
            .O(N__61036),
            .I(N__60995));
    InMux I__15007 (
            .O(N__61035),
            .I(N__60995));
    InMux I__15006 (
            .O(N__61034),
            .I(N__60995));
    InMux I__15005 (
            .O(N__61033),
            .I(N__60995));
    InMux I__15004 (
            .O(N__61032),
            .I(N__60986));
    LocalMux I__15003 (
            .O(N__61029),
            .I(N__60981));
    LocalMux I__15002 (
            .O(N__61026),
            .I(N__60981));
    InMux I__15001 (
            .O(N__61025),
            .I(N__60970));
    InMux I__15000 (
            .O(N__61024),
            .I(N__60970));
    InMux I__14999 (
            .O(N__61023),
            .I(N__60963));
    InMux I__14998 (
            .O(N__61022),
            .I(N__60963));
    InMux I__14997 (
            .O(N__61021),
            .I(N__60963));
    InMux I__14996 (
            .O(N__61020),
            .I(N__60958));
    InMux I__14995 (
            .O(N__61019),
            .I(N__60958));
    CascadeMux I__14994 (
            .O(N__61018),
            .I(N__60949));
    InMux I__14993 (
            .O(N__61017),
            .I(N__60945));
    LocalMux I__14992 (
            .O(N__61014),
            .I(N__60942));
    InMux I__14991 (
            .O(N__61013),
            .I(N__60939));
    Span4Mux_v I__14990 (
            .O(N__61010),
            .I(N__60932));
    Span4Mux_v I__14989 (
            .O(N__61007),
            .I(N__60932));
    Span4Mux_h I__14988 (
            .O(N__61004),
            .I(N__60932));
    LocalMux I__14987 (
            .O(N__60995),
            .I(N__60929));
    InMux I__14986 (
            .O(N__60994),
            .I(N__60926));
    InMux I__14985 (
            .O(N__60993),
            .I(N__60921));
    InMux I__14984 (
            .O(N__60992),
            .I(N__60921));
    InMux I__14983 (
            .O(N__60991),
            .I(N__60918));
    InMux I__14982 (
            .O(N__60990),
            .I(N__60915));
    InMux I__14981 (
            .O(N__60989),
            .I(N__60912));
    LocalMux I__14980 (
            .O(N__60986),
            .I(N__60909));
    Span4Mux_v I__14979 (
            .O(N__60981),
            .I(N__60906));
    InMux I__14978 (
            .O(N__60980),
            .I(N__60903));
    InMux I__14977 (
            .O(N__60979),
            .I(N__60899));
    InMux I__14976 (
            .O(N__60978),
            .I(N__60894));
    InMux I__14975 (
            .O(N__60977),
            .I(N__60894));
    InMux I__14974 (
            .O(N__60976),
            .I(N__60889));
    InMux I__14973 (
            .O(N__60975),
            .I(N__60889));
    LocalMux I__14972 (
            .O(N__60970),
            .I(N__60884));
    LocalMux I__14971 (
            .O(N__60963),
            .I(N__60884));
    LocalMux I__14970 (
            .O(N__60958),
            .I(N__60881));
    InMux I__14969 (
            .O(N__60957),
            .I(N__60876));
    InMux I__14968 (
            .O(N__60956),
            .I(N__60871));
    InMux I__14967 (
            .O(N__60955),
            .I(N__60871));
    InMux I__14966 (
            .O(N__60954),
            .I(N__60866));
    InMux I__14965 (
            .O(N__60953),
            .I(N__60866));
    InMux I__14964 (
            .O(N__60952),
            .I(N__60862));
    InMux I__14963 (
            .O(N__60949),
            .I(N__60859));
    InMux I__14962 (
            .O(N__60948),
            .I(N__60856));
    LocalMux I__14961 (
            .O(N__60945),
            .I(N__60853));
    Span12Mux_v I__14960 (
            .O(N__60942),
            .I(N__60850));
    LocalMux I__14959 (
            .O(N__60939),
            .I(N__60847));
    Span4Mux_h I__14958 (
            .O(N__60932),
            .I(N__60842));
    Span4Mux_h I__14957 (
            .O(N__60929),
            .I(N__60842));
    LocalMux I__14956 (
            .O(N__60926),
            .I(N__60837));
    LocalMux I__14955 (
            .O(N__60921),
            .I(N__60837));
    LocalMux I__14954 (
            .O(N__60918),
            .I(N__60834));
    LocalMux I__14953 (
            .O(N__60915),
            .I(N__60831));
    LocalMux I__14952 (
            .O(N__60912),
            .I(N__60822));
    Span4Mux_v I__14951 (
            .O(N__60909),
            .I(N__60822));
    Span4Mux_h I__14950 (
            .O(N__60906),
            .I(N__60822));
    LocalMux I__14949 (
            .O(N__60903),
            .I(N__60822));
    InMux I__14948 (
            .O(N__60902),
            .I(N__60819));
    LocalMux I__14947 (
            .O(N__60899),
            .I(N__60810));
    LocalMux I__14946 (
            .O(N__60894),
            .I(N__60810));
    LocalMux I__14945 (
            .O(N__60889),
            .I(N__60810));
    Span4Mux_v I__14944 (
            .O(N__60884),
            .I(N__60810));
    Span4Mux_h I__14943 (
            .O(N__60881),
            .I(N__60807));
    InMux I__14942 (
            .O(N__60880),
            .I(N__60804));
    InMux I__14941 (
            .O(N__60879),
            .I(N__60801));
    LocalMux I__14940 (
            .O(N__60876),
            .I(N__60794));
    LocalMux I__14939 (
            .O(N__60871),
            .I(N__60794));
    LocalMux I__14938 (
            .O(N__60866),
            .I(N__60794));
    InMux I__14937 (
            .O(N__60865),
            .I(N__60789));
    LocalMux I__14936 (
            .O(N__60862),
            .I(N__60786));
    LocalMux I__14935 (
            .O(N__60859),
            .I(N__60781));
    LocalMux I__14934 (
            .O(N__60856),
            .I(N__60781));
    Span12Mux_h I__14933 (
            .O(N__60853),
            .I(N__60778));
    Span12Mux_h I__14932 (
            .O(N__60850),
            .I(N__60775));
    Span4Mux_h I__14931 (
            .O(N__60847),
            .I(N__60770));
    Span4Mux_h I__14930 (
            .O(N__60842),
            .I(N__60770));
    Span4Mux_v I__14929 (
            .O(N__60837),
            .I(N__60757));
    Span4Mux_v I__14928 (
            .O(N__60834),
            .I(N__60757));
    Span4Mux_v I__14927 (
            .O(N__60831),
            .I(N__60757));
    Span4Mux_h I__14926 (
            .O(N__60822),
            .I(N__60757));
    LocalMux I__14925 (
            .O(N__60819),
            .I(N__60757));
    Span4Mux_v I__14924 (
            .O(N__60810),
            .I(N__60757));
    Span4Mux_h I__14923 (
            .O(N__60807),
            .I(N__60750));
    LocalMux I__14922 (
            .O(N__60804),
            .I(N__60750));
    LocalMux I__14921 (
            .O(N__60801),
            .I(N__60750));
    Span4Mux_v I__14920 (
            .O(N__60794),
            .I(N__60747));
    InMux I__14919 (
            .O(N__60793),
            .I(N__60742));
    InMux I__14918 (
            .O(N__60792),
            .I(N__60742));
    LocalMux I__14917 (
            .O(N__60789),
            .I(comm_cmd_3));
    Odrv4 I__14916 (
            .O(N__60786),
            .I(comm_cmd_3));
    Odrv12 I__14915 (
            .O(N__60781),
            .I(comm_cmd_3));
    Odrv12 I__14914 (
            .O(N__60778),
            .I(comm_cmd_3));
    Odrv12 I__14913 (
            .O(N__60775),
            .I(comm_cmd_3));
    Odrv4 I__14912 (
            .O(N__60770),
            .I(comm_cmd_3));
    Odrv4 I__14911 (
            .O(N__60757),
            .I(comm_cmd_3));
    Odrv4 I__14910 (
            .O(N__60750),
            .I(comm_cmd_3));
    Odrv4 I__14909 (
            .O(N__60747),
            .I(comm_cmd_3));
    LocalMux I__14908 (
            .O(N__60742),
            .I(comm_cmd_3));
    InMux I__14907 (
            .O(N__60721),
            .I(N__60718));
    LocalMux I__14906 (
            .O(N__60718),
            .I(N__60715));
    Odrv4 I__14905 (
            .O(N__60715),
            .I(n23492));
    CascadeMux I__14904 (
            .O(N__60712),
            .I(N__60709));
    InMux I__14903 (
            .O(N__60709),
            .I(N__60706));
    LocalMux I__14902 (
            .O(N__60706),
            .I(N__60703));
    Sp12to4 I__14901 (
            .O(N__60703),
            .I(N__60700));
    Odrv12 I__14900 (
            .O(N__60700),
            .I(n23_adj_1773));
    InMux I__14899 (
            .O(N__60697),
            .I(N__60694));
    LocalMux I__14898 (
            .O(N__60694),
            .I(N__60691));
    Span12Mux_h I__14897 (
            .O(N__60691),
            .I(N__60686));
    InMux I__14896 (
            .O(N__60690),
            .I(N__60681));
    InMux I__14895 (
            .O(N__60689),
            .I(N__60681));
    Odrv12 I__14894 (
            .O(N__60686),
            .I(req_data_cnt_13));
    LocalMux I__14893 (
            .O(N__60681),
            .I(req_data_cnt_13));
    InMux I__14892 (
            .O(N__60676),
            .I(N__60673));
    LocalMux I__14891 (
            .O(N__60673),
            .I(n25_adj_1774));
    InMux I__14890 (
            .O(N__60670),
            .I(N__60660));
    InMux I__14889 (
            .O(N__60669),
            .I(N__60657));
    InMux I__14888 (
            .O(N__60668),
            .I(N__60650));
    InMux I__14887 (
            .O(N__60667),
            .I(N__60650));
    InMux I__14886 (
            .O(N__60666),
            .I(N__60650));
    InMux I__14885 (
            .O(N__60665),
            .I(N__60643));
    InMux I__14884 (
            .O(N__60664),
            .I(N__60637));
    CascadeMux I__14883 (
            .O(N__60663),
            .I(N__60632));
    LocalMux I__14882 (
            .O(N__60660),
            .I(N__60628));
    LocalMux I__14881 (
            .O(N__60657),
            .I(N__60624));
    LocalMux I__14880 (
            .O(N__60650),
            .I(N__60621));
    InMux I__14879 (
            .O(N__60649),
            .I(N__60616));
    InMux I__14878 (
            .O(N__60648),
            .I(N__60612));
    InMux I__14877 (
            .O(N__60647),
            .I(N__60604));
    InMux I__14876 (
            .O(N__60646),
            .I(N__60604));
    LocalMux I__14875 (
            .O(N__60643),
            .I(N__60584));
    InMux I__14874 (
            .O(N__60642),
            .I(N__60579));
    InMux I__14873 (
            .O(N__60641),
            .I(N__60579));
    InMux I__14872 (
            .O(N__60640),
            .I(N__60576));
    LocalMux I__14871 (
            .O(N__60637),
            .I(N__60573));
    InMux I__14870 (
            .O(N__60636),
            .I(N__60568));
    InMux I__14869 (
            .O(N__60635),
            .I(N__60568));
    InMux I__14868 (
            .O(N__60632),
            .I(N__60565));
    InMux I__14867 (
            .O(N__60631),
            .I(N__60561));
    Span4Mux_h I__14866 (
            .O(N__60628),
            .I(N__60558));
    InMux I__14865 (
            .O(N__60627),
            .I(N__60555));
    Span4Mux_h I__14864 (
            .O(N__60624),
            .I(N__60550));
    Span4Mux_h I__14863 (
            .O(N__60621),
            .I(N__60550));
    InMux I__14862 (
            .O(N__60620),
            .I(N__60547));
    InMux I__14861 (
            .O(N__60619),
            .I(N__60540));
    LocalMux I__14860 (
            .O(N__60616),
            .I(N__60537));
    InMux I__14859 (
            .O(N__60615),
            .I(N__60534));
    LocalMux I__14858 (
            .O(N__60612),
            .I(N__60531));
    InMux I__14857 (
            .O(N__60611),
            .I(N__60528));
    InMux I__14856 (
            .O(N__60610),
            .I(N__60523));
    InMux I__14855 (
            .O(N__60609),
            .I(N__60523));
    LocalMux I__14854 (
            .O(N__60604),
            .I(N__60513));
    InMux I__14853 (
            .O(N__60603),
            .I(N__60510));
    InMux I__14852 (
            .O(N__60602),
            .I(N__60507));
    InMux I__14851 (
            .O(N__60601),
            .I(N__60502));
    InMux I__14850 (
            .O(N__60600),
            .I(N__60502));
    InMux I__14849 (
            .O(N__60599),
            .I(N__60490));
    InMux I__14848 (
            .O(N__60598),
            .I(N__60490));
    InMux I__14847 (
            .O(N__60597),
            .I(N__60487));
    InMux I__14846 (
            .O(N__60596),
            .I(N__60480));
    InMux I__14845 (
            .O(N__60595),
            .I(N__60480));
    InMux I__14844 (
            .O(N__60594),
            .I(N__60480));
    InMux I__14843 (
            .O(N__60593),
            .I(N__60475));
    InMux I__14842 (
            .O(N__60592),
            .I(N__60470));
    InMux I__14841 (
            .O(N__60591),
            .I(N__60470));
    InMux I__14840 (
            .O(N__60590),
            .I(N__60464));
    InMux I__14839 (
            .O(N__60589),
            .I(N__60458));
    InMux I__14838 (
            .O(N__60588),
            .I(N__60453));
    InMux I__14837 (
            .O(N__60587),
            .I(N__60453));
    Span4Mux_h I__14836 (
            .O(N__60584),
            .I(N__60446));
    LocalMux I__14835 (
            .O(N__60579),
            .I(N__60446));
    LocalMux I__14834 (
            .O(N__60576),
            .I(N__60446));
    Span4Mux_v I__14833 (
            .O(N__60573),
            .I(N__60439));
    LocalMux I__14832 (
            .O(N__60568),
            .I(N__60439));
    LocalMux I__14831 (
            .O(N__60565),
            .I(N__60439));
    InMux I__14830 (
            .O(N__60564),
            .I(N__60436));
    LocalMux I__14829 (
            .O(N__60561),
            .I(N__60433));
    Span4Mux_h I__14828 (
            .O(N__60558),
            .I(N__60426));
    LocalMux I__14827 (
            .O(N__60555),
            .I(N__60426));
    Span4Mux_h I__14826 (
            .O(N__60550),
            .I(N__60426));
    LocalMux I__14825 (
            .O(N__60547),
            .I(N__60423));
    InMux I__14824 (
            .O(N__60546),
            .I(N__60416));
    InMux I__14823 (
            .O(N__60545),
            .I(N__60416));
    InMux I__14822 (
            .O(N__60544),
            .I(N__60416));
    InMux I__14821 (
            .O(N__60543),
            .I(N__60413));
    LocalMux I__14820 (
            .O(N__60540),
            .I(N__60410));
    Span4Mux_v I__14819 (
            .O(N__60537),
            .I(N__60407));
    LocalMux I__14818 (
            .O(N__60534),
            .I(N__60398));
    Span4Mux_v I__14817 (
            .O(N__60531),
            .I(N__60398));
    LocalMux I__14816 (
            .O(N__60528),
            .I(N__60398));
    LocalMux I__14815 (
            .O(N__60523),
            .I(N__60398));
    InMux I__14814 (
            .O(N__60522),
            .I(N__60392));
    InMux I__14813 (
            .O(N__60521),
            .I(N__60389));
    InMux I__14812 (
            .O(N__60520),
            .I(N__60386));
    InMux I__14811 (
            .O(N__60519),
            .I(N__60381));
    InMux I__14810 (
            .O(N__60518),
            .I(N__60381));
    InMux I__14809 (
            .O(N__60517),
            .I(N__60376));
    InMux I__14808 (
            .O(N__60516),
            .I(N__60376));
    Span4Mux_h I__14807 (
            .O(N__60513),
            .I(N__60371));
    LocalMux I__14806 (
            .O(N__60510),
            .I(N__60371));
    LocalMux I__14805 (
            .O(N__60507),
            .I(N__60366));
    LocalMux I__14804 (
            .O(N__60502),
            .I(N__60366));
    InMux I__14803 (
            .O(N__60501),
            .I(N__60359));
    InMux I__14802 (
            .O(N__60500),
            .I(N__60359));
    InMux I__14801 (
            .O(N__60499),
            .I(N__60359));
    InMux I__14800 (
            .O(N__60498),
            .I(N__60354));
    InMux I__14799 (
            .O(N__60497),
            .I(N__60349));
    InMux I__14798 (
            .O(N__60496),
            .I(N__60344));
    InMux I__14797 (
            .O(N__60495),
            .I(N__60344));
    LocalMux I__14796 (
            .O(N__60490),
            .I(N__60341));
    LocalMux I__14795 (
            .O(N__60487),
            .I(N__60336));
    LocalMux I__14794 (
            .O(N__60480),
            .I(N__60336));
    InMux I__14793 (
            .O(N__60479),
            .I(N__60331));
    InMux I__14792 (
            .O(N__60478),
            .I(N__60331));
    LocalMux I__14791 (
            .O(N__60475),
            .I(N__60326));
    LocalMux I__14790 (
            .O(N__60470),
            .I(N__60326));
    InMux I__14789 (
            .O(N__60469),
            .I(N__60321));
    InMux I__14788 (
            .O(N__60468),
            .I(N__60321));
    InMux I__14787 (
            .O(N__60467),
            .I(N__60318));
    LocalMux I__14786 (
            .O(N__60464),
            .I(N__60315));
    CascadeMux I__14785 (
            .O(N__60463),
            .I(N__60310));
    InMux I__14784 (
            .O(N__60462),
            .I(N__60304));
    InMux I__14783 (
            .O(N__60461),
            .I(N__60304));
    LocalMux I__14782 (
            .O(N__60458),
            .I(N__60301));
    LocalMux I__14781 (
            .O(N__60453),
            .I(N__60294));
    Span4Mux_h I__14780 (
            .O(N__60446),
            .I(N__60294));
    Span4Mux_h I__14779 (
            .O(N__60439),
            .I(N__60294));
    LocalMux I__14778 (
            .O(N__60436),
            .I(N__60285));
    Span4Mux_h I__14777 (
            .O(N__60433),
            .I(N__60285));
    Span4Mux_v I__14776 (
            .O(N__60426),
            .I(N__60285));
    Span4Mux_h I__14775 (
            .O(N__60423),
            .I(N__60285));
    LocalMux I__14774 (
            .O(N__60416),
            .I(N__60282));
    LocalMux I__14773 (
            .O(N__60413),
            .I(N__60273));
    Span4Mux_h I__14772 (
            .O(N__60410),
            .I(N__60273));
    Span4Mux_v I__14771 (
            .O(N__60407),
            .I(N__60273));
    Span4Mux_v I__14770 (
            .O(N__60398),
            .I(N__60273));
    CascadeMux I__14769 (
            .O(N__60397),
            .I(N__60270));
    InMux I__14768 (
            .O(N__60396),
            .I(N__60266));
    InMux I__14767 (
            .O(N__60395),
            .I(N__60263));
    LocalMux I__14766 (
            .O(N__60392),
            .I(N__60251));
    LocalMux I__14765 (
            .O(N__60389),
            .I(N__60251));
    LocalMux I__14764 (
            .O(N__60386),
            .I(N__60251));
    LocalMux I__14763 (
            .O(N__60381),
            .I(N__60251));
    LocalMux I__14762 (
            .O(N__60376),
            .I(N__60251));
    Span4Mux_v I__14761 (
            .O(N__60371),
            .I(N__60240));
    Span4Mux_v I__14760 (
            .O(N__60366),
            .I(N__60240));
    LocalMux I__14759 (
            .O(N__60359),
            .I(N__60240));
    InMux I__14758 (
            .O(N__60358),
            .I(N__60237));
    CascadeMux I__14757 (
            .O(N__60357),
            .I(N__60234));
    LocalMux I__14756 (
            .O(N__60354),
            .I(N__60230));
    InMux I__14755 (
            .O(N__60353),
            .I(N__60225));
    InMux I__14754 (
            .O(N__60352),
            .I(N__60225));
    LocalMux I__14753 (
            .O(N__60349),
            .I(N__60212));
    LocalMux I__14752 (
            .O(N__60344),
            .I(N__60212));
    Span4Mux_h I__14751 (
            .O(N__60341),
            .I(N__60212));
    Span4Mux_h I__14750 (
            .O(N__60336),
            .I(N__60212));
    LocalMux I__14749 (
            .O(N__60331),
            .I(N__60212));
    Span4Mux_h I__14748 (
            .O(N__60326),
            .I(N__60212));
    LocalMux I__14747 (
            .O(N__60321),
            .I(N__60209));
    LocalMux I__14746 (
            .O(N__60318),
            .I(N__60204));
    Span4Mux_v I__14745 (
            .O(N__60315),
            .I(N__60204));
    InMux I__14744 (
            .O(N__60314),
            .I(N__60195));
    InMux I__14743 (
            .O(N__60313),
            .I(N__60195));
    InMux I__14742 (
            .O(N__60310),
            .I(N__60195));
    InMux I__14741 (
            .O(N__60309),
            .I(N__60195));
    LocalMux I__14740 (
            .O(N__60304),
            .I(N__60186));
    Sp12to4 I__14739 (
            .O(N__60301),
            .I(N__60186));
    Sp12to4 I__14738 (
            .O(N__60294),
            .I(N__60186));
    Sp12to4 I__14737 (
            .O(N__60285),
            .I(N__60186));
    Span4Mux_v I__14736 (
            .O(N__60282),
            .I(N__60181));
    Span4Mux_h I__14735 (
            .O(N__60273),
            .I(N__60181));
    InMux I__14734 (
            .O(N__60270),
            .I(N__60176));
    InMux I__14733 (
            .O(N__60269),
            .I(N__60176));
    LocalMux I__14732 (
            .O(N__60266),
            .I(N__60173));
    LocalMux I__14731 (
            .O(N__60263),
            .I(N__60170));
    InMux I__14730 (
            .O(N__60262),
            .I(N__60167));
    Span4Mux_v I__14729 (
            .O(N__60251),
            .I(N__60164));
    InMux I__14728 (
            .O(N__60250),
            .I(N__60157));
    InMux I__14727 (
            .O(N__60249),
            .I(N__60157));
    InMux I__14726 (
            .O(N__60248),
            .I(N__60157));
    InMux I__14725 (
            .O(N__60247),
            .I(N__60154));
    Span4Mux_h I__14724 (
            .O(N__60240),
            .I(N__60151));
    LocalMux I__14723 (
            .O(N__60237),
            .I(N__60148));
    InMux I__14722 (
            .O(N__60234),
            .I(N__60143));
    InMux I__14721 (
            .O(N__60233),
            .I(N__60143));
    Span4Mux_v I__14720 (
            .O(N__60230),
            .I(N__60132));
    LocalMux I__14719 (
            .O(N__60225),
            .I(N__60132));
    Span4Mux_v I__14718 (
            .O(N__60212),
            .I(N__60132));
    Span4Mux_h I__14717 (
            .O(N__60209),
            .I(N__60132));
    Span4Mux_h I__14716 (
            .O(N__60204),
            .I(N__60132));
    LocalMux I__14715 (
            .O(N__60195),
            .I(N__60123));
    Span12Mux_v I__14714 (
            .O(N__60186),
            .I(N__60123));
    Sp12to4 I__14713 (
            .O(N__60181),
            .I(N__60123));
    LocalMux I__14712 (
            .O(N__60176),
            .I(N__60123));
    Odrv4 I__14711 (
            .O(N__60173),
            .I(comm_cmd_1));
    Odrv12 I__14710 (
            .O(N__60170),
            .I(comm_cmd_1));
    LocalMux I__14709 (
            .O(N__60167),
            .I(comm_cmd_1));
    Odrv4 I__14708 (
            .O(N__60164),
            .I(comm_cmd_1));
    LocalMux I__14707 (
            .O(N__60157),
            .I(comm_cmd_1));
    LocalMux I__14706 (
            .O(N__60154),
            .I(comm_cmd_1));
    Odrv4 I__14705 (
            .O(N__60151),
            .I(comm_cmd_1));
    Odrv12 I__14704 (
            .O(N__60148),
            .I(comm_cmd_1));
    LocalMux I__14703 (
            .O(N__60143),
            .I(comm_cmd_1));
    Odrv4 I__14702 (
            .O(N__60132),
            .I(comm_cmd_1));
    Odrv12 I__14701 (
            .O(N__60123),
            .I(comm_cmd_1));
    InMux I__14700 (
            .O(N__60100),
            .I(N__60087));
    InMux I__14699 (
            .O(N__60099),
            .I(N__60084));
    InMux I__14698 (
            .O(N__60098),
            .I(N__60077));
    CascadeMux I__14697 (
            .O(N__60097),
            .I(N__60073));
    InMux I__14696 (
            .O(N__60096),
            .I(N__60069));
    InMux I__14695 (
            .O(N__60095),
            .I(N__60066));
    InMux I__14694 (
            .O(N__60094),
            .I(N__60060));
    InMux I__14693 (
            .O(N__60093),
            .I(N__60053));
    InMux I__14692 (
            .O(N__60092),
            .I(N__60053));
    CascadeMux I__14691 (
            .O(N__60091),
            .I(N__60049));
    CascadeMux I__14690 (
            .O(N__60090),
            .I(N__60037));
    LocalMux I__14689 (
            .O(N__60087),
            .I(N__60031));
    LocalMux I__14688 (
            .O(N__60084),
            .I(N__60031));
    InMux I__14687 (
            .O(N__60083),
            .I(N__60026));
    InMux I__14686 (
            .O(N__60082),
            .I(N__60026));
    InMux I__14685 (
            .O(N__60081),
            .I(N__60021));
    InMux I__14684 (
            .O(N__60080),
            .I(N__60021));
    LocalMux I__14683 (
            .O(N__60077),
            .I(N__60018));
    InMux I__14682 (
            .O(N__60076),
            .I(N__60015));
    InMux I__14681 (
            .O(N__60073),
            .I(N__60009));
    InMux I__14680 (
            .O(N__60072),
            .I(N__60009));
    LocalMux I__14679 (
            .O(N__60069),
            .I(N__60003));
    LocalMux I__14678 (
            .O(N__60066),
            .I(N__59996));
    InMux I__14677 (
            .O(N__60065),
            .I(N__59988));
    InMux I__14676 (
            .O(N__60064),
            .I(N__59979));
    InMux I__14675 (
            .O(N__60063),
            .I(N__59970));
    LocalMux I__14674 (
            .O(N__60060),
            .I(N__59966));
    InMux I__14673 (
            .O(N__60059),
            .I(N__59955));
    InMux I__14672 (
            .O(N__60058),
            .I(N__59955));
    LocalMux I__14671 (
            .O(N__60053),
            .I(N__59951));
    InMux I__14670 (
            .O(N__60052),
            .I(N__59944));
    InMux I__14669 (
            .O(N__60049),
            .I(N__59944));
    InMux I__14668 (
            .O(N__60048),
            .I(N__59944));
    InMux I__14667 (
            .O(N__60047),
            .I(N__59937));
    InMux I__14666 (
            .O(N__60046),
            .I(N__59937));
    InMux I__14665 (
            .O(N__60045),
            .I(N__59937));
    CascadeMux I__14664 (
            .O(N__60044),
            .I(N__59933));
    CascadeMux I__14663 (
            .O(N__60043),
            .I(N__59930));
    InMux I__14662 (
            .O(N__60042),
            .I(N__59925));
    InMux I__14661 (
            .O(N__60041),
            .I(N__59925));
    InMux I__14660 (
            .O(N__60040),
            .I(N__59922));
    InMux I__14659 (
            .O(N__60037),
            .I(N__59917));
    InMux I__14658 (
            .O(N__60036),
            .I(N__59917));
    Span4Mux_v I__14657 (
            .O(N__60031),
            .I(N__59912));
    LocalMux I__14656 (
            .O(N__60026),
            .I(N__59912));
    LocalMux I__14655 (
            .O(N__60021),
            .I(N__59905));
    Span4Mux_v I__14654 (
            .O(N__60018),
            .I(N__59905));
    LocalMux I__14653 (
            .O(N__60015),
            .I(N__59905));
    CascadeMux I__14652 (
            .O(N__60014),
            .I(N__59901));
    LocalMux I__14651 (
            .O(N__60009),
            .I(N__59897));
    InMux I__14650 (
            .O(N__60008),
            .I(N__59894));
    InMux I__14649 (
            .O(N__60007),
            .I(N__59891));
    InMux I__14648 (
            .O(N__60006),
            .I(N__59888));
    Span4Mux_v I__14647 (
            .O(N__60003),
            .I(N__59884));
    InMux I__14646 (
            .O(N__60002),
            .I(N__59881));
    InMux I__14645 (
            .O(N__60001),
            .I(N__59874));
    InMux I__14644 (
            .O(N__60000),
            .I(N__59874));
    InMux I__14643 (
            .O(N__59999),
            .I(N__59874));
    Span4Mux_v I__14642 (
            .O(N__59996),
            .I(N__59871));
    InMux I__14641 (
            .O(N__59995),
            .I(N__59868));
    InMux I__14640 (
            .O(N__59994),
            .I(N__59862));
    InMux I__14639 (
            .O(N__59993),
            .I(N__59862));
    InMux I__14638 (
            .O(N__59992),
            .I(N__59857));
    InMux I__14637 (
            .O(N__59991),
            .I(N__59857));
    LocalMux I__14636 (
            .O(N__59988),
            .I(N__59854));
    InMux I__14635 (
            .O(N__59987),
            .I(N__59851));
    InMux I__14634 (
            .O(N__59986),
            .I(N__59846));
    InMux I__14633 (
            .O(N__59985),
            .I(N__59846));
    InMux I__14632 (
            .O(N__59984),
            .I(N__59839));
    InMux I__14631 (
            .O(N__59983),
            .I(N__59839));
    InMux I__14630 (
            .O(N__59982),
            .I(N__59839));
    LocalMux I__14629 (
            .O(N__59979),
            .I(N__59836));
    InMux I__14628 (
            .O(N__59978),
            .I(N__59831));
    InMux I__14627 (
            .O(N__59977),
            .I(N__59831));
    InMux I__14626 (
            .O(N__59976),
            .I(N__59828));
    InMux I__14625 (
            .O(N__59975),
            .I(N__59823));
    InMux I__14624 (
            .O(N__59974),
            .I(N__59823));
    CascadeMux I__14623 (
            .O(N__59973),
            .I(N__59819));
    LocalMux I__14622 (
            .O(N__59970),
            .I(N__59816));
    InMux I__14621 (
            .O(N__59969),
            .I(N__59813));
    Span4Mux_h I__14620 (
            .O(N__59966),
            .I(N__59809));
    InMux I__14619 (
            .O(N__59965),
            .I(N__59802));
    InMux I__14618 (
            .O(N__59964),
            .I(N__59802));
    InMux I__14617 (
            .O(N__59963),
            .I(N__59802));
    InMux I__14616 (
            .O(N__59962),
            .I(N__59797));
    InMux I__14615 (
            .O(N__59961),
            .I(N__59797));
    InMux I__14614 (
            .O(N__59960),
            .I(N__59794));
    LocalMux I__14613 (
            .O(N__59955),
            .I(N__59791));
    InMux I__14612 (
            .O(N__59954),
            .I(N__59788));
    Span4Mux_v I__14611 (
            .O(N__59951),
            .I(N__59785));
    LocalMux I__14610 (
            .O(N__59944),
            .I(N__59780));
    LocalMux I__14609 (
            .O(N__59937),
            .I(N__59780));
    InMux I__14608 (
            .O(N__59936),
            .I(N__59777));
    InMux I__14607 (
            .O(N__59933),
            .I(N__59772));
    InMux I__14606 (
            .O(N__59930),
            .I(N__59772));
    LocalMux I__14605 (
            .O(N__59925),
            .I(N__59769));
    LocalMux I__14604 (
            .O(N__59922),
            .I(N__59764));
    LocalMux I__14603 (
            .O(N__59917),
            .I(N__59764));
    Span4Mux_h I__14602 (
            .O(N__59912),
            .I(N__59759));
    Span4Mux_v I__14601 (
            .O(N__59905),
            .I(N__59759));
    InMux I__14600 (
            .O(N__59904),
            .I(N__59756));
    InMux I__14599 (
            .O(N__59901),
            .I(N__59751));
    InMux I__14598 (
            .O(N__59900),
            .I(N__59751));
    Span4Mux_h I__14597 (
            .O(N__59897),
            .I(N__59748));
    LocalMux I__14596 (
            .O(N__59894),
            .I(N__59743));
    LocalMux I__14595 (
            .O(N__59891),
            .I(N__59743));
    LocalMux I__14594 (
            .O(N__59888),
            .I(N__59740));
    InMux I__14593 (
            .O(N__59887),
            .I(N__59737));
    Span4Mux_h I__14592 (
            .O(N__59884),
            .I(N__59734));
    LocalMux I__14591 (
            .O(N__59881),
            .I(N__59725));
    LocalMux I__14590 (
            .O(N__59874),
            .I(N__59725));
    Span4Mux_h I__14589 (
            .O(N__59871),
            .I(N__59725));
    LocalMux I__14588 (
            .O(N__59868),
            .I(N__59725));
    InMux I__14587 (
            .O(N__59867),
            .I(N__59722));
    LocalMux I__14586 (
            .O(N__59862),
            .I(N__59717));
    LocalMux I__14585 (
            .O(N__59857),
            .I(N__59717));
    Span4Mux_v I__14584 (
            .O(N__59854),
            .I(N__59704));
    LocalMux I__14583 (
            .O(N__59851),
            .I(N__59704));
    LocalMux I__14582 (
            .O(N__59846),
            .I(N__59704));
    LocalMux I__14581 (
            .O(N__59839),
            .I(N__59704));
    Span4Mux_h I__14580 (
            .O(N__59836),
            .I(N__59704));
    LocalMux I__14579 (
            .O(N__59831),
            .I(N__59704));
    LocalMux I__14578 (
            .O(N__59828),
            .I(N__59697));
    LocalMux I__14577 (
            .O(N__59823),
            .I(N__59697));
    InMux I__14576 (
            .O(N__59822),
            .I(N__59692));
    InMux I__14575 (
            .O(N__59819),
            .I(N__59692));
    Span4Mux_h I__14574 (
            .O(N__59816),
            .I(N__59687));
    LocalMux I__14573 (
            .O(N__59813),
            .I(N__59687));
    InMux I__14572 (
            .O(N__59812),
            .I(N__59684));
    Span4Mux_h I__14571 (
            .O(N__59809),
            .I(N__59673));
    LocalMux I__14570 (
            .O(N__59802),
            .I(N__59673));
    LocalMux I__14569 (
            .O(N__59797),
            .I(N__59673));
    LocalMux I__14568 (
            .O(N__59794),
            .I(N__59673));
    Span4Mux_h I__14567 (
            .O(N__59791),
            .I(N__59673));
    LocalMux I__14566 (
            .O(N__59788),
            .I(N__59661));
    Sp12to4 I__14565 (
            .O(N__59785),
            .I(N__59661));
    Span12Mux_h I__14564 (
            .O(N__59780),
            .I(N__59661));
    LocalMux I__14563 (
            .O(N__59777),
            .I(N__59661));
    LocalMux I__14562 (
            .O(N__59772),
            .I(N__59661));
    Span4Mux_v I__14561 (
            .O(N__59769),
            .I(N__59654));
    Span4Mux_v I__14560 (
            .O(N__59764),
            .I(N__59654));
    Span4Mux_h I__14559 (
            .O(N__59759),
            .I(N__59654));
    LocalMux I__14558 (
            .O(N__59756),
            .I(N__59649));
    LocalMux I__14557 (
            .O(N__59751),
            .I(N__59649));
    Span4Mux_v I__14556 (
            .O(N__59748),
            .I(N__59644));
    Span4Mux_h I__14555 (
            .O(N__59743),
            .I(N__59644));
    Span4Mux_v I__14554 (
            .O(N__59740),
            .I(N__59629));
    LocalMux I__14553 (
            .O(N__59737),
            .I(N__59629));
    Span4Mux_h I__14552 (
            .O(N__59734),
            .I(N__59629));
    Span4Mux_v I__14551 (
            .O(N__59725),
            .I(N__59629));
    LocalMux I__14550 (
            .O(N__59722),
            .I(N__59629));
    Span4Mux_v I__14549 (
            .O(N__59717),
            .I(N__59629));
    Span4Mux_v I__14548 (
            .O(N__59704),
            .I(N__59629));
    InMux I__14547 (
            .O(N__59703),
            .I(N__59624));
    InMux I__14546 (
            .O(N__59702),
            .I(N__59624));
    Span4Mux_v I__14545 (
            .O(N__59697),
            .I(N__59619));
    LocalMux I__14544 (
            .O(N__59692),
            .I(N__59619));
    Span4Mux_v I__14543 (
            .O(N__59687),
            .I(N__59612));
    LocalMux I__14542 (
            .O(N__59684),
            .I(N__59612));
    Span4Mux_v I__14541 (
            .O(N__59673),
            .I(N__59612));
    InMux I__14540 (
            .O(N__59672),
            .I(N__59609));
    Span12Mux_h I__14539 (
            .O(N__59661),
            .I(N__59606));
    Span4Mux_h I__14538 (
            .O(N__59654),
            .I(N__59601));
    Span4Mux_v I__14537 (
            .O(N__59649),
            .I(N__59601));
    Odrv4 I__14536 (
            .O(N__59644),
            .I(comm_cmd_2));
    Odrv4 I__14535 (
            .O(N__59629),
            .I(comm_cmd_2));
    LocalMux I__14534 (
            .O(N__59624),
            .I(comm_cmd_2));
    Odrv4 I__14533 (
            .O(N__59619),
            .I(comm_cmd_2));
    Odrv4 I__14532 (
            .O(N__59612),
            .I(comm_cmd_2));
    LocalMux I__14531 (
            .O(N__59609),
            .I(comm_cmd_2));
    Odrv12 I__14530 (
            .O(N__59606),
            .I(comm_cmd_2));
    Odrv4 I__14529 (
            .O(N__59601),
            .I(comm_cmd_2));
    CascadeMux I__14528 (
            .O(N__59584),
            .I(N__59581));
    InMux I__14527 (
            .O(N__59581),
            .I(N__59578));
    LocalMux I__14526 (
            .O(N__59578),
            .I(N__59575));
    Odrv4 I__14525 (
            .O(N__59575),
            .I(n22316));
    InMux I__14524 (
            .O(N__59572),
            .I(N__59569));
    LocalMux I__14523 (
            .O(N__59569),
            .I(n26_adj_1792));
    InMux I__14522 (
            .O(N__59566),
            .I(N__59563));
    LocalMux I__14521 (
            .O(N__59563),
            .I(n23456));
    InMux I__14520 (
            .O(N__59560),
            .I(N__59557));
    LocalMux I__14519 (
            .O(N__59557),
            .I(buf_data_iac_13));
    InMux I__14518 (
            .O(N__59554),
            .I(N__59551));
    LocalMux I__14517 (
            .O(N__59551),
            .I(N__59548));
    Span4Mux_h I__14516 (
            .O(N__59548),
            .I(N__59545));
    Odrv4 I__14515 (
            .O(N__59545),
            .I(n22313));
    InMux I__14514 (
            .O(N__59542),
            .I(N__59539));
    LocalMux I__14513 (
            .O(N__59539),
            .I(buf_data_iac_11));
    InMux I__14512 (
            .O(N__59536),
            .I(N__59533));
    LocalMux I__14511 (
            .O(N__59533),
            .I(N__59530));
    Odrv12 I__14510 (
            .O(N__59530),
            .I(n22300));
    InMux I__14509 (
            .O(N__59527),
            .I(N__59524));
    LocalMux I__14508 (
            .O(N__59524),
            .I(N__59521));
    Odrv4 I__14507 (
            .O(N__59521),
            .I(buf_data_iac_8));
    CascadeMux I__14506 (
            .O(N__59518),
            .I(N__59510));
    CascadeMux I__14505 (
            .O(N__59517),
            .I(N__59498));
    InMux I__14504 (
            .O(N__59516),
            .I(N__59493));
    InMux I__14503 (
            .O(N__59515),
            .I(N__59485));
    CascadeMux I__14502 (
            .O(N__59514),
            .I(N__59480));
    CascadeMux I__14501 (
            .O(N__59513),
            .I(N__59476));
    InMux I__14500 (
            .O(N__59510),
            .I(N__59472));
    InMux I__14499 (
            .O(N__59509),
            .I(N__59469));
    InMux I__14498 (
            .O(N__59508),
            .I(N__59461));
    InMux I__14497 (
            .O(N__59507),
            .I(N__59461));
    InMux I__14496 (
            .O(N__59506),
            .I(N__59458));
    InMux I__14495 (
            .O(N__59505),
            .I(N__59455));
    InMux I__14494 (
            .O(N__59504),
            .I(N__59450));
    InMux I__14493 (
            .O(N__59503),
            .I(N__59450));
    InMux I__14492 (
            .O(N__59502),
            .I(N__59447));
    InMux I__14491 (
            .O(N__59501),
            .I(N__59417));
    InMux I__14490 (
            .O(N__59498),
            .I(N__59414));
    InMux I__14489 (
            .O(N__59497),
            .I(N__59411));
    InMux I__14488 (
            .O(N__59496),
            .I(N__59402));
    LocalMux I__14487 (
            .O(N__59493),
            .I(N__59394));
    InMux I__14486 (
            .O(N__59492),
            .I(N__59391));
    InMux I__14485 (
            .O(N__59491),
            .I(N__59388));
    InMux I__14484 (
            .O(N__59490),
            .I(N__59381));
    InMux I__14483 (
            .O(N__59489),
            .I(N__59381));
    InMux I__14482 (
            .O(N__59488),
            .I(N__59381));
    LocalMux I__14481 (
            .O(N__59485),
            .I(N__59378));
    InMux I__14480 (
            .O(N__59484),
            .I(N__59373));
    InMux I__14479 (
            .O(N__59483),
            .I(N__59373));
    InMux I__14478 (
            .O(N__59480),
            .I(N__59368));
    InMux I__14477 (
            .O(N__59479),
            .I(N__59359));
    InMux I__14476 (
            .O(N__59476),
            .I(N__59356));
    InMux I__14475 (
            .O(N__59475),
            .I(N__59347));
    LocalMux I__14474 (
            .O(N__59472),
            .I(N__59342));
    LocalMux I__14473 (
            .O(N__59469),
            .I(N__59342));
    InMux I__14472 (
            .O(N__59468),
            .I(N__59337));
    InMux I__14471 (
            .O(N__59467),
            .I(N__59337));
    InMux I__14470 (
            .O(N__59466),
            .I(N__59332));
    LocalMux I__14469 (
            .O(N__59461),
            .I(N__59317));
    LocalMux I__14468 (
            .O(N__59458),
            .I(N__59308));
    LocalMux I__14467 (
            .O(N__59455),
            .I(N__59308));
    LocalMux I__14466 (
            .O(N__59450),
            .I(N__59308));
    LocalMux I__14465 (
            .O(N__59447),
            .I(N__59308));
    InMux I__14464 (
            .O(N__59446),
            .I(N__59298));
    InMux I__14463 (
            .O(N__59445),
            .I(N__59298));
    InMux I__14462 (
            .O(N__59444),
            .I(N__59298));
    InMux I__14461 (
            .O(N__59443),
            .I(N__59293));
    InMux I__14460 (
            .O(N__59442),
            .I(N__59293));
    InMux I__14459 (
            .O(N__59441),
            .I(N__59288));
    InMux I__14458 (
            .O(N__59440),
            .I(N__59288));
    InMux I__14457 (
            .O(N__59439),
            .I(N__59283));
    InMux I__14456 (
            .O(N__59438),
            .I(N__59283));
    InMux I__14455 (
            .O(N__59437),
            .I(N__59278));
    InMux I__14454 (
            .O(N__59436),
            .I(N__59278));
    InMux I__14453 (
            .O(N__59435),
            .I(N__59269));
    InMux I__14452 (
            .O(N__59434),
            .I(N__59269));
    InMux I__14451 (
            .O(N__59433),
            .I(N__59269));
    InMux I__14450 (
            .O(N__59432),
            .I(N__59269));
    InMux I__14449 (
            .O(N__59431),
            .I(N__59258));
    InMux I__14448 (
            .O(N__59430),
            .I(N__59251));
    InMux I__14447 (
            .O(N__59429),
            .I(N__59251));
    InMux I__14446 (
            .O(N__59428),
            .I(N__59251));
    InMux I__14445 (
            .O(N__59427),
            .I(N__59247));
    InMux I__14444 (
            .O(N__59426),
            .I(N__59241));
    InMux I__14443 (
            .O(N__59425),
            .I(N__59241));
    InMux I__14442 (
            .O(N__59424),
            .I(N__59238));
    InMux I__14441 (
            .O(N__59423),
            .I(N__59231));
    InMux I__14440 (
            .O(N__59422),
            .I(N__59231));
    InMux I__14439 (
            .O(N__59421),
            .I(N__59231));
    InMux I__14438 (
            .O(N__59420),
            .I(N__59228));
    LocalMux I__14437 (
            .O(N__59417),
            .I(N__59218));
    LocalMux I__14436 (
            .O(N__59414),
            .I(N__59218));
    LocalMux I__14435 (
            .O(N__59411),
            .I(N__59218));
    InMux I__14434 (
            .O(N__59410),
            .I(N__59215));
    InMux I__14433 (
            .O(N__59409),
            .I(N__59210));
    InMux I__14432 (
            .O(N__59408),
            .I(N__59210));
    InMux I__14431 (
            .O(N__59407),
            .I(N__59206));
    InMux I__14430 (
            .O(N__59406),
            .I(N__59201));
    InMux I__14429 (
            .O(N__59405),
            .I(N__59201));
    LocalMux I__14428 (
            .O(N__59402),
            .I(N__59198));
    InMux I__14427 (
            .O(N__59401),
            .I(N__59193));
    InMux I__14426 (
            .O(N__59400),
            .I(N__59193));
    InMux I__14425 (
            .O(N__59399),
            .I(N__59186));
    InMux I__14424 (
            .O(N__59398),
            .I(N__59182));
    InMux I__14423 (
            .O(N__59397),
            .I(N__59178));
    Span4Mux_v I__14422 (
            .O(N__59394),
            .I(N__59165));
    LocalMux I__14421 (
            .O(N__59391),
            .I(N__59165));
    LocalMux I__14420 (
            .O(N__59388),
            .I(N__59165));
    LocalMux I__14419 (
            .O(N__59381),
            .I(N__59165));
    Span4Mux_h I__14418 (
            .O(N__59378),
            .I(N__59165));
    LocalMux I__14417 (
            .O(N__59373),
            .I(N__59165));
    InMux I__14416 (
            .O(N__59372),
            .I(N__59160));
    InMux I__14415 (
            .O(N__59371),
            .I(N__59160));
    LocalMux I__14414 (
            .O(N__59368),
            .I(N__59157));
    InMux I__14413 (
            .O(N__59367),
            .I(N__59148));
    InMux I__14412 (
            .O(N__59366),
            .I(N__59148));
    InMux I__14411 (
            .O(N__59365),
            .I(N__59148));
    InMux I__14410 (
            .O(N__59364),
            .I(N__59148));
    InMux I__14409 (
            .O(N__59363),
            .I(N__59143));
    InMux I__14408 (
            .O(N__59362),
            .I(N__59143));
    LocalMux I__14407 (
            .O(N__59359),
            .I(N__59138));
    LocalMux I__14406 (
            .O(N__59356),
            .I(N__59138));
    InMux I__14405 (
            .O(N__59355),
            .I(N__59127));
    InMux I__14404 (
            .O(N__59354),
            .I(N__59127));
    InMux I__14403 (
            .O(N__59353),
            .I(N__59127));
    InMux I__14402 (
            .O(N__59352),
            .I(N__59127));
    InMux I__14401 (
            .O(N__59351),
            .I(N__59127));
    InMux I__14400 (
            .O(N__59350),
            .I(N__59124));
    LocalMux I__14399 (
            .O(N__59347),
            .I(N__59121));
    Span4Mux_v I__14398 (
            .O(N__59342),
            .I(N__59116));
    LocalMux I__14397 (
            .O(N__59337),
            .I(N__59116));
    InMux I__14396 (
            .O(N__59336),
            .I(N__59106));
    InMux I__14395 (
            .O(N__59335),
            .I(N__59106));
    LocalMux I__14394 (
            .O(N__59332),
            .I(N__59103));
    InMux I__14393 (
            .O(N__59331),
            .I(N__59094));
    InMux I__14392 (
            .O(N__59330),
            .I(N__59094));
    InMux I__14391 (
            .O(N__59329),
            .I(N__59094));
    InMux I__14390 (
            .O(N__59328),
            .I(N__59094));
    InMux I__14389 (
            .O(N__59327),
            .I(N__59091));
    InMux I__14388 (
            .O(N__59326),
            .I(N__59082));
    InMux I__14387 (
            .O(N__59325),
            .I(N__59082));
    InMux I__14386 (
            .O(N__59324),
            .I(N__59082));
    InMux I__14385 (
            .O(N__59323),
            .I(N__59082));
    InMux I__14384 (
            .O(N__59322),
            .I(N__59079));
    InMux I__14383 (
            .O(N__59321),
            .I(N__59074));
    InMux I__14382 (
            .O(N__59320),
            .I(N__59074));
    Span4Mux_v I__14381 (
            .O(N__59317),
            .I(N__59069));
    Span4Mux_v I__14380 (
            .O(N__59308),
            .I(N__59069));
    InMux I__14379 (
            .O(N__59307),
            .I(N__59066));
    InMux I__14378 (
            .O(N__59306),
            .I(N__59063));
    InMux I__14377 (
            .O(N__59305),
            .I(N__59060));
    LocalMux I__14376 (
            .O(N__59298),
            .I(N__59057));
    LocalMux I__14375 (
            .O(N__59293),
            .I(N__59050));
    LocalMux I__14374 (
            .O(N__59288),
            .I(N__59050));
    LocalMux I__14373 (
            .O(N__59283),
            .I(N__59050));
    LocalMux I__14372 (
            .O(N__59278),
            .I(N__59045));
    LocalMux I__14371 (
            .O(N__59269),
            .I(N__59045));
    InMux I__14370 (
            .O(N__59268),
            .I(N__59042));
    InMux I__14369 (
            .O(N__59267),
            .I(N__59035));
    InMux I__14368 (
            .O(N__59266),
            .I(N__59035));
    InMux I__14367 (
            .O(N__59265),
            .I(N__59035));
    InMux I__14366 (
            .O(N__59264),
            .I(N__59026));
    InMux I__14365 (
            .O(N__59263),
            .I(N__59026));
    InMux I__14364 (
            .O(N__59262),
            .I(N__59026));
    InMux I__14363 (
            .O(N__59261),
            .I(N__59026));
    LocalMux I__14362 (
            .O(N__59258),
            .I(N__59021));
    LocalMux I__14361 (
            .O(N__59251),
            .I(N__59021));
    InMux I__14360 (
            .O(N__59250),
            .I(N__59017));
    LocalMux I__14359 (
            .O(N__59247),
            .I(N__59011));
    InMux I__14358 (
            .O(N__59246),
            .I(N__59006));
    LocalMux I__14357 (
            .O(N__59241),
            .I(N__58999));
    LocalMux I__14356 (
            .O(N__59238),
            .I(N__58999));
    LocalMux I__14355 (
            .O(N__59231),
            .I(N__58999));
    LocalMux I__14354 (
            .O(N__59228),
            .I(N__58996));
    InMux I__14353 (
            .O(N__59227),
            .I(N__58993));
    InMux I__14352 (
            .O(N__59226),
            .I(N__58988));
    InMux I__14351 (
            .O(N__59225),
            .I(N__58988));
    Span4Mux_v I__14350 (
            .O(N__59218),
            .I(N__58981));
    LocalMux I__14349 (
            .O(N__59215),
            .I(N__58981));
    LocalMux I__14348 (
            .O(N__59210),
            .I(N__58981));
    InMux I__14347 (
            .O(N__59209),
            .I(N__58978));
    LocalMux I__14346 (
            .O(N__59206),
            .I(N__58973));
    LocalMux I__14345 (
            .O(N__59201),
            .I(N__58973));
    Span4Mux_v I__14344 (
            .O(N__59198),
            .I(N__58968));
    LocalMux I__14343 (
            .O(N__59193),
            .I(N__58968));
    InMux I__14342 (
            .O(N__59192),
            .I(N__58963));
    InMux I__14341 (
            .O(N__59191),
            .I(N__58963));
    InMux I__14340 (
            .O(N__59190),
            .I(N__58960));
    InMux I__14339 (
            .O(N__59189),
            .I(N__58957));
    LocalMux I__14338 (
            .O(N__59186),
            .I(N__58954));
    InMux I__14337 (
            .O(N__59185),
            .I(N__58951));
    LocalMux I__14336 (
            .O(N__59182),
            .I(N__58945));
    InMux I__14335 (
            .O(N__59181),
            .I(N__58942));
    LocalMux I__14334 (
            .O(N__59178),
            .I(N__58939));
    Span4Mux_v I__14333 (
            .O(N__59165),
            .I(N__58934));
    LocalMux I__14332 (
            .O(N__59160),
            .I(N__58934));
    Span4Mux_v I__14331 (
            .O(N__59157),
            .I(N__58923));
    LocalMux I__14330 (
            .O(N__59148),
            .I(N__58923));
    LocalMux I__14329 (
            .O(N__59143),
            .I(N__58923));
    Span4Mux_v I__14328 (
            .O(N__59138),
            .I(N__58923));
    LocalMux I__14327 (
            .O(N__59127),
            .I(N__58923));
    LocalMux I__14326 (
            .O(N__59124),
            .I(N__58916));
    Span4Mux_h I__14325 (
            .O(N__59121),
            .I(N__58916));
    Span4Mux_h I__14324 (
            .O(N__59116),
            .I(N__58916));
    InMux I__14323 (
            .O(N__59115),
            .I(N__58908));
    InMux I__14322 (
            .O(N__59114),
            .I(N__58908));
    InMux I__14321 (
            .O(N__59113),
            .I(N__58908));
    InMux I__14320 (
            .O(N__59112),
            .I(N__58905));
    InMux I__14319 (
            .O(N__59111),
            .I(N__58902));
    LocalMux I__14318 (
            .O(N__59106),
            .I(N__58899));
    Span4Mux_v I__14317 (
            .O(N__59103),
            .I(N__58896));
    LocalMux I__14316 (
            .O(N__59094),
            .I(N__58889));
    LocalMux I__14315 (
            .O(N__59091),
            .I(N__58889));
    LocalMux I__14314 (
            .O(N__59082),
            .I(N__58889));
    LocalMux I__14313 (
            .O(N__59079),
            .I(N__58870));
    LocalMux I__14312 (
            .O(N__59074),
            .I(N__58870));
    Span4Mux_h I__14311 (
            .O(N__59069),
            .I(N__58870));
    LocalMux I__14310 (
            .O(N__59066),
            .I(N__58870));
    LocalMux I__14309 (
            .O(N__59063),
            .I(N__58870));
    LocalMux I__14308 (
            .O(N__59060),
            .I(N__58870));
    Span4Mux_h I__14307 (
            .O(N__59057),
            .I(N__58870));
    Span4Mux_v I__14306 (
            .O(N__59050),
            .I(N__58870));
    Span4Mux_v I__14305 (
            .O(N__59045),
            .I(N__58870));
    LocalMux I__14304 (
            .O(N__59042),
            .I(N__58861));
    LocalMux I__14303 (
            .O(N__59035),
            .I(N__58861));
    LocalMux I__14302 (
            .O(N__59026),
            .I(N__58861));
    Span4Mux_v I__14301 (
            .O(N__59021),
            .I(N__58861));
    InMux I__14300 (
            .O(N__59020),
            .I(N__58858));
    LocalMux I__14299 (
            .O(N__59017),
            .I(N__58852));
    InMux I__14298 (
            .O(N__59016),
            .I(N__58845));
    InMux I__14297 (
            .O(N__59015),
            .I(N__58845));
    InMux I__14296 (
            .O(N__59014),
            .I(N__58845));
    Span4Mux_h I__14295 (
            .O(N__59011),
            .I(N__58837));
    InMux I__14294 (
            .O(N__59010),
            .I(N__58831));
    InMux I__14293 (
            .O(N__59009),
            .I(N__58831));
    LocalMux I__14292 (
            .O(N__59006),
            .I(N__58828));
    Span4Mux_v I__14291 (
            .O(N__58999),
            .I(N__58823));
    Span4Mux_v I__14290 (
            .O(N__58996),
            .I(N__58823));
    LocalMux I__14289 (
            .O(N__58993),
            .I(N__58814));
    LocalMux I__14288 (
            .O(N__58988),
            .I(N__58814));
    Span4Mux_h I__14287 (
            .O(N__58981),
            .I(N__58814));
    LocalMux I__14286 (
            .O(N__58978),
            .I(N__58814));
    Span4Mux_v I__14285 (
            .O(N__58973),
            .I(N__58807));
    Span4Mux_v I__14284 (
            .O(N__58968),
            .I(N__58807));
    LocalMux I__14283 (
            .O(N__58963),
            .I(N__58807));
    LocalMux I__14282 (
            .O(N__58960),
            .I(N__58798));
    LocalMux I__14281 (
            .O(N__58957),
            .I(N__58798));
    Span4Mux_h I__14280 (
            .O(N__58954),
            .I(N__58798));
    LocalMux I__14279 (
            .O(N__58951),
            .I(N__58798));
    InMux I__14278 (
            .O(N__58950),
            .I(N__58791));
    InMux I__14277 (
            .O(N__58949),
            .I(N__58791));
    InMux I__14276 (
            .O(N__58948),
            .I(N__58791));
    Span4Mux_h I__14275 (
            .O(N__58945),
            .I(N__58784));
    LocalMux I__14274 (
            .O(N__58942),
            .I(N__58784));
    Span4Mux_v I__14273 (
            .O(N__58939),
            .I(N__58784));
    Span4Mux_h I__14272 (
            .O(N__58934),
            .I(N__58777));
    Span4Mux_v I__14271 (
            .O(N__58923),
            .I(N__58777));
    Span4Mux_h I__14270 (
            .O(N__58916),
            .I(N__58777));
    InMux I__14269 (
            .O(N__58915),
            .I(N__58774));
    LocalMux I__14268 (
            .O(N__58908),
            .I(N__58771));
    LocalMux I__14267 (
            .O(N__58905),
            .I(N__58766));
    LocalMux I__14266 (
            .O(N__58902),
            .I(N__58766));
    Span4Mux_h I__14265 (
            .O(N__58899),
            .I(N__58753));
    Span4Mux_h I__14264 (
            .O(N__58896),
            .I(N__58753));
    Span4Mux_v I__14263 (
            .O(N__58889),
            .I(N__58753));
    Span4Mux_v I__14262 (
            .O(N__58870),
            .I(N__58753));
    Span4Mux_v I__14261 (
            .O(N__58861),
            .I(N__58753));
    LocalMux I__14260 (
            .O(N__58858),
            .I(N__58753));
    InMux I__14259 (
            .O(N__58857),
            .I(N__58746));
    InMux I__14258 (
            .O(N__58856),
            .I(N__58746));
    InMux I__14257 (
            .O(N__58855),
            .I(N__58746));
    Span4Mux_h I__14256 (
            .O(N__58852),
            .I(N__58743));
    LocalMux I__14255 (
            .O(N__58845),
            .I(N__58740));
    InMux I__14254 (
            .O(N__58844),
            .I(N__58733));
    InMux I__14253 (
            .O(N__58843),
            .I(N__58733));
    InMux I__14252 (
            .O(N__58842),
            .I(N__58733));
    InMux I__14251 (
            .O(N__58841),
            .I(N__58730));
    InMux I__14250 (
            .O(N__58840),
            .I(N__58727));
    Span4Mux_v I__14249 (
            .O(N__58837),
            .I(N__58724));
    InMux I__14248 (
            .O(N__58836),
            .I(N__58721));
    LocalMux I__14247 (
            .O(N__58831),
            .I(N__58716));
    Span12Mux_h I__14246 (
            .O(N__58828),
            .I(N__58716));
    Span4Mux_h I__14245 (
            .O(N__58823),
            .I(N__58709));
    Span4Mux_v I__14244 (
            .O(N__58814),
            .I(N__58709));
    Span4Mux_h I__14243 (
            .O(N__58807),
            .I(N__58709));
    Span4Mux_v I__14242 (
            .O(N__58798),
            .I(N__58700));
    LocalMux I__14241 (
            .O(N__58791),
            .I(N__58700));
    Span4Mux_h I__14240 (
            .O(N__58784),
            .I(N__58700));
    Span4Mux_h I__14239 (
            .O(N__58777),
            .I(N__58700));
    LocalMux I__14238 (
            .O(N__58774),
            .I(N__58689));
    Span12Mux_v I__14237 (
            .O(N__58771),
            .I(N__58689));
    Span12Mux_h I__14236 (
            .O(N__58766),
            .I(N__58689));
    Sp12to4 I__14235 (
            .O(N__58753),
            .I(N__58689));
    LocalMux I__14234 (
            .O(N__58746),
            .I(N__58689));
    Odrv4 I__14233 (
            .O(N__58743),
            .I(comm_cmd_0));
    Odrv4 I__14232 (
            .O(N__58740),
            .I(comm_cmd_0));
    LocalMux I__14231 (
            .O(N__58733),
            .I(comm_cmd_0));
    LocalMux I__14230 (
            .O(N__58730),
            .I(comm_cmd_0));
    LocalMux I__14229 (
            .O(N__58727),
            .I(comm_cmd_0));
    Odrv4 I__14228 (
            .O(N__58724),
            .I(comm_cmd_0));
    LocalMux I__14227 (
            .O(N__58721),
            .I(comm_cmd_0));
    Odrv12 I__14226 (
            .O(N__58716),
            .I(comm_cmd_0));
    Odrv4 I__14225 (
            .O(N__58709),
            .I(comm_cmd_0));
    Odrv4 I__14224 (
            .O(N__58700),
            .I(comm_cmd_0));
    Odrv12 I__14223 (
            .O(N__58689),
            .I(comm_cmd_0));
    InMux I__14222 (
            .O(N__58666),
            .I(N__58663));
    LocalMux I__14221 (
            .O(N__58663),
            .I(N__58660));
    Span4Mux_h I__14220 (
            .O(N__58660),
            .I(N__58657));
    Odrv4 I__14219 (
            .O(N__58657),
            .I(n22649));
    InMux I__14218 (
            .O(N__58654),
            .I(N__58643));
    InMux I__14217 (
            .O(N__58653),
            .I(N__58643));
    InMux I__14216 (
            .O(N__58652),
            .I(N__58638));
    InMux I__14215 (
            .O(N__58651),
            .I(N__58635));
    InMux I__14214 (
            .O(N__58650),
            .I(N__58630));
    InMux I__14213 (
            .O(N__58649),
            .I(N__58630));
    InMux I__14212 (
            .O(N__58648),
            .I(N__58627));
    LocalMux I__14211 (
            .O(N__58643),
            .I(N__58621));
    InMux I__14210 (
            .O(N__58642),
            .I(N__58616));
    InMux I__14209 (
            .O(N__58641),
            .I(N__58616));
    LocalMux I__14208 (
            .O(N__58638),
            .I(N__58611));
    LocalMux I__14207 (
            .O(N__58635),
            .I(N__58602));
    LocalMux I__14206 (
            .O(N__58630),
            .I(N__58602));
    LocalMux I__14205 (
            .O(N__58627),
            .I(N__58599));
    InMux I__14204 (
            .O(N__58626),
            .I(N__58594));
    InMux I__14203 (
            .O(N__58625),
            .I(N__58594));
    InMux I__14202 (
            .O(N__58624),
            .I(N__58591));
    Span4Mux_v I__14201 (
            .O(N__58621),
            .I(N__58586));
    LocalMux I__14200 (
            .O(N__58616),
            .I(N__58586));
    InMux I__14199 (
            .O(N__58615),
            .I(N__58581));
    InMux I__14198 (
            .O(N__58614),
            .I(N__58578));
    Span4Mux_h I__14197 (
            .O(N__58611),
            .I(N__58575));
    InMux I__14196 (
            .O(N__58610),
            .I(N__58572));
    InMux I__14195 (
            .O(N__58609),
            .I(N__58567));
    InMux I__14194 (
            .O(N__58608),
            .I(N__58567));
    InMux I__14193 (
            .O(N__58607),
            .I(N__58564));
    Span4Mux_v I__14192 (
            .O(N__58602),
            .I(N__58557));
    Span4Mux_v I__14191 (
            .O(N__58599),
            .I(N__58557));
    LocalMux I__14190 (
            .O(N__58594),
            .I(N__58557));
    LocalMux I__14189 (
            .O(N__58591),
            .I(N__58552));
    Span4Mux_h I__14188 (
            .O(N__58586),
            .I(N__58552));
    InMux I__14187 (
            .O(N__58585),
            .I(N__58547));
    InMux I__14186 (
            .O(N__58584),
            .I(N__58547));
    LocalMux I__14185 (
            .O(N__58581),
            .I(comm_cmd_5));
    LocalMux I__14184 (
            .O(N__58578),
            .I(comm_cmd_5));
    Odrv4 I__14183 (
            .O(N__58575),
            .I(comm_cmd_5));
    LocalMux I__14182 (
            .O(N__58572),
            .I(comm_cmd_5));
    LocalMux I__14181 (
            .O(N__58567),
            .I(comm_cmd_5));
    LocalMux I__14180 (
            .O(N__58564),
            .I(comm_cmd_5));
    Odrv4 I__14179 (
            .O(N__58557),
            .I(comm_cmd_5));
    Odrv4 I__14178 (
            .O(N__58552),
            .I(comm_cmd_5));
    LocalMux I__14177 (
            .O(N__58547),
            .I(comm_cmd_5));
    InMux I__14176 (
            .O(N__58528),
            .I(N__58523));
    InMux I__14175 (
            .O(N__58527),
            .I(N__58516));
    InMux I__14174 (
            .O(N__58526),
            .I(N__58516));
    LocalMux I__14173 (
            .O(N__58523),
            .I(N__58512));
    InMux I__14172 (
            .O(N__58522),
            .I(N__58508));
    CascadeMux I__14171 (
            .O(N__58521),
            .I(N__58505));
    LocalMux I__14170 (
            .O(N__58516),
            .I(N__58502));
    InMux I__14169 (
            .O(N__58515),
            .I(N__58499));
    Span4Mux_v I__14168 (
            .O(N__58512),
            .I(N__58496));
    CascadeMux I__14167 (
            .O(N__58511),
            .I(N__58493));
    LocalMux I__14166 (
            .O(N__58508),
            .I(N__58488));
    InMux I__14165 (
            .O(N__58505),
            .I(N__58484));
    Span4Mux_v I__14164 (
            .O(N__58502),
            .I(N__58475));
    LocalMux I__14163 (
            .O(N__58499),
            .I(N__58475));
    Span4Mux_v I__14162 (
            .O(N__58496),
            .I(N__58475));
    InMux I__14161 (
            .O(N__58493),
            .I(N__58470));
    InMux I__14160 (
            .O(N__58492),
            .I(N__58470));
    CascadeMux I__14159 (
            .O(N__58491),
            .I(N__58466));
    Span4Mux_h I__14158 (
            .O(N__58488),
            .I(N__58463));
    InMux I__14157 (
            .O(N__58487),
            .I(N__58460));
    LocalMux I__14156 (
            .O(N__58484),
            .I(N__58457));
    InMux I__14155 (
            .O(N__58483),
            .I(N__58452));
    InMux I__14154 (
            .O(N__58482),
            .I(N__58452));
    Sp12to4 I__14153 (
            .O(N__58475),
            .I(N__58447));
    LocalMux I__14152 (
            .O(N__58470),
            .I(N__58447));
    InMux I__14151 (
            .O(N__58469),
            .I(N__58442));
    InMux I__14150 (
            .O(N__58466),
            .I(N__58442));
    Odrv4 I__14149 (
            .O(N__58463),
            .I(comm_cmd_4));
    LocalMux I__14148 (
            .O(N__58460),
            .I(comm_cmd_4));
    Odrv4 I__14147 (
            .O(N__58457),
            .I(comm_cmd_4));
    LocalMux I__14146 (
            .O(N__58452),
            .I(comm_cmd_4));
    Odrv12 I__14145 (
            .O(N__58447),
            .I(comm_cmd_4));
    LocalMux I__14144 (
            .O(N__58442),
            .I(comm_cmd_4));
    InMux I__14143 (
            .O(N__58429),
            .I(N__58426));
    LocalMux I__14142 (
            .O(N__58426),
            .I(n22365));
    CascadeMux I__14141 (
            .O(N__58423),
            .I(n22364_cascade_));
    InMux I__14140 (
            .O(N__58420),
            .I(N__58417));
    LocalMux I__14139 (
            .O(N__58417),
            .I(n48));
    CascadeMux I__14138 (
            .O(N__58414),
            .I(n22370_cascade_));
    InMux I__14137 (
            .O(N__58411),
            .I(N__58408));
    LocalMux I__14136 (
            .O(N__58408),
            .I(N__58404));
    InMux I__14135 (
            .O(N__58407),
            .I(N__58400));
    Span4Mux_h I__14134 (
            .O(N__58404),
            .I(N__58396));
    InMux I__14133 (
            .O(N__58403),
            .I(N__58393));
    LocalMux I__14132 (
            .O(N__58400),
            .I(N__58390));
    InMux I__14131 (
            .O(N__58399),
            .I(N__58387));
    Odrv4 I__14130 (
            .O(N__58396),
            .I(n7148));
    LocalMux I__14129 (
            .O(N__58393),
            .I(n7148));
    Odrv4 I__14128 (
            .O(N__58390),
            .I(n7148));
    LocalMux I__14127 (
            .O(N__58387),
            .I(n7148));
    InMux I__14126 (
            .O(N__58378),
            .I(N__58375));
    LocalMux I__14125 (
            .O(N__58375),
            .I(N__58372));
    Odrv4 I__14124 (
            .O(N__58372),
            .I(n22368));
    InMux I__14123 (
            .O(N__58369),
            .I(N__58366));
    LocalMux I__14122 (
            .O(N__58366),
            .I(N__58362));
    InMux I__14121 (
            .O(N__58365),
            .I(N__58359));
    Span4Mux_h I__14120 (
            .O(N__58362),
            .I(N__58356));
    LocalMux I__14119 (
            .O(N__58359),
            .I(N__58353));
    Odrv4 I__14118 (
            .O(N__58356),
            .I(n9_adj_1507));
    Odrv12 I__14117 (
            .O(N__58353),
            .I(n9_adj_1507));
    InMux I__14116 (
            .O(N__58348),
            .I(N__58345));
    LocalMux I__14115 (
            .O(N__58345),
            .I(N__58342));
    Span4Mux_v I__14114 (
            .O(N__58342),
            .I(N__58339));
    Span4Mux_h I__14113 (
            .O(N__58339),
            .I(N__58336));
    Span4Mux_h I__14112 (
            .O(N__58336),
            .I(N__58333));
    Odrv4 I__14111 (
            .O(N__58333),
            .I(n23387));
    CascadeMux I__14110 (
            .O(N__58330),
            .I(N__58327));
    InMux I__14109 (
            .O(N__58327),
            .I(N__58324));
    LocalMux I__14108 (
            .O(N__58324),
            .I(N__58321));
    Odrv4 I__14107 (
            .O(N__58321),
            .I(n23351));
    InMux I__14106 (
            .O(N__58318),
            .I(N__58315));
    LocalMux I__14105 (
            .O(N__58315),
            .I(n23495));
    InMux I__14104 (
            .O(N__58312),
            .I(N__58309));
    LocalMux I__14103 (
            .O(N__58309),
            .I(N__58306));
    Span4Mux_v I__14102 (
            .O(N__58306),
            .I(N__58303));
    Odrv4 I__14101 (
            .O(N__58303),
            .I(buf_data_iac_19));
    InMux I__14100 (
            .O(N__58300),
            .I(N__58297));
    LocalMux I__14099 (
            .O(N__58297),
            .I(N__58294));
    Odrv12 I__14098 (
            .O(N__58294),
            .I(n22642));
    CascadeMux I__14097 (
            .O(N__58291),
            .I(N__58288));
    InMux I__14096 (
            .O(N__58288),
            .I(N__58285));
    LocalMux I__14095 (
            .O(N__58285),
            .I(N__58282));
    Span4Mux_h I__14094 (
            .O(N__58282),
            .I(N__58279));
    Odrv4 I__14093 (
            .O(N__58279),
            .I(n23_adj_1791));
    InMux I__14092 (
            .O(N__58276),
            .I(N__58273));
    LocalMux I__14091 (
            .O(N__58273),
            .I(N__58270));
    Span4Mux_v I__14090 (
            .O(N__58270),
            .I(N__58267));
    Sp12to4 I__14089 (
            .O(N__58267),
            .I(N__58264));
    Span12Mux_h I__14088 (
            .O(N__58264),
            .I(N__58261));
    Odrv12 I__14087 (
            .O(N__58261),
            .I(n23501));
    CascadeMux I__14086 (
            .O(N__58258),
            .I(n23459_cascade_));
    InMux I__14085 (
            .O(N__58255),
            .I(N__58252));
    LocalMux I__14084 (
            .O(N__58252),
            .I(N__58249));
    Span4Mux_v I__14083 (
            .O(N__58249),
            .I(N__58246));
    Sp12to4 I__14082 (
            .O(N__58246),
            .I(N__58243));
    Span12Mux_h I__14081 (
            .O(N__58243),
            .I(N__58240));
    Odrv12 I__14080 (
            .O(N__58240),
            .I(n112_adj_1795));
    InMux I__14079 (
            .O(N__58237),
            .I(N__58234));
    LocalMux I__14078 (
            .O(N__58234),
            .I(n22492));
    CascadeMux I__14077 (
            .O(N__58231),
            .I(n6_adj_1657_cascade_));
    CascadeMux I__14076 (
            .O(N__58228),
            .I(n26_adj_1597_cascade_));
    CEMux I__14075 (
            .O(N__58225),
            .I(N__58222));
    LocalMux I__14074 (
            .O(N__58222),
            .I(N__58219));
    Odrv4 I__14073 (
            .O(N__58219),
            .I(n18_adj_1595));
    InMux I__14072 (
            .O(N__58216),
            .I(N__58213));
    LocalMux I__14071 (
            .O(N__58213),
            .I(n21908));
    InMux I__14070 (
            .O(N__58210),
            .I(N__58201));
    InMux I__14069 (
            .O(N__58209),
            .I(N__58194));
    InMux I__14068 (
            .O(N__58208),
            .I(N__58194));
    InMux I__14067 (
            .O(N__58207),
            .I(N__58194));
    CascadeMux I__14066 (
            .O(N__58206),
            .I(N__58189));
    CascadeMux I__14065 (
            .O(N__58205),
            .I(N__58182));
    InMux I__14064 (
            .O(N__58204),
            .I(N__58178));
    LocalMux I__14063 (
            .O(N__58201),
            .I(N__58173));
    LocalMux I__14062 (
            .O(N__58194),
            .I(N__58173));
    InMux I__14061 (
            .O(N__58193),
            .I(N__58170));
    InMux I__14060 (
            .O(N__58192),
            .I(N__58161));
    InMux I__14059 (
            .O(N__58189),
            .I(N__58161));
    InMux I__14058 (
            .O(N__58188),
            .I(N__58161));
    InMux I__14057 (
            .O(N__58187),
            .I(N__58161));
    InMux I__14056 (
            .O(N__58186),
            .I(N__58154));
    InMux I__14055 (
            .O(N__58185),
            .I(N__58154));
    InMux I__14054 (
            .O(N__58182),
            .I(N__58154));
    CascadeMux I__14053 (
            .O(N__58181),
            .I(N__58148));
    LocalMux I__14052 (
            .O(N__58178),
            .I(N__58144));
    Span4Mux_v I__14051 (
            .O(N__58173),
            .I(N__58141));
    LocalMux I__14050 (
            .O(N__58170),
            .I(N__58138));
    LocalMux I__14049 (
            .O(N__58161),
            .I(N__58133));
    LocalMux I__14048 (
            .O(N__58154),
            .I(N__58133));
    InMux I__14047 (
            .O(N__58153),
            .I(N__58129));
    InMux I__14046 (
            .O(N__58152),
            .I(N__58126));
    InMux I__14045 (
            .O(N__58151),
            .I(N__58119));
    InMux I__14044 (
            .O(N__58148),
            .I(N__58119));
    InMux I__14043 (
            .O(N__58147),
            .I(N__58119));
    Span4Mux_v I__14042 (
            .O(N__58144),
            .I(N__58114));
    Span4Mux_h I__14041 (
            .O(N__58141),
            .I(N__58107));
    Span4Mux_h I__14040 (
            .O(N__58138),
            .I(N__58107));
    Span4Mux_v I__14039 (
            .O(N__58133),
            .I(N__58107));
    CascadeMux I__14038 (
            .O(N__58132),
            .I(N__58104));
    LocalMux I__14037 (
            .O(N__58129),
            .I(N__58097));
    LocalMux I__14036 (
            .O(N__58126),
            .I(N__58097));
    LocalMux I__14035 (
            .O(N__58119),
            .I(N__58097));
    InMux I__14034 (
            .O(N__58118),
            .I(N__58092));
    InMux I__14033 (
            .O(N__58117),
            .I(N__58092));
    Span4Mux_v I__14032 (
            .O(N__58114),
            .I(N__58089));
    Span4Mux_h I__14031 (
            .O(N__58107),
            .I(N__58086));
    InMux I__14030 (
            .O(N__58104),
            .I(N__58083));
    Span4Mux_v I__14029 (
            .O(N__58097),
            .I(N__58080));
    LocalMux I__14028 (
            .O(N__58092),
            .I(N__58077));
    Span4Mux_v I__14027 (
            .O(N__58089),
            .I(N__58074));
    Sp12to4 I__14026 (
            .O(N__58086),
            .I(N__58071));
    LocalMux I__14025 (
            .O(N__58083),
            .I(N__58068));
    Sp12to4 I__14024 (
            .O(N__58080),
            .I(N__58063));
    Span12Mux_v I__14023 (
            .O(N__58077),
            .I(N__58063));
    Sp12to4 I__14022 (
            .O(N__58074),
            .I(N__58060));
    Span12Mux_s2_h I__14021 (
            .O(N__58071),
            .I(N__58055));
    Span12Mux_h I__14020 (
            .O(N__58068),
            .I(N__58055));
    Span12Mux_v I__14019 (
            .O(N__58063),
            .I(N__58052));
    Span12Mux_h I__14018 (
            .O(N__58060),
            .I(N__58047));
    Span12Mux_v I__14017 (
            .O(N__58055),
            .I(N__58047));
    Odrv12 I__14016 (
            .O(N__58052),
            .I(ICE_SPI_CE0));
    Odrv12 I__14015 (
            .O(N__58047),
            .I(ICE_SPI_CE0));
    InMux I__14014 (
            .O(N__58042),
            .I(N__58023));
    InMux I__14013 (
            .O(N__58041),
            .I(N__58023));
    InMux I__14012 (
            .O(N__58040),
            .I(N__58023));
    CascadeMux I__14011 (
            .O(N__58039),
            .I(N__58019));
    InMux I__14010 (
            .O(N__58038),
            .I(N__58011));
    InMux I__14009 (
            .O(N__58037),
            .I(N__58011));
    InMux I__14008 (
            .O(N__58036),
            .I(N__58011));
    InMux I__14007 (
            .O(N__58035),
            .I(N__58002));
    InMux I__14006 (
            .O(N__58034),
            .I(N__58002));
    InMux I__14005 (
            .O(N__58033),
            .I(N__58002));
    InMux I__14004 (
            .O(N__58032),
            .I(N__58002));
    InMux I__14003 (
            .O(N__58031),
            .I(N__57999));
    InMux I__14002 (
            .O(N__58030),
            .I(N__57996));
    LocalMux I__14001 (
            .O(N__58023),
            .I(N__57993));
    InMux I__14000 (
            .O(N__58022),
            .I(N__57990));
    InMux I__13999 (
            .O(N__58019),
            .I(N__57985));
    InMux I__13998 (
            .O(N__58018),
            .I(N__57985));
    LocalMux I__13997 (
            .O(N__58011),
            .I(comm_data_vld));
    LocalMux I__13996 (
            .O(N__58002),
            .I(comm_data_vld));
    LocalMux I__13995 (
            .O(N__57999),
            .I(comm_data_vld));
    LocalMux I__13994 (
            .O(N__57996),
            .I(comm_data_vld));
    Odrv4 I__13993 (
            .O(N__57993),
            .I(comm_data_vld));
    LocalMux I__13992 (
            .O(N__57990),
            .I(comm_data_vld));
    LocalMux I__13991 (
            .O(N__57985),
            .I(comm_data_vld));
    InMux I__13990 (
            .O(N__57970),
            .I(N__57967));
    LocalMux I__13989 (
            .O(N__57967),
            .I(N__57964));
    Span4Mux_h I__13988 (
            .O(N__57964),
            .I(N__57961));
    Odrv4 I__13987 (
            .O(N__57961),
            .I(n4_adj_1718));
    InMux I__13986 (
            .O(N__57958),
            .I(N__57954));
    CascadeMux I__13985 (
            .O(N__57957),
            .I(N__57950));
    LocalMux I__13984 (
            .O(N__57954),
            .I(N__57947));
    InMux I__13983 (
            .O(N__57953),
            .I(N__57942));
    InMux I__13982 (
            .O(N__57950),
            .I(N__57942));
    Odrv4 I__13981 (
            .O(N__57947),
            .I(req_data_cnt_11));
    LocalMux I__13980 (
            .O(N__57942),
            .I(req_data_cnt_11));
    InMux I__13979 (
            .O(N__57937),
            .I(N__57934));
    LocalMux I__13978 (
            .O(N__57934),
            .I(N__57931));
    Span4Mux_h I__13977 (
            .O(N__57931),
            .I(N__57928));
    Span4Mux_h I__13976 (
            .O(N__57928),
            .I(N__57925));
    Span4Mux_v I__13975 (
            .O(N__57925),
            .I(N__57922));
    Odrv4 I__13974 (
            .O(N__57922),
            .I(n112_adj_1777));
    InMux I__13973 (
            .O(N__57919),
            .I(N__57916));
    LocalMux I__13972 (
            .O(N__57916),
            .I(N__57913));
    Span12Mux_h I__13971 (
            .O(N__57913),
            .I(N__57910));
    Odrv12 I__13970 (
            .O(N__57910),
            .I(comm_buf_0_7_N_543_5));
    InMux I__13969 (
            .O(N__57907),
            .I(N__57900));
    InMux I__13968 (
            .O(N__57906),
            .I(N__57900));
    InMux I__13967 (
            .O(N__57905),
            .I(N__57897));
    LocalMux I__13966 (
            .O(N__57900),
            .I(n1373));
    LocalMux I__13965 (
            .O(N__57897),
            .I(n1373));
    CascadeMux I__13964 (
            .O(N__57892),
            .I(n2_cascade_));
    InMux I__13963 (
            .O(N__57889),
            .I(N__57886));
    LocalMux I__13962 (
            .O(N__57886),
            .I(N__57883));
    Odrv4 I__13961 (
            .O(N__57883),
            .I(n23342));
    CascadeMux I__13960 (
            .O(N__57880),
            .I(N__57873));
    InMux I__13959 (
            .O(N__57879),
            .I(N__57864));
    InMux I__13958 (
            .O(N__57878),
            .I(N__57864));
    InMux I__13957 (
            .O(N__57877),
            .I(N__57857));
    InMux I__13956 (
            .O(N__57876),
            .I(N__57845));
    InMux I__13955 (
            .O(N__57873),
            .I(N__57841));
    CascadeMux I__13954 (
            .O(N__57872),
            .I(N__57838));
    CascadeMux I__13953 (
            .O(N__57871),
            .I(N__57835));
    InMux I__13952 (
            .O(N__57870),
            .I(N__57830));
    CascadeMux I__13951 (
            .O(N__57869),
            .I(N__57827));
    LocalMux I__13950 (
            .O(N__57864),
            .I(N__57824));
    InMux I__13949 (
            .O(N__57863),
            .I(N__57821));
    InMux I__13948 (
            .O(N__57862),
            .I(N__57814));
    InMux I__13947 (
            .O(N__57861),
            .I(N__57814));
    InMux I__13946 (
            .O(N__57860),
            .I(N__57814));
    LocalMux I__13945 (
            .O(N__57857),
            .I(N__57811));
    InMux I__13944 (
            .O(N__57856),
            .I(N__57808));
    CascadeMux I__13943 (
            .O(N__57855),
            .I(N__57805));
    CascadeMux I__13942 (
            .O(N__57854),
            .I(N__57802));
    InMux I__13941 (
            .O(N__57853),
            .I(N__57799));
    InMux I__13940 (
            .O(N__57852),
            .I(N__57794));
    InMux I__13939 (
            .O(N__57851),
            .I(N__57794));
    InMux I__13938 (
            .O(N__57850),
            .I(N__57789));
    InMux I__13937 (
            .O(N__57849),
            .I(N__57789));
    InMux I__13936 (
            .O(N__57848),
            .I(N__57786));
    LocalMux I__13935 (
            .O(N__57845),
            .I(N__57783));
    CascadeMux I__13934 (
            .O(N__57844),
            .I(N__57780));
    LocalMux I__13933 (
            .O(N__57841),
            .I(N__57775));
    InMux I__13932 (
            .O(N__57838),
            .I(N__57772));
    InMux I__13931 (
            .O(N__57835),
            .I(N__57765));
    InMux I__13930 (
            .O(N__57834),
            .I(N__57765));
    InMux I__13929 (
            .O(N__57833),
            .I(N__57765));
    LocalMux I__13928 (
            .O(N__57830),
            .I(N__57760));
    InMux I__13927 (
            .O(N__57827),
            .I(N__57757));
    Span4Mux_v I__13926 (
            .O(N__57824),
            .I(N__57754));
    LocalMux I__13925 (
            .O(N__57821),
            .I(N__57751));
    LocalMux I__13924 (
            .O(N__57814),
            .I(N__57748));
    Span4Mux_h I__13923 (
            .O(N__57811),
            .I(N__57742));
    LocalMux I__13922 (
            .O(N__57808),
            .I(N__57736));
    InMux I__13921 (
            .O(N__57805),
            .I(N__57731));
    InMux I__13920 (
            .O(N__57802),
            .I(N__57731));
    LocalMux I__13919 (
            .O(N__57799),
            .I(N__57723));
    LocalMux I__13918 (
            .O(N__57794),
            .I(N__57723));
    LocalMux I__13917 (
            .O(N__57789),
            .I(N__57716));
    LocalMux I__13916 (
            .O(N__57786),
            .I(N__57716));
    Span4Mux_h I__13915 (
            .O(N__57783),
            .I(N__57716));
    InMux I__13914 (
            .O(N__57780),
            .I(N__57713));
    CascadeMux I__13913 (
            .O(N__57779),
            .I(N__57697));
    CascadeMux I__13912 (
            .O(N__57778),
            .I(N__57694));
    Span4Mux_h I__13911 (
            .O(N__57775),
            .I(N__57687));
    LocalMux I__13910 (
            .O(N__57772),
            .I(N__57687));
    LocalMux I__13909 (
            .O(N__57765),
            .I(N__57684));
    InMux I__13908 (
            .O(N__57764),
            .I(N__57681));
    CascadeMux I__13907 (
            .O(N__57763),
            .I(N__57678));
    Span4Mux_v I__13906 (
            .O(N__57760),
            .I(N__57673));
    LocalMux I__13905 (
            .O(N__57757),
            .I(N__57673));
    Span4Mux_v I__13904 (
            .O(N__57754),
            .I(N__57666));
    Span4Mux_v I__13903 (
            .O(N__57751),
            .I(N__57666));
    Span4Mux_v I__13902 (
            .O(N__57748),
            .I(N__57666));
    CascadeMux I__13901 (
            .O(N__57747),
            .I(N__57662));
    CascadeMux I__13900 (
            .O(N__57746),
            .I(N__57658));
    InMux I__13899 (
            .O(N__57745),
            .I(N__57655));
    Span4Mux_h I__13898 (
            .O(N__57742),
            .I(N__57652));
    InMux I__13897 (
            .O(N__57741),
            .I(N__57647));
    InMux I__13896 (
            .O(N__57740),
            .I(N__57647));
    InMux I__13895 (
            .O(N__57739),
            .I(N__57644));
    Span4Mux_h I__13894 (
            .O(N__57736),
            .I(N__57639));
    LocalMux I__13893 (
            .O(N__57731),
            .I(N__57639));
    InMux I__13892 (
            .O(N__57730),
            .I(N__57632));
    InMux I__13891 (
            .O(N__57729),
            .I(N__57632));
    InMux I__13890 (
            .O(N__57728),
            .I(N__57632));
    Span4Mux_v I__13889 (
            .O(N__57723),
            .I(N__57625));
    Span4Mux_v I__13888 (
            .O(N__57716),
            .I(N__57625));
    LocalMux I__13887 (
            .O(N__57713),
            .I(N__57625));
    InMux I__13886 (
            .O(N__57712),
            .I(N__57622));
    CascadeMux I__13885 (
            .O(N__57711),
            .I(N__57614));
    CascadeMux I__13884 (
            .O(N__57710),
            .I(N__57611));
    CascadeMux I__13883 (
            .O(N__57709),
            .I(N__57607));
    CascadeMux I__13882 (
            .O(N__57708),
            .I(N__57604));
    CascadeMux I__13881 (
            .O(N__57707),
            .I(N__57600));
    InMux I__13880 (
            .O(N__57706),
            .I(N__57591));
    InMux I__13879 (
            .O(N__57705),
            .I(N__57591));
    InMux I__13878 (
            .O(N__57704),
            .I(N__57591));
    InMux I__13877 (
            .O(N__57703),
            .I(N__57591));
    InMux I__13876 (
            .O(N__57702),
            .I(N__57588));
    CascadeMux I__13875 (
            .O(N__57701),
            .I(N__57584));
    InMux I__13874 (
            .O(N__57700),
            .I(N__57571));
    InMux I__13873 (
            .O(N__57697),
            .I(N__57571));
    InMux I__13872 (
            .O(N__57694),
            .I(N__57571));
    InMux I__13871 (
            .O(N__57693),
            .I(N__57571));
    InMux I__13870 (
            .O(N__57692),
            .I(N__57571));
    Span4Mux_h I__13869 (
            .O(N__57687),
            .I(N__57566));
    Span4Mux_h I__13868 (
            .O(N__57684),
            .I(N__57566));
    LocalMux I__13867 (
            .O(N__57681),
            .I(N__57563));
    InMux I__13866 (
            .O(N__57678),
            .I(N__57560));
    Sp12to4 I__13865 (
            .O(N__57673),
            .I(N__57557));
    Span4Mux_h I__13864 (
            .O(N__57666),
            .I(N__57554));
    InMux I__13863 (
            .O(N__57665),
            .I(N__57551));
    InMux I__13862 (
            .O(N__57662),
            .I(N__57546));
    InMux I__13861 (
            .O(N__57661),
            .I(N__57546));
    InMux I__13860 (
            .O(N__57658),
            .I(N__57543));
    LocalMux I__13859 (
            .O(N__57655),
            .I(N__57540));
    Span4Mux_h I__13858 (
            .O(N__57652),
            .I(N__57535));
    LocalMux I__13857 (
            .O(N__57647),
            .I(N__57535));
    LocalMux I__13856 (
            .O(N__57644),
            .I(N__57532));
    Span4Mux_h I__13855 (
            .O(N__57639),
            .I(N__57527));
    LocalMux I__13854 (
            .O(N__57632),
            .I(N__57527));
    Span4Mux_h I__13853 (
            .O(N__57625),
            .I(N__57522));
    LocalMux I__13852 (
            .O(N__57622),
            .I(N__57522));
    InMux I__13851 (
            .O(N__57621),
            .I(N__57517));
    InMux I__13850 (
            .O(N__57620),
            .I(N__57514));
    InMux I__13849 (
            .O(N__57619),
            .I(N__57509));
    InMux I__13848 (
            .O(N__57618),
            .I(N__57509));
    InMux I__13847 (
            .O(N__57617),
            .I(N__57506));
    InMux I__13846 (
            .O(N__57614),
            .I(N__57501));
    InMux I__13845 (
            .O(N__57611),
            .I(N__57501));
    InMux I__13844 (
            .O(N__57610),
            .I(N__57498));
    InMux I__13843 (
            .O(N__57607),
            .I(N__57489));
    InMux I__13842 (
            .O(N__57604),
            .I(N__57489));
    InMux I__13841 (
            .O(N__57603),
            .I(N__57489));
    InMux I__13840 (
            .O(N__57600),
            .I(N__57489));
    LocalMux I__13839 (
            .O(N__57591),
            .I(N__57484));
    LocalMux I__13838 (
            .O(N__57588),
            .I(N__57484));
    InMux I__13837 (
            .O(N__57587),
            .I(N__57475));
    InMux I__13836 (
            .O(N__57584),
            .I(N__57475));
    InMux I__13835 (
            .O(N__57583),
            .I(N__57475));
    InMux I__13834 (
            .O(N__57582),
            .I(N__57475));
    LocalMux I__13833 (
            .O(N__57571),
            .I(N__57472));
    Sp12to4 I__13832 (
            .O(N__57566),
            .I(N__57469));
    Span4Mux_h I__13831 (
            .O(N__57563),
            .I(N__57465));
    LocalMux I__13830 (
            .O(N__57560),
            .I(N__57462));
    Span12Mux_v I__13829 (
            .O(N__57557),
            .I(N__57455));
    Sp12to4 I__13828 (
            .O(N__57554),
            .I(N__57455));
    LocalMux I__13827 (
            .O(N__57551),
            .I(N__57455));
    LocalMux I__13826 (
            .O(N__57546),
            .I(N__57450));
    LocalMux I__13825 (
            .O(N__57543),
            .I(N__57450));
    Span4Mux_v I__13824 (
            .O(N__57540),
            .I(N__57445));
    Span4Mux_h I__13823 (
            .O(N__57535),
            .I(N__57445));
    Span4Mux_h I__13822 (
            .O(N__57532),
            .I(N__57438));
    Span4Mux_v I__13821 (
            .O(N__57527),
            .I(N__57438));
    Span4Mux_h I__13820 (
            .O(N__57522),
            .I(N__57438));
    InMux I__13819 (
            .O(N__57521),
            .I(N__57435));
    InMux I__13818 (
            .O(N__57520),
            .I(N__57432));
    LocalMux I__13817 (
            .O(N__57517),
            .I(N__57429));
    LocalMux I__13816 (
            .O(N__57514),
            .I(N__57408));
    LocalMux I__13815 (
            .O(N__57509),
            .I(N__57408));
    LocalMux I__13814 (
            .O(N__57506),
            .I(N__57408));
    LocalMux I__13813 (
            .O(N__57501),
            .I(N__57408));
    LocalMux I__13812 (
            .O(N__57498),
            .I(N__57408));
    LocalMux I__13811 (
            .O(N__57489),
            .I(N__57408));
    Sp12to4 I__13810 (
            .O(N__57484),
            .I(N__57408));
    LocalMux I__13809 (
            .O(N__57475),
            .I(N__57408));
    Sp12to4 I__13808 (
            .O(N__57472),
            .I(N__57408));
    Span12Mux_s6_v I__13807 (
            .O(N__57469),
            .I(N__57408));
    InMux I__13806 (
            .O(N__57468),
            .I(N__57405));
    Span4Mux_h I__13805 (
            .O(N__57465),
            .I(N__57400));
    Span4Mux_v I__13804 (
            .O(N__57462),
            .I(N__57400));
    Span12Mux_h I__13803 (
            .O(N__57455),
            .I(N__57397));
    Span12Mux_h I__13802 (
            .O(N__57450),
            .I(N__57394));
    Span4Mux_h I__13801 (
            .O(N__57445),
            .I(N__57389));
    Span4Mux_v I__13800 (
            .O(N__57438),
            .I(N__57389));
    LocalMux I__13799 (
            .O(N__57435),
            .I(N__57380));
    LocalMux I__13798 (
            .O(N__57432),
            .I(N__57380));
    Span12Mux_h I__13797 (
            .O(N__57429),
            .I(N__57380));
    Span12Mux_v I__13796 (
            .O(N__57408),
            .I(N__57380));
    LocalMux I__13795 (
            .O(N__57405),
            .I(n9837));
    Odrv4 I__13794 (
            .O(N__57400),
            .I(n9837));
    Odrv12 I__13793 (
            .O(N__57397),
            .I(n9837));
    Odrv12 I__13792 (
            .O(N__57394),
            .I(n9837));
    Odrv4 I__13791 (
            .O(N__57389),
            .I(n9837));
    Odrv12 I__13790 (
            .O(N__57380),
            .I(n9837));
    CascadeMux I__13789 (
            .O(N__57367),
            .I(n23345_cascade_));
    InMux I__13788 (
            .O(N__57364),
            .I(N__57361));
    LocalMux I__13787 (
            .O(N__57361),
            .I(n8_adj_1659));
    InMux I__13786 (
            .O(N__57358),
            .I(N__57355));
    LocalMux I__13785 (
            .O(N__57355),
            .I(N__57350));
    InMux I__13784 (
            .O(N__57354),
            .I(N__57347));
    InMux I__13783 (
            .O(N__57353),
            .I(N__57344));
    Odrv4 I__13782 (
            .O(N__57350),
            .I(n2562));
    LocalMux I__13781 (
            .O(N__57347),
            .I(n2562));
    LocalMux I__13780 (
            .O(N__57344),
            .I(n2562));
    InMux I__13779 (
            .O(N__57337),
            .I(N__57334));
    LocalMux I__13778 (
            .O(N__57334),
            .I(N__57331));
    Odrv4 I__13777 (
            .O(N__57331),
            .I(n22339));
    CascadeMux I__13776 (
            .O(N__57328),
            .I(n22340_cascade_));
    CEMux I__13775 (
            .O(N__57325),
            .I(N__57322));
    LocalMux I__13774 (
            .O(N__57322),
            .I(N__57319));
    Span4Mux_h I__13773 (
            .O(N__57319),
            .I(N__57316));
    Span4Mux_h I__13772 (
            .O(N__57316),
            .I(N__57313));
    Odrv4 I__13771 (
            .O(N__57313),
            .I(n14_adj_1593));
    CascadeMux I__13770 (
            .O(N__57310),
            .I(N__57307));
    InMux I__13769 (
            .O(N__57307),
            .I(N__57304));
    LocalMux I__13768 (
            .O(N__57304),
            .I(N__57301));
    Span4Mux_h I__13767 (
            .O(N__57301),
            .I(N__57296));
    InMux I__13766 (
            .O(N__57300),
            .I(N__57293));
    InMux I__13765 (
            .O(N__57299),
            .I(N__57290));
    Odrv4 I__13764 (
            .O(N__57296),
            .I(n5));
    LocalMux I__13763 (
            .O(N__57293),
            .I(n5));
    LocalMux I__13762 (
            .O(N__57290),
            .I(n5));
    CascadeMux I__13761 (
            .O(N__57283),
            .I(n9725_cascade_));
    InMux I__13760 (
            .O(N__57280),
            .I(N__57277));
    LocalMux I__13759 (
            .O(N__57277),
            .I(N__57274));
    Span4Mux_h I__13758 (
            .O(N__57274),
            .I(N__57271));
    Odrv4 I__13757 (
            .O(N__57271),
            .I(n4));
    InMux I__13756 (
            .O(N__57268),
            .I(N__57265));
    LocalMux I__13755 (
            .O(N__57265),
            .I(\ADC_VDC.genclk.n28_adj_1481 ));
    CascadeMux I__13754 (
            .O(N__57262),
            .I(N__57258));
    InMux I__13753 (
            .O(N__57261),
            .I(N__57255));
    InMux I__13752 (
            .O(N__57258),
            .I(N__57252));
    LocalMux I__13751 (
            .O(N__57255),
            .I(N__57249));
    LocalMux I__13750 (
            .O(N__57252),
            .I(\ADC_VDC.genclk.t0on_13 ));
    Odrv4 I__13749 (
            .O(N__57249),
            .I(\ADC_VDC.genclk.t0on_13 ));
    InMux I__13748 (
            .O(N__57244),
            .I(N__57240));
    InMux I__13747 (
            .O(N__57243),
            .I(N__57237));
    LocalMux I__13746 (
            .O(N__57240),
            .I(\ADC_VDC.genclk.t0on_3 ));
    LocalMux I__13745 (
            .O(N__57237),
            .I(\ADC_VDC.genclk.t0on_3 ));
    CascadeMux I__13744 (
            .O(N__57232),
            .I(N__57228));
    InMux I__13743 (
            .O(N__57231),
            .I(N__57225));
    InMux I__13742 (
            .O(N__57228),
            .I(N__57222));
    LocalMux I__13741 (
            .O(N__57225),
            .I(\ADC_VDC.genclk.t0on_5 ));
    LocalMux I__13740 (
            .O(N__57222),
            .I(\ADC_VDC.genclk.t0on_5 ));
    InMux I__13739 (
            .O(N__57217),
            .I(N__57213));
    InMux I__13738 (
            .O(N__57216),
            .I(N__57210));
    LocalMux I__13737 (
            .O(N__57213),
            .I(\ADC_VDC.genclk.t0on_8 ));
    LocalMux I__13736 (
            .O(N__57210),
            .I(\ADC_VDC.genclk.t0on_8 ));
    InMux I__13735 (
            .O(N__57205),
            .I(N__57202));
    LocalMux I__13734 (
            .O(N__57202),
            .I(\ADC_VDC.genclk.n26_adj_1482 ));
    CEMux I__13733 (
            .O(N__57199),
            .I(N__57196));
    LocalMux I__13732 (
            .O(N__57196),
            .I(N__57192));
    CEMux I__13731 (
            .O(N__57195),
            .I(N__57189));
    Span4Mux_h I__13730 (
            .O(N__57192),
            .I(N__57186));
    LocalMux I__13729 (
            .O(N__57189),
            .I(N__57183));
    Odrv4 I__13728 (
            .O(N__57186),
            .I(\ADC_VDC.genclk.div_state_1__N_1480 ));
    Odrv12 I__13727 (
            .O(N__57183),
            .I(\ADC_VDC.genclk.div_state_1__N_1480 ));
    InMux I__13726 (
            .O(N__57178),
            .I(N__57167));
    InMux I__13725 (
            .O(N__57177),
            .I(N__57164));
    InMux I__13724 (
            .O(N__57176),
            .I(N__57161));
    InMux I__13723 (
            .O(N__57175),
            .I(N__57148));
    InMux I__13722 (
            .O(N__57174),
            .I(N__57148));
    InMux I__13721 (
            .O(N__57173),
            .I(N__57148));
    InMux I__13720 (
            .O(N__57172),
            .I(N__57148));
    InMux I__13719 (
            .O(N__57171),
            .I(N__57148));
    InMux I__13718 (
            .O(N__57170),
            .I(N__57148));
    LocalMux I__13717 (
            .O(N__57167),
            .I(N__57138));
    LocalMux I__13716 (
            .O(N__57164),
            .I(N__57138));
    LocalMux I__13715 (
            .O(N__57161),
            .I(N__57138));
    LocalMux I__13714 (
            .O(N__57148),
            .I(N__57138));
    CascadeMux I__13713 (
            .O(N__57147),
            .I(N__57132));
    Span4Mux_v I__13712 (
            .O(N__57138),
            .I(N__57126));
    InMux I__13711 (
            .O(N__57137),
            .I(N__57123));
    InMux I__13710 (
            .O(N__57136),
            .I(N__57100));
    InMux I__13709 (
            .O(N__57135),
            .I(N__57100));
    InMux I__13708 (
            .O(N__57132),
            .I(N__57100));
    InMux I__13707 (
            .O(N__57131),
            .I(N__57100));
    InMux I__13706 (
            .O(N__57130),
            .I(N__57097));
    InMux I__13705 (
            .O(N__57129),
            .I(N__57093));
    Span4Mux_h I__13704 (
            .O(N__57126),
            .I(N__57087));
    LocalMux I__13703 (
            .O(N__57123),
            .I(N__57087));
    SRMux I__13702 (
            .O(N__57122),
            .I(N__57084));
    InMux I__13701 (
            .O(N__57121),
            .I(N__57079));
    InMux I__13700 (
            .O(N__57120),
            .I(N__57079));
    InMux I__13699 (
            .O(N__57119),
            .I(N__57074));
    InMux I__13698 (
            .O(N__57118),
            .I(N__57071));
    InMux I__13697 (
            .O(N__57117),
            .I(N__57063));
    InMux I__13696 (
            .O(N__57116),
            .I(N__57063));
    InMux I__13695 (
            .O(N__57115),
            .I(N__57063));
    InMux I__13694 (
            .O(N__57114),
            .I(N__57058));
    InMux I__13693 (
            .O(N__57113),
            .I(N__57058));
    InMux I__13692 (
            .O(N__57112),
            .I(N__57053));
    InMux I__13691 (
            .O(N__57111),
            .I(N__57053));
    InMux I__13690 (
            .O(N__57110),
            .I(N__57050));
    InMux I__13689 (
            .O(N__57109),
            .I(N__57046));
    LocalMux I__13688 (
            .O(N__57100),
            .I(N__57043));
    LocalMux I__13687 (
            .O(N__57097),
            .I(N__57040));
    InMux I__13686 (
            .O(N__57096),
            .I(N__57037));
    LocalMux I__13685 (
            .O(N__57093),
            .I(N__57034));
    SRMux I__13684 (
            .O(N__57092),
            .I(N__57031));
    Span4Mux_v I__13683 (
            .O(N__57087),
            .I(N__57028));
    LocalMux I__13682 (
            .O(N__57084),
            .I(N__57025));
    LocalMux I__13681 (
            .O(N__57079),
            .I(N__57022));
    SRMux I__13680 (
            .O(N__57078),
            .I(N__57019));
    InMux I__13679 (
            .O(N__57077),
            .I(N__57016));
    LocalMux I__13678 (
            .O(N__57074),
            .I(N__57011));
    LocalMux I__13677 (
            .O(N__57071),
            .I(N__57011));
    InMux I__13676 (
            .O(N__57070),
            .I(N__57008));
    LocalMux I__13675 (
            .O(N__57063),
            .I(N__57003));
    LocalMux I__13674 (
            .O(N__57058),
            .I(N__57003));
    LocalMux I__13673 (
            .O(N__57053),
            .I(N__57000));
    LocalMux I__13672 (
            .O(N__57050),
            .I(N__56997));
    InMux I__13671 (
            .O(N__57049),
            .I(N__56994));
    LocalMux I__13670 (
            .O(N__57046),
            .I(N__56989));
    Span4Mux_v I__13669 (
            .O(N__57043),
            .I(N__56989));
    Span4Mux_h I__13668 (
            .O(N__57040),
            .I(N__56984));
    LocalMux I__13667 (
            .O(N__57037),
            .I(N__56984));
    Span4Mux_h I__13666 (
            .O(N__57034),
            .I(N__56979));
    LocalMux I__13665 (
            .O(N__57031),
            .I(N__56979));
    Span4Mux_h I__13664 (
            .O(N__57028),
            .I(N__56972));
    Span4Mux_v I__13663 (
            .O(N__57025),
            .I(N__56972));
    Span4Mux_v I__13662 (
            .O(N__57022),
            .I(N__56972));
    LocalMux I__13661 (
            .O(N__57019),
            .I(N__56969));
    LocalMux I__13660 (
            .O(N__57016),
            .I(N__56962));
    Span4Mux_v I__13659 (
            .O(N__57011),
            .I(N__56962));
    LocalMux I__13658 (
            .O(N__57008),
            .I(N__56962));
    Span4Mux_v I__13657 (
            .O(N__57003),
            .I(N__56957));
    Span4Mux_v I__13656 (
            .O(N__57000),
            .I(N__56957));
    Span4Mux_v I__13655 (
            .O(N__56997),
            .I(N__56950));
    LocalMux I__13654 (
            .O(N__56994),
            .I(N__56950));
    Span4Mux_h I__13653 (
            .O(N__56989),
            .I(N__56950));
    Span4Mux_h I__13652 (
            .O(N__56984),
            .I(N__56947));
    Span4Mux_v I__13651 (
            .O(N__56979),
            .I(N__56938));
    Span4Mux_h I__13650 (
            .O(N__56972),
            .I(N__56938));
    Span4Mux_v I__13649 (
            .O(N__56969),
            .I(N__56938));
    Span4Mux_h I__13648 (
            .O(N__56962),
            .I(N__56938));
    Span4Mux_h I__13647 (
            .O(N__56957),
            .I(N__56933));
    Span4Mux_h I__13646 (
            .O(N__56950),
            .I(N__56933));
    Odrv4 I__13645 (
            .O(N__56947),
            .I(comm_clear));
    Odrv4 I__13644 (
            .O(N__56938),
            .I(comm_clear));
    Odrv4 I__13643 (
            .O(N__56933),
            .I(comm_clear));
    InMux I__13642 (
            .O(N__56926),
            .I(N__56923));
    LocalMux I__13641 (
            .O(N__56923),
            .I(N__56920));
    Odrv4 I__13640 (
            .O(N__56920),
            .I(buf_data_iac_18));
    CascadeMux I__13639 (
            .O(N__56917),
            .I(N__56914));
    InMux I__13638 (
            .O(N__56914),
            .I(N__56911));
    LocalMux I__13637 (
            .O(N__56911),
            .I(N__56908));
    Span4Mux_h I__13636 (
            .O(N__56908),
            .I(N__56905));
    Span4Mux_h I__13635 (
            .O(N__56905),
            .I(N__56902));
    Span4Mux_v I__13634 (
            .O(N__56902),
            .I(N__56899));
    Odrv4 I__13633 (
            .O(N__56899),
            .I(n22170));
    CEMux I__13632 (
            .O(N__56896),
            .I(N__56893));
    LocalMux I__13631 (
            .O(N__56893),
            .I(N__56890));
    Span4Mux_h I__13630 (
            .O(N__56890),
            .I(N__56887));
    Odrv4 I__13629 (
            .O(N__56887),
            .I(n12035));
    InMux I__13628 (
            .O(N__56884),
            .I(N__56881));
    LocalMux I__13627 (
            .O(N__56881),
            .I(N__56878));
    Odrv12 I__13626 (
            .O(N__56878),
            .I(n7_adj_1687));
    InMux I__13625 (
            .O(N__56875),
            .I(N__56872));
    LocalMux I__13624 (
            .O(N__56872),
            .I(N__56868));
    InMux I__13623 (
            .O(N__56871),
            .I(N__56865));
    Span4Mux_h I__13622 (
            .O(N__56868),
            .I(N__56862));
    LocalMux I__13621 (
            .O(N__56865),
            .I(N__56859));
    Odrv4 I__13620 (
            .O(N__56862),
            .I(comm_state_3_N_484_3));
    Odrv4 I__13619 (
            .O(N__56859),
            .I(comm_state_3_N_484_3));
    InMux I__13618 (
            .O(N__56854),
            .I(N__56851));
    LocalMux I__13617 (
            .O(N__56851),
            .I(N__56846));
    InMux I__13616 (
            .O(N__56850),
            .I(N__56843));
    InMux I__13615 (
            .O(N__56849),
            .I(N__56840));
    Span4Mux_h I__13614 (
            .O(N__56846),
            .I(N__56835));
    LocalMux I__13613 (
            .O(N__56843),
            .I(N__56831));
    LocalMux I__13612 (
            .O(N__56840),
            .I(N__56828));
    InMux I__13611 (
            .O(N__56839),
            .I(N__56825));
    InMux I__13610 (
            .O(N__56838),
            .I(N__56822));
    Span4Mux_h I__13609 (
            .O(N__56835),
            .I(N__56819));
    InMux I__13608 (
            .O(N__56834),
            .I(N__56816));
    Span12Mux_v I__13607 (
            .O(N__56831),
            .I(N__56813));
    Span4Mux_h I__13606 (
            .O(N__56828),
            .I(N__56810));
    LocalMux I__13605 (
            .O(N__56825),
            .I(N__56807));
    LocalMux I__13604 (
            .O(N__56822),
            .I(N__56804));
    Span4Mux_v I__13603 (
            .O(N__56819),
            .I(N__56799));
    LocalMux I__13602 (
            .O(N__56816),
            .I(N__56799));
    Span12Mux_h I__13601 (
            .O(N__56813),
            .I(N__56796));
    Span4Mux_h I__13600 (
            .O(N__56810),
            .I(N__56793));
    Span4Mux_h I__13599 (
            .O(N__56807),
            .I(N__56790));
    Span4Mux_v I__13598 (
            .O(N__56804),
            .I(N__56785));
    Span4Mux_h I__13597 (
            .O(N__56799),
            .I(N__56785));
    Odrv12 I__13596 (
            .O(N__56796),
            .I(n14_adj_1654));
    Odrv4 I__13595 (
            .O(N__56793),
            .I(n14_adj_1654));
    Odrv4 I__13594 (
            .O(N__56790),
            .I(n14_adj_1654));
    Odrv4 I__13593 (
            .O(N__56785),
            .I(n14_adj_1654));
    CEMux I__13592 (
            .O(N__56776),
            .I(N__56773));
    LocalMux I__13591 (
            .O(N__56773),
            .I(N__56770));
    Odrv4 I__13590 (
            .O(N__56770),
            .I(\ADC_VDC.genclk.n6 ));
    CascadeMux I__13589 (
            .O(N__56767),
            .I(N__56764));
    InMux I__13588 (
            .O(N__56764),
            .I(N__56760));
    InMux I__13587 (
            .O(N__56763),
            .I(N__56757));
    LocalMux I__13586 (
            .O(N__56760),
            .I(\ADC_VDC.genclk.t0on_6 ));
    LocalMux I__13585 (
            .O(N__56757),
            .I(\ADC_VDC.genclk.t0on_6 ));
    InMux I__13584 (
            .O(N__56752),
            .I(N__56748));
    InMux I__13583 (
            .O(N__56751),
            .I(N__56745));
    LocalMux I__13582 (
            .O(N__56748),
            .I(\ADC_VDC.genclk.t0on_1 ));
    LocalMux I__13581 (
            .O(N__56745),
            .I(\ADC_VDC.genclk.t0on_1 ));
    CascadeMux I__13580 (
            .O(N__56740),
            .I(N__56736));
    CascadeMux I__13579 (
            .O(N__56739),
            .I(N__56733));
    InMux I__13578 (
            .O(N__56736),
            .I(N__56730));
    InMux I__13577 (
            .O(N__56733),
            .I(N__56727));
    LocalMux I__13576 (
            .O(N__56730),
            .I(\ADC_VDC.genclk.t0on_4 ));
    LocalMux I__13575 (
            .O(N__56727),
            .I(\ADC_VDC.genclk.t0on_4 ));
    InMux I__13574 (
            .O(N__56722),
            .I(N__56718));
    InMux I__13573 (
            .O(N__56721),
            .I(N__56715));
    LocalMux I__13572 (
            .O(N__56718),
            .I(\ADC_VDC.genclk.t0on_0 ));
    LocalMux I__13571 (
            .O(N__56715),
            .I(\ADC_VDC.genclk.t0on_0 ));
    CascadeMux I__13570 (
            .O(N__56710),
            .I(\ADC_VDC.genclk.n22308_cascade_ ));
    InMux I__13569 (
            .O(N__56707),
            .I(N__56703));
    InMux I__13568 (
            .O(N__56706),
            .I(N__56700));
    LocalMux I__13567 (
            .O(N__56703),
            .I(N__56697));
    LocalMux I__13566 (
            .O(N__56700),
            .I(\ADC_VDC.genclk.t0on_12 ));
    Odrv4 I__13565 (
            .O(N__56697),
            .I(\ADC_VDC.genclk.t0on_12 ));
    CascadeMux I__13564 (
            .O(N__56692),
            .I(N__56689));
    InMux I__13563 (
            .O(N__56689),
            .I(N__56685));
    InMux I__13562 (
            .O(N__56688),
            .I(N__56682));
    LocalMux I__13561 (
            .O(N__56685),
            .I(\ADC_VDC.genclk.t0on_2 ));
    LocalMux I__13560 (
            .O(N__56682),
            .I(\ADC_VDC.genclk.t0on_2 ));
    CascadeMux I__13559 (
            .O(N__56677),
            .I(N__56673));
    InMux I__13558 (
            .O(N__56676),
            .I(N__56670));
    InMux I__13557 (
            .O(N__56673),
            .I(N__56667));
    LocalMux I__13556 (
            .O(N__56670),
            .I(\ADC_VDC.genclk.t0on_7 ));
    LocalMux I__13555 (
            .O(N__56667),
            .I(\ADC_VDC.genclk.t0on_7 ));
    InMux I__13554 (
            .O(N__56662),
            .I(N__56658));
    InMux I__13553 (
            .O(N__56661),
            .I(N__56655));
    LocalMux I__13552 (
            .O(N__56658),
            .I(\ADC_VDC.genclk.t0on_10 ));
    LocalMux I__13551 (
            .O(N__56655),
            .I(\ADC_VDC.genclk.t0on_10 ));
    InMux I__13550 (
            .O(N__56650),
            .I(N__56647));
    LocalMux I__13549 (
            .O(N__56647),
            .I(\ADC_VDC.genclk.n27_adj_1483 ));
    InMux I__13548 (
            .O(N__56644),
            .I(N__56640));
    InMux I__13547 (
            .O(N__56643),
            .I(N__56637));
    LocalMux I__13546 (
            .O(N__56640),
            .I(\ADC_VDC.genclk.t0on_14 ));
    LocalMux I__13545 (
            .O(N__56637),
            .I(\ADC_VDC.genclk.t0on_14 ));
    CascadeMux I__13544 (
            .O(N__56632),
            .I(N__56629));
    InMux I__13543 (
            .O(N__56629),
            .I(N__56625));
    InMux I__13542 (
            .O(N__56628),
            .I(N__56622));
    LocalMux I__13541 (
            .O(N__56625),
            .I(\ADC_VDC.genclk.t0on_9 ));
    LocalMux I__13540 (
            .O(N__56622),
            .I(\ADC_VDC.genclk.t0on_9 ));
    CascadeMux I__13539 (
            .O(N__56617),
            .I(N__56613));
    InMux I__13538 (
            .O(N__56616),
            .I(N__56610));
    InMux I__13537 (
            .O(N__56613),
            .I(N__56607));
    LocalMux I__13536 (
            .O(N__56610),
            .I(\ADC_VDC.genclk.t0on_15 ));
    LocalMux I__13535 (
            .O(N__56607),
            .I(\ADC_VDC.genclk.t0on_15 ));
    CascadeMux I__13534 (
            .O(N__56602),
            .I(N__56599));
    InMux I__13533 (
            .O(N__56599),
            .I(N__56595));
    InMux I__13532 (
            .O(N__56598),
            .I(N__56592));
    LocalMux I__13531 (
            .O(N__56595),
            .I(\ADC_VDC.genclk.t0on_11 ));
    LocalMux I__13530 (
            .O(N__56592),
            .I(\ADC_VDC.genclk.t0on_11 ));
    InMux I__13529 (
            .O(N__56587),
            .I(N__56584));
    LocalMux I__13528 (
            .O(N__56584),
            .I(N__56579));
    InMux I__13527 (
            .O(N__56583),
            .I(N__56574));
    CascadeMux I__13526 (
            .O(N__56582),
            .I(N__56571));
    Span4Mux_v I__13525 (
            .O(N__56579),
            .I(N__56566));
    InMux I__13524 (
            .O(N__56578),
            .I(N__56563));
    InMux I__13523 (
            .O(N__56577),
            .I(N__56560));
    LocalMux I__13522 (
            .O(N__56574),
            .I(N__56557));
    InMux I__13521 (
            .O(N__56571),
            .I(N__56554));
    InMux I__13520 (
            .O(N__56570),
            .I(N__56551));
    InMux I__13519 (
            .O(N__56569),
            .I(N__56548));
    Span4Mux_h I__13518 (
            .O(N__56566),
            .I(N__56543));
    LocalMux I__13517 (
            .O(N__56563),
            .I(N__56543));
    LocalMux I__13516 (
            .O(N__56560),
            .I(N__56540));
    Span4Mux_v I__13515 (
            .O(N__56557),
            .I(N__56533));
    LocalMux I__13514 (
            .O(N__56554),
            .I(N__56533));
    LocalMux I__13513 (
            .O(N__56551),
            .I(N__56533));
    LocalMux I__13512 (
            .O(N__56548),
            .I(N__56529));
    Span4Mux_h I__13511 (
            .O(N__56543),
            .I(N__56526));
    Span4Mux_v I__13510 (
            .O(N__56540),
            .I(N__56521));
    Span4Mux_h I__13509 (
            .O(N__56533),
            .I(N__56521));
    InMux I__13508 (
            .O(N__56532),
            .I(N__56518));
    Span12Mux_h I__13507 (
            .O(N__56529),
            .I(N__56515));
    Span4Mux_v I__13506 (
            .O(N__56526),
            .I(N__56508));
    Span4Mux_h I__13505 (
            .O(N__56521),
            .I(N__56508));
    LocalMux I__13504 (
            .O(N__56518),
            .I(N__56508));
    Odrv12 I__13503 (
            .O(N__56515),
            .I(comm_buf_1_5));
    Odrv4 I__13502 (
            .O(N__56508),
            .I(comm_buf_1_5));
    InMux I__13501 (
            .O(N__56503),
            .I(N__56499));
    InMux I__13500 (
            .O(N__56502),
            .I(N__56496));
    LocalMux I__13499 (
            .O(N__56499),
            .I(N__56490));
    LocalMux I__13498 (
            .O(N__56496),
            .I(N__56490));
    InMux I__13497 (
            .O(N__56495),
            .I(N__56487));
    Span12Mux_h I__13496 (
            .O(N__56490),
            .I(N__56484));
    LocalMux I__13495 (
            .O(N__56487),
            .I(data_index_5));
    Odrv12 I__13494 (
            .O(N__56484),
            .I(data_index_5));
    InMux I__13493 (
            .O(N__56479),
            .I(N__56475));
    InMux I__13492 (
            .O(N__56478),
            .I(N__56470));
    LocalMux I__13491 (
            .O(N__56475),
            .I(N__56466));
    InMux I__13490 (
            .O(N__56474),
            .I(N__56463));
    InMux I__13489 (
            .O(N__56473),
            .I(N__56455));
    LocalMux I__13488 (
            .O(N__56470),
            .I(N__56452));
    InMux I__13487 (
            .O(N__56469),
            .I(N__56448));
    Span4Mux_h I__13486 (
            .O(N__56466),
            .I(N__56445));
    LocalMux I__13485 (
            .O(N__56463),
            .I(N__56442));
    InMux I__13484 (
            .O(N__56462),
            .I(N__56439));
    InMux I__13483 (
            .O(N__56461),
            .I(N__56434));
    InMux I__13482 (
            .O(N__56460),
            .I(N__56434));
    InMux I__13481 (
            .O(N__56459),
            .I(N__56429));
    InMux I__13480 (
            .O(N__56458),
            .I(N__56429));
    LocalMux I__13479 (
            .O(N__56455),
            .I(N__56426));
    Span4Mux_v I__13478 (
            .O(N__56452),
            .I(N__56423));
    InMux I__13477 (
            .O(N__56451),
            .I(N__56420));
    LocalMux I__13476 (
            .O(N__56448),
            .I(N__56417));
    Span4Mux_v I__13475 (
            .O(N__56445),
            .I(N__56414));
    Sp12to4 I__13474 (
            .O(N__56442),
            .I(N__56405));
    LocalMux I__13473 (
            .O(N__56439),
            .I(N__56405));
    LocalMux I__13472 (
            .O(N__56434),
            .I(N__56405));
    LocalMux I__13471 (
            .O(N__56429),
            .I(N__56405));
    Span4Mux_v I__13470 (
            .O(N__56426),
            .I(N__56396));
    Span4Mux_h I__13469 (
            .O(N__56423),
            .I(N__56396));
    LocalMux I__13468 (
            .O(N__56420),
            .I(N__56396));
    Span4Mux_h I__13467 (
            .O(N__56417),
            .I(N__56396));
    Odrv4 I__13466 (
            .O(N__56414),
            .I(n9324));
    Odrv12 I__13465 (
            .O(N__56405),
            .I(n9324));
    Odrv4 I__13464 (
            .O(N__56396),
            .I(n9324));
    InMux I__13463 (
            .O(N__56389),
            .I(N__56386));
    LocalMux I__13462 (
            .O(N__56386),
            .I(n8_adj_1623));
    CascadeMux I__13461 (
            .O(N__56383),
            .I(n8_adj_1623_cascade_));
    CascadeMux I__13460 (
            .O(N__56380),
            .I(N__56377));
    InMux I__13459 (
            .O(N__56377),
            .I(N__56373));
    InMux I__13458 (
            .O(N__56376),
            .I(N__56370));
    LocalMux I__13457 (
            .O(N__56373),
            .I(N__56365));
    LocalMux I__13456 (
            .O(N__56370),
            .I(N__56365));
    Odrv12 I__13455 (
            .O(N__56365),
            .I(n7_adj_1622));
    CascadeMux I__13454 (
            .O(N__56362),
            .I(N__56359));
    CascadeBuf I__13453 (
            .O(N__56359),
            .I(N__56356));
    CascadeMux I__13452 (
            .O(N__56356),
            .I(N__56353));
    CascadeBuf I__13451 (
            .O(N__56353),
            .I(N__56350));
    CascadeMux I__13450 (
            .O(N__56350),
            .I(N__56347));
    CascadeBuf I__13449 (
            .O(N__56347),
            .I(N__56344));
    CascadeMux I__13448 (
            .O(N__56344),
            .I(N__56341));
    CascadeBuf I__13447 (
            .O(N__56341),
            .I(N__56338));
    CascadeMux I__13446 (
            .O(N__56338),
            .I(N__56335));
    CascadeBuf I__13445 (
            .O(N__56335),
            .I(N__56332));
    CascadeMux I__13444 (
            .O(N__56332),
            .I(N__56329));
    CascadeBuf I__13443 (
            .O(N__56329),
            .I(N__56325));
    CascadeMux I__13442 (
            .O(N__56328),
            .I(N__56322));
    CascadeMux I__13441 (
            .O(N__56325),
            .I(N__56319));
    CascadeBuf I__13440 (
            .O(N__56322),
            .I(N__56316));
    CascadeBuf I__13439 (
            .O(N__56319),
            .I(N__56313));
    CascadeMux I__13438 (
            .O(N__56316),
            .I(N__56310));
    CascadeMux I__13437 (
            .O(N__56313),
            .I(N__56307));
    InMux I__13436 (
            .O(N__56310),
            .I(N__56304));
    CascadeBuf I__13435 (
            .O(N__56307),
            .I(N__56301));
    LocalMux I__13434 (
            .O(N__56304),
            .I(N__56298));
    CascadeMux I__13433 (
            .O(N__56301),
            .I(N__56295));
    Span4Mux_h I__13432 (
            .O(N__56298),
            .I(N__56292));
    CascadeBuf I__13431 (
            .O(N__56295),
            .I(N__56289));
    Span4Mux_v I__13430 (
            .O(N__56292),
            .I(N__56286));
    CascadeMux I__13429 (
            .O(N__56289),
            .I(N__56283));
    Span4Mux_v I__13428 (
            .O(N__56286),
            .I(N__56280));
    InMux I__13427 (
            .O(N__56283),
            .I(N__56277));
    Span4Mux_h I__13426 (
            .O(N__56280),
            .I(N__56274));
    LocalMux I__13425 (
            .O(N__56277),
            .I(N__56271));
    Span4Mux_h I__13424 (
            .O(N__56274),
            .I(N__56268));
    Span4Mux_h I__13423 (
            .O(N__56271),
            .I(N__56265));
    Span4Mux_h I__13422 (
            .O(N__56268),
            .I(N__56260));
    Span4Mux_v I__13421 (
            .O(N__56265),
            .I(N__56260));
    Odrv4 I__13420 (
            .O(N__56260),
            .I(data_index_9_N_236_5));
    InMux I__13419 (
            .O(N__56257),
            .I(N__56254));
    LocalMux I__13418 (
            .O(N__56254),
            .I(N__56251));
    Span4Mux_h I__13417 (
            .O(N__56251),
            .I(N__56248));
    Span4Mux_v I__13416 (
            .O(N__56248),
            .I(N__56244));
    InMux I__13415 (
            .O(N__56247),
            .I(N__56241));
    Odrv4 I__13414 (
            .O(N__56244),
            .I(n21966));
    LocalMux I__13413 (
            .O(N__56241),
            .I(n21966));
    CascadeMux I__13412 (
            .O(N__56236),
            .I(N__56233));
    InMux I__13411 (
            .O(N__56233),
            .I(N__56229));
    CascadeMux I__13410 (
            .O(N__56232),
            .I(N__56225));
    LocalMux I__13409 (
            .O(N__56229),
            .I(N__56222));
    InMux I__13408 (
            .O(N__56228),
            .I(N__56217));
    InMux I__13407 (
            .O(N__56225),
            .I(N__56217));
    Span4Mux_v I__13406 (
            .O(N__56222),
            .I(N__56212));
    LocalMux I__13405 (
            .O(N__56217),
            .I(N__56212));
    Span4Mux_v I__13404 (
            .O(N__56212),
            .I(N__56209));
    Span4Mux_h I__13403 (
            .O(N__56209),
            .I(N__56206));
    Sp12to4 I__13402 (
            .O(N__56206),
            .I(N__56202));
    CascadeMux I__13401 (
            .O(N__56205),
            .I(N__56199));
    Span12Mux_h I__13400 (
            .O(N__56202),
            .I(N__56196));
    InMux I__13399 (
            .O(N__56199),
            .I(N__56193));
    Span12Mux_v I__13398 (
            .O(N__56196),
            .I(N__56190));
    LocalMux I__13397 (
            .O(N__56193),
            .I(trig_dds1));
    Odrv12 I__13396 (
            .O(N__56190),
            .I(trig_dds1));
    InMux I__13395 (
            .O(N__56185),
            .I(N__56181));
    InMux I__13394 (
            .O(N__56184),
            .I(N__56178));
    LocalMux I__13393 (
            .O(N__56181),
            .I(n21920));
    LocalMux I__13392 (
            .O(N__56178),
            .I(n21920));
    CascadeMux I__13391 (
            .O(N__56173),
            .I(n22399_cascade_));
    InMux I__13390 (
            .O(N__56170),
            .I(N__56167));
    LocalMux I__13389 (
            .O(N__56167),
            .I(N__56164));
    Span4Mux_h I__13388 (
            .O(N__56164),
            .I(N__56161));
    Odrv4 I__13387 (
            .O(N__56161),
            .I(n40_adj_1689));
    InMux I__13386 (
            .O(N__56158),
            .I(N__56154));
    CascadeMux I__13385 (
            .O(N__56157),
            .I(N__56151));
    LocalMux I__13384 (
            .O(N__56154),
            .I(N__56148));
    InMux I__13383 (
            .O(N__56151),
            .I(N__56145));
    Span4Mux_h I__13382 (
            .O(N__56148),
            .I(N__56142));
    LocalMux I__13381 (
            .O(N__56145),
            .I(data_idxvec_11));
    Odrv4 I__13380 (
            .O(N__56142),
            .I(data_idxvec_11));
    InMux I__13379 (
            .O(N__56137),
            .I(N__56134));
    LocalMux I__13378 (
            .O(N__56134),
            .I(N__56129));
    InMux I__13377 (
            .O(N__56133),
            .I(N__56126));
    InMux I__13376 (
            .O(N__56132),
            .I(N__56123));
    Span4Mux_v I__13375 (
            .O(N__56129),
            .I(N__56120));
    LocalMux I__13374 (
            .O(N__56126),
            .I(N__56117));
    LocalMux I__13373 (
            .O(N__56123),
            .I(data_cntvec_11));
    Odrv4 I__13372 (
            .O(N__56120),
            .I(data_cntvec_11));
    Odrv4 I__13371 (
            .O(N__56117),
            .I(data_cntvec_11));
    InMux I__13370 (
            .O(N__56110),
            .I(N__56106));
    CascadeMux I__13369 (
            .O(N__56109),
            .I(N__56103));
    LocalMux I__13368 (
            .O(N__56106),
            .I(N__56100));
    InMux I__13367 (
            .O(N__56103),
            .I(N__56097));
    Span4Mux_v I__13366 (
            .O(N__56100),
            .I(N__56093));
    LocalMux I__13365 (
            .O(N__56097),
            .I(N__56090));
    InMux I__13364 (
            .O(N__56096),
            .I(N__56087));
    Span4Mux_h I__13363 (
            .O(N__56093),
            .I(N__56079));
    Span4Mux_v I__13362 (
            .O(N__56090),
            .I(N__56079));
    LocalMux I__13361 (
            .O(N__56087),
            .I(N__56079));
    CascadeMux I__13360 (
            .O(N__56086),
            .I(N__56075));
    Span4Mux_h I__13359 (
            .O(N__56079),
            .I(N__56071));
    CascadeMux I__13358 (
            .O(N__56078),
            .I(N__56066));
    InMux I__13357 (
            .O(N__56075),
            .I(N__56062));
    InMux I__13356 (
            .O(N__56074),
            .I(N__56059));
    Span4Mux_h I__13355 (
            .O(N__56071),
            .I(N__56056));
    InMux I__13354 (
            .O(N__56070),
            .I(N__56051));
    InMux I__13353 (
            .O(N__56069),
            .I(N__56051));
    InMux I__13352 (
            .O(N__56066),
            .I(N__56048));
    InMux I__13351 (
            .O(N__56065),
            .I(N__56045));
    LocalMux I__13350 (
            .O(N__56062),
            .I(N__56042));
    LocalMux I__13349 (
            .O(N__56059),
            .I(N__56037));
    Span4Mux_v I__13348 (
            .O(N__56056),
            .I(N__56037));
    LocalMux I__13347 (
            .O(N__56051),
            .I(N__56030));
    LocalMux I__13346 (
            .O(N__56048),
            .I(N__56030));
    LocalMux I__13345 (
            .O(N__56045),
            .I(N__56030));
    Odrv4 I__13344 (
            .O(N__56042),
            .I(comm_buf_1_4));
    Odrv4 I__13343 (
            .O(N__56037),
            .I(comm_buf_1_4));
    Odrv12 I__13342 (
            .O(N__56030),
            .I(comm_buf_1_4));
    InMux I__13341 (
            .O(N__56023),
            .I(N__56019));
    InMux I__13340 (
            .O(N__56022),
            .I(N__56016));
    LocalMux I__13339 (
            .O(N__56019),
            .I(N__56013));
    LocalMux I__13338 (
            .O(N__56016),
            .I(N__56010));
    Span4Mux_h I__13337 (
            .O(N__56013),
            .I(N__56007));
    Span4Mux_h I__13336 (
            .O(N__56010),
            .I(N__56004));
    Odrv4 I__13335 (
            .O(N__56007),
            .I(n14_adj_1611));
    Odrv4 I__13334 (
            .O(N__56004),
            .I(n14_adj_1611));
    InMux I__13333 (
            .O(N__55999),
            .I(N__55996));
    LocalMux I__13332 (
            .O(N__55996),
            .I(N__55993));
    Span4Mux_v I__13331 (
            .O(N__55993),
            .I(N__55990));
    Sp12to4 I__13330 (
            .O(N__55990),
            .I(N__55987));
    Span12Mux_h I__13329 (
            .O(N__55987),
            .I(N__55984));
    Odrv12 I__13328 (
            .O(N__55984),
            .I(n22272));
    CascadeMux I__13327 (
            .O(N__55981),
            .I(n23420_cascade_));
    InMux I__13326 (
            .O(N__55978),
            .I(N__55975));
    LocalMux I__13325 (
            .O(N__55975),
            .I(N__55972));
    Span4Mux_h I__13324 (
            .O(N__55972),
            .I(N__55969));
    Odrv4 I__13323 (
            .O(N__55969),
            .I(n22271));
    InMux I__13322 (
            .O(N__55966),
            .I(N__55963));
    LocalMux I__13321 (
            .O(N__55963),
            .I(N__55960));
    Span4Mux_v I__13320 (
            .O(N__55960),
            .I(N__55957));
    Span4Mux_v I__13319 (
            .O(N__55957),
            .I(N__55954));
    Sp12to4 I__13318 (
            .O(N__55954),
            .I(N__55951));
    Odrv12 I__13317 (
            .O(N__55951),
            .I(n111_adj_1719));
    CascadeMux I__13316 (
            .O(N__55948),
            .I(n23423_cascade_));
    CascadeMux I__13315 (
            .O(N__55945),
            .I(N__55942));
    InMux I__13314 (
            .O(N__55942),
            .I(N__55938));
    CascadeMux I__13313 (
            .O(N__55941),
            .I(N__55932));
    LocalMux I__13312 (
            .O(N__55938),
            .I(N__55928));
    InMux I__13311 (
            .O(N__55937),
            .I(N__55925));
    CascadeMux I__13310 (
            .O(N__55936),
            .I(N__55922));
    InMux I__13309 (
            .O(N__55935),
            .I(N__55917));
    InMux I__13308 (
            .O(N__55932),
            .I(N__55917));
    CascadeMux I__13307 (
            .O(N__55931),
            .I(N__55914));
    Span4Mux_v I__13306 (
            .O(N__55928),
            .I(N__55909));
    LocalMux I__13305 (
            .O(N__55925),
            .I(N__55909));
    InMux I__13304 (
            .O(N__55922),
            .I(N__55906));
    LocalMux I__13303 (
            .O(N__55917),
            .I(N__55903));
    InMux I__13302 (
            .O(N__55914),
            .I(N__55900));
    Span4Mux_v I__13301 (
            .O(N__55909),
            .I(N__55896));
    LocalMux I__13300 (
            .O(N__55906),
            .I(N__55893));
    Span4Mux_v I__13299 (
            .O(N__55903),
            .I(N__55888));
    LocalMux I__13298 (
            .O(N__55900),
            .I(N__55888));
    InMux I__13297 (
            .O(N__55899),
            .I(N__55885));
    Span4Mux_h I__13296 (
            .O(N__55896),
            .I(N__55881));
    Span4Mux_v I__13295 (
            .O(N__55893),
            .I(N__55878));
    Span4Mux_h I__13294 (
            .O(N__55888),
            .I(N__55873));
    LocalMux I__13293 (
            .O(N__55885),
            .I(N__55873));
    InMux I__13292 (
            .O(N__55884),
            .I(N__55870));
    Span4Mux_h I__13291 (
            .O(N__55881),
            .I(N__55867));
    Span4Mux_h I__13290 (
            .O(N__55878),
            .I(N__55862));
    Span4Mux_v I__13289 (
            .O(N__55873),
            .I(N__55862));
    LocalMux I__13288 (
            .O(N__55870),
            .I(N__55859));
    Odrv4 I__13287 (
            .O(N__55867),
            .I(comm_rx_buf_7));
    Odrv4 I__13286 (
            .O(N__55862),
            .I(comm_rx_buf_7));
    Odrv4 I__13285 (
            .O(N__55859),
            .I(comm_rx_buf_7));
    CascadeMux I__13284 (
            .O(N__55852),
            .I(comm_buf_1_7_N_559_7_cascade_));
    CascadeMux I__13283 (
            .O(N__55849),
            .I(N__55845));
    InMux I__13282 (
            .O(N__55848),
            .I(N__55842));
    InMux I__13281 (
            .O(N__55845),
            .I(N__55838));
    LocalMux I__13280 (
            .O(N__55842),
            .I(N__55834));
    InMux I__13279 (
            .O(N__55841),
            .I(N__55831));
    LocalMux I__13278 (
            .O(N__55838),
            .I(N__55828));
    CascadeMux I__13277 (
            .O(N__55837),
            .I(N__55824));
    Span4Mux_v I__13276 (
            .O(N__55834),
            .I(N__55817));
    LocalMux I__13275 (
            .O(N__55831),
            .I(N__55817));
    Sp12to4 I__13274 (
            .O(N__55828),
            .I(N__55814));
    InMux I__13273 (
            .O(N__55827),
            .I(N__55811));
    InMux I__13272 (
            .O(N__55824),
            .I(N__55808));
    InMux I__13271 (
            .O(N__55823),
            .I(N__55805));
    InMux I__13270 (
            .O(N__55822),
            .I(N__55802));
    Span4Mux_h I__13269 (
            .O(N__55817),
            .I(N__55799));
    Span12Mux_v I__13268 (
            .O(N__55814),
            .I(N__55792));
    LocalMux I__13267 (
            .O(N__55811),
            .I(N__55792));
    LocalMux I__13266 (
            .O(N__55808),
            .I(N__55792));
    LocalMux I__13265 (
            .O(N__55805),
            .I(N__55787));
    LocalMux I__13264 (
            .O(N__55802),
            .I(N__55787));
    Span4Mux_h I__13263 (
            .O(N__55799),
            .I(N__55784));
    Span12Mux_h I__13262 (
            .O(N__55792),
            .I(N__55781));
    Odrv12 I__13261 (
            .O(N__55787),
            .I(comm_buf_1_7));
    Odrv4 I__13260 (
            .O(N__55784),
            .I(comm_buf_1_7));
    Odrv12 I__13259 (
            .O(N__55781),
            .I(comm_buf_1_7));
    CEMux I__13258 (
            .O(N__55774),
            .I(N__55771));
    LocalMux I__13257 (
            .O(N__55771),
            .I(N__55764));
    CEMux I__13256 (
            .O(N__55770),
            .I(N__55761));
    CEMux I__13255 (
            .O(N__55769),
            .I(N__55758));
    CEMux I__13254 (
            .O(N__55768),
            .I(N__55755));
    CEMux I__13253 (
            .O(N__55767),
            .I(N__55752));
    Span4Mux_v I__13252 (
            .O(N__55764),
            .I(N__55746));
    LocalMux I__13251 (
            .O(N__55761),
            .I(N__55746));
    LocalMux I__13250 (
            .O(N__55758),
            .I(N__55743));
    LocalMux I__13249 (
            .O(N__55755),
            .I(N__55740));
    LocalMux I__13248 (
            .O(N__55752),
            .I(N__55737));
    CEMux I__13247 (
            .O(N__55751),
            .I(N__55734));
    Span4Mux_h I__13246 (
            .O(N__55746),
            .I(N__55729));
    Span4Mux_h I__13245 (
            .O(N__55743),
            .I(N__55729));
    Span4Mux_v I__13244 (
            .O(N__55740),
            .I(N__55724));
    Span4Mux_h I__13243 (
            .O(N__55737),
            .I(N__55724));
    LocalMux I__13242 (
            .O(N__55734),
            .I(N__55721));
    Odrv4 I__13241 (
            .O(N__55729),
            .I(n12761));
    Odrv4 I__13240 (
            .O(N__55724),
            .I(n12761));
    Odrv12 I__13239 (
            .O(N__55721),
            .I(n12761));
    SRMux I__13238 (
            .O(N__55714),
            .I(N__55711));
    LocalMux I__13237 (
            .O(N__55711),
            .I(N__55704));
    SRMux I__13236 (
            .O(N__55710),
            .I(N__55701));
    SRMux I__13235 (
            .O(N__55709),
            .I(N__55697));
    SRMux I__13234 (
            .O(N__55708),
            .I(N__55694));
    SRMux I__13233 (
            .O(N__55707),
            .I(N__55691));
    Span4Mux_h I__13232 (
            .O(N__55704),
            .I(N__55686));
    LocalMux I__13231 (
            .O(N__55701),
            .I(N__55686));
    SRMux I__13230 (
            .O(N__55700),
            .I(N__55683));
    LocalMux I__13229 (
            .O(N__55697),
            .I(N__55678));
    LocalMux I__13228 (
            .O(N__55694),
            .I(N__55678));
    LocalMux I__13227 (
            .O(N__55691),
            .I(N__55675));
    Span4Mux_h I__13226 (
            .O(N__55686),
            .I(N__55670));
    LocalMux I__13225 (
            .O(N__55683),
            .I(N__55670));
    Span4Mux_v I__13224 (
            .O(N__55678),
            .I(N__55667));
    Span4Mux_h I__13223 (
            .O(N__55675),
            .I(N__55664));
    Span4Mux_v I__13222 (
            .O(N__55670),
            .I(N__55661));
    Span4Mux_h I__13221 (
            .O(N__55667),
            .I(N__55658));
    Odrv4 I__13220 (
            .O(N__55664),
            .I(n15489));
    Odrv4 I__13219 (
            .O(N__55661),
            .I(n15489));
    Odrv4 I__13218 (
            .O(N__55658),
            .I(n15489));
    CascadeMux I__13217 (
            .O(N__55651),
            .I(N__55646));
    InMux I__13216 (
            .O(N__55650),
            .I(N__55641));
    InMux I__13215 (
            .O(N__55649),
            .I(N__55641));
    InMux I__13214 (
            .O(N__55646),
            .I(N__55637));
    LocalMux I__13213 (
            .O(N__55641),
            .I(N__55631));
    InMux I__13212 (
            .O(N__55640),
            .I(N__55627));
    LocalMux I__13211 (
            .O(N__55637),
            .I(N__55623));
    InMux I__13210 (
            .O(N__55636),
            .I(N__55616));
    InMux I__13209 (
            .O(N__55635),
            .I(N__55616));
    InMux I__13208 (
            .O(N__55634),
            .I(N__55616));
    Span4Mux_h I__13207 (
            .O(N__55631),
            .I(N__55613));
    InMux I__13206 (
            .O(N__55630),
            .I(N__55610));
    LocalMux I__13205 (
            .O(N__55627),
            .I(N__55607));
    InMux I__13204 (
            .O(N__55626),
            .I(N__55604));
    Span4Mux_v I__13203 (
            .O(N__55623),
            .I(N__55599));
    LocalMux I__13202 (
            .O(N__55616),
            .I(N__55599));
    Span4Mux_h I__13201 (
            .O(N__55613),
            .I(N__55595));
    LocalMux I__13200 (
            .O(N__55610),
            .I(N__55592));
    Span4Mux_h I__13199 (
            .O(N__55607),
            .I(N__55589));
    LocalMux I__13198 (
            .O(N__55604),
            .I(N__55584));
    Sp12to4 I__13197 (
            .O(N__55599),
            .I(N__55584));
    InMux I__13196 (
            .O(N__55598),
            .I(N__55581));
    Span4Mux_v I__13195 (
            .O(N__55595),
            .I(N__55576));
    Span4Mux_v I__13194 (
            .O(N__55592),
            .I(N__55576));
    Span4Mux_v I__13193 (
            .O(N__55589),
            .I(N__55573));
    Span12Mux_v I__13192 (
            .O(N__55584),
            .I(N__55570));
    LocalMux I__13191 (
            .O(N__55581),
            .I(N__55565));
    Span4Mux_h I__13190 (
            .O(N__55576),
            .I(N__55565));
    Odrv4 I__13189 (
            .O(N__55573),
            .I(n18955));
    Odrv12 I__13188 (
            .O(N__55570),
            .I(n18955));
    Odrv4 I__13187 (
            .O(N__55565),
            .I(n18955));
    InMux I__13186 (
            .O(N__55558),
            .I(N__55555));
    LocalMux I__13185 (
            .O(N__55555),
            .I(N__55552));
    Odrv4 I__13184 (
            .O(N__55552),
            .I(n22356));
    InMux I__13183 (
            .O(N__55549),
            .I(N__55545));
    CascadeMux I__13182 (
            .O(N__55548),
            .I(N__55542));
    LocalMux I__13181 (
            .O(N__55545),
            .I(N__55539));
    InMux I__13180 (
            .O(N__55542),
            .I(N__55536));
    Span4Mux_v I__13179 (
            .O(N__55539),
            .I(N__55533));
    LocalMux I__13178 (
            .O(N__55536),
            .I(N__55530));
    Span4Mux_h I__13177 (
            .O(N__55533),
            .I(N__55526));
    Span4Mux_v I__13176 (
            .O(N__55530),
            .I(N__55523));
    InMux I__13175 (
            .O(N__55529),
            .I(N__55520));
    Span4Mux_v I__13174 (
            .O(N__55526),
            .I(N__55515));
    Span4Mux_h I__13173 (
            .O(N__55523),
            .I(N__55515));
    LocalMux I__13172 (
            .O(N__55520),
            .I(buf_dds0_13));
    Odrv4 I__13171 (
            .O(N__55515),
            .I(buf_dds0_13));
    InMux I__13170 (
            .O(N__55510),
            .I(N__55507));
    LocalMux I__13169 (
            .O(N__55507),
            .I(N__55504));
    Odrv12 I__13168 (
            .O(N__55504),
            .I(n23348));
    InMux I__13167 (
            .O(N__55501),
            .I(N__55498));
    LocalMux I__13166 (
            .O(N__55498),
            .I(N__55494));
    CascadeMux I__13165 (
            .O(N__55497),
            .I(N__55491));
    Span4Mux_h I__13164 (
            .O(N__55494),
            .I(N__55487));
    InMux I__13163 (
            .O(N__55491),
            .I(N__55482));
    InMux I__13162 (
            .O(N__55490),
            .I(N__55482));
    Odrv4 I__13161 (
            .O(N__55487),
            .I(req_data_cnt_7));
    LocalMux I__13160 (
            .O(N__55482),
            .I(req_data_cnt_7));
    InMux I__13159 (
            .O(N__55477),
            .I(N__55474));
    LocalMux I__13158 (
            .O(N__55474),
            .I(N__55471));
    Span12Mux_v I__13157 (
            .O(N__55471),
            .I(N__55466));
    InMux I__13156 (
            .O(N__55470),
            .I(N__55461));
    InMux I__13155 (
            .O(N__55469),
            .I(N__55461));
    Odrv12 I__13154 (
            .O(N__55466),
            .I(acadc_skipCount_7));
    LocalMux I__13153 (
            .O(N__55461),
            .I(acadc_skipCount_7));
    InMux I__13152 (
            .O(N__55456),
            .I(N__55453));
    LocalMux I__13151 (
            .O(N__55453),
            .I(n22262));
    InMux I__13150 (
            .O(N__55450),
            .I(N__55447));
    LocalMux I__13149 (
            .O(N__55447),
            .I(N__55444));
    Odrv12 I__13148 (
            .O(N__55444),
            .I(buf_data_iac_14));
    InMux I__13147 (
            .O(N__55441),
            .I(N__55438));
    LocalMux I__13146 (
            .O(N__55438),
            .I(N__55435));
    Odrv4 I__13145 (
            .O(N__55435),
            .I(n22391));
    InMux I__13144 (
            .O(N__55432),
            .I(N__55427));
    InMux I__13143 (
            .O(N__55431),
            .I(N__55424));
    InMux I__13142 (
            .O(N__55430),
            .I(N__55420));
    LocalMux I__13141 (
            .O(N__55427),
            .I(N__55415));
    LocalMux I__13140 (
            .O(N__55424),
            .I(N__55415));
    InMux I__13139 (
            .O(N__55423),
            .I(N__55412));
    LocalMux I__13138 (
            .O(N__55420),
            .I(N__55409));
    Span4Mux_v I__13137 (
            .O(N__55415),
            .I(N__55404));
    LocalMux I__13136 (
            .O(N__55412),
            .I(N__55404));
    Span4Mux_v I__13135 (
            .O(N__55409),
            .I(N__55394));
    Span4Mux_v I__13134 (
            .O(N__55404),
            .I(N__55394));
    InMux I__13133 (
            .O(N__55403),
            .I(N__55389));
    InMux I__13132 (
            .O(N__55402),
            .I(N__55389));
    InMux I__13131 (
            .O(N__55401),
            .I(N__55385));
    CascadeMux I__13130 (
            .O(N__55400),
            .I(N__55382));
    InMux I__13129 (
            .O(N__55399),
            .I(N__55377));
    Span4Mux_h I__13128 (
            .O(N__55394),
            .I(N__55372));
    LocalMux I__13127 (
            .O(N__55389),
            .I(N__55372));
    InMux I__13126 (
            .O(N__55388),
            .I(N__55365));
    LocalMux I__13125 (
            .O(N__55385),
            .I(N__55362));
    InMux I__13124 (
            .O(N__55382),
            .I(N__55359));
    InMux I__13123 (
            .O(N__55381),
            .I(N__55356));
    InMux I__13122 (
            .O(N__55380),
            .I(N__55353));
    LocalMux I__13121 (
            .O(N__55377),
            .I(N__55348));
    Span4Mux_v I__13120 (
            .O(N__55372),
            .I(N__55348));
    InMux I__13119 (
            .O(N__55371),
            .I(N__55345));
    InMux I__13118 (
            .O(N__55370),
            .I(N__55338));
    InMux I__13117 (
            .O(N__55369),
            .I(N__55338));
    InMux I__13116 (
            .O(N__55368),
            .I(N__55338));
    LocalMux I__13115 (
            .O(N__55365),
            .I(N__55335));
    Span4Mux_h I__13114 (
            .O(N__55362),
            .I(N__55332));
    LocalMux I__13113 (
            .O(N__55359),
            .I(N__55329));
    LocalMux I__13112 (
            .O(N__55356),
            .I(N__55326));
    LocalMux I__13111 (
            .O(N__55353),
            .I(N__55323));
    Span4Mux_h I__13110 (
            .O(N__55348),
            .I(N__55320));
    LocalMux I__13109 (
            .O(N__55345),
            .I(N__55313));
    LocalMux I__13108 (
            .O(N__55338),
            .I(N__55313));
    Sp12to4 I__13107 (
            .O(N__55335),
            .I(N__55313));
    Span4Mux_h I__13106 (
            .O(N__55332),
            .I(N__55310));
    Span12Mux_h I__13105 (
            .O(N__55329),
            .I(N__55307));
    Span4Mux_v I__13104 (
            .O(N__55326),
            .I(N__55304));
    Span12Mux_v I__13103 (
            .O(N__55323),
            .I(N__55297));
    Sp12to4 I__13102 (
            .O(N__55320),
            .I(N__55297));
    Span12Mux_v I__13101 (
            .O(N__55313),
            .I(N__55297));
    Odrv4 I__13100 (
            .O(N__55310),
            .I(n12509));
    Odrv12 I__13099 (
            .O(N__55307),
            .I(n12509));
    Odrv4 I__13098 (
            .O(N__55304),
            .I(n12509));
    Odrv12 I__13097 (
            .O(N__55297),
            .I(n12509));
    InMux I__13096 (
            .O(N__55288),
            .I(N__55284));
    InMux I__13095 (
            .O(N__55287),
            .I(N__55280));
    LocalMux I__13094 (
            .O(N__55284),
            .I(N__55277));
    CascadeMux I__13093 (
            .O(N__55283),
            .I(N__55273));
    LocalMux I__13092 (
            .O(N__55280),
            .I(N__55270));
    Sp12to4 I__13091 (
            .O(N__55277),
            .I(N__55267));
    InMux I__13090 (
            .O(N__55276),
            .I(N__55264));
    InMux I__13089 (
            .O(N__55273),
            .I(N__55261));
    Span4Mux_v I__13088 (
            .O(N__55270),
            .I(N__55258));
    Span12Mux_v I__13087 (
            .O(N__55267),
            .I(N__55255));
    LocalMux I__13086 (
            .O(N__55264),
            .I(N__55252));
    LocalMux I__13085 (
            .O(N__55261),
            .I(N__55249));
    Span4Mux_h I__13084 (
            .O(N__55258),
            .I(N__55246));
    Odrv12 I__13083 (
            .O(N__55255),
            .I(n14_adj_1660));
    Odrv4 I__13082 (
            .O(N__55252),
            .I(n14_adj_1660));
    Odrv4 I__13081 (
            .O(N__55249),
            .I(n14_adj_1660));
    Odrv4 I__13080 (
            .O(N__55246),
            .I(n14_adj_1660));
    InMux I__13079 (
            .O(N__55237),
            .I(N__55234));
    LocalMux I__13078 (
            .O(N__55234),
            .I(N__55231));
    Span4Mux_v I__13077 (
            .O(N__55231),
            .I(N__55228));
    Sp12to4 I__13076 (
            .O(N__55228),
            .I(N__55224));
    InMux I__13075 (
            .O(N__55227),
            .I(N__55220));
    Span12Mux_h I__13074 (
            .O(N__55224),
            .I(N__55217));
    InMux I__13073 (
            .O(N__55223),
            .I(N__55214));
    LocalMux I__13072 (
            .O(N__55220),
            .I(buf_dds1_13));
    Odrv12 I__13071 (
            .O(N__55217),
            .I(buf_dds1_13));
    LocalMux I__13070 (
            .O(N__55214),
            .I(buf_dds1_13));
    InMux I__13069 (
            .O(N__55207),
            .I(N__55203));
    InMux I__13068 (
            .O(N__55206),
            .I(N__55200));
    LocalMux I__13067 (
            .O(N__55203),
            .I(N__55195));
    LocalMux I__13066 (
            .O(N__55200),
            .I(N__55195));
    Span4Mux_v I__13065 (
            .O(N__55195),
            .I(N__55190));
    CascadeMux I__13064 (
            .O(N__55194),
            .I(N__55186));
    CascadeMux I__13063 (
            .O(N__55193),
            .I(N__55183));
    Span4Mux_h I__13062 (
            .O(N__55190),
            .I(N__55180));
    InMux I__13061 (
            .O(N__55189),
            .I(N__55177));
    InMux I__13060 (
            .O(N__55186),
            .I(N__55174));
    InMux I__13059 (
            .O(N__55183),
            .I(N__55171));
    Span4Mux_v I__13058 (
            .O(N__55180),
            .I(N__55164));
    LocalMux I__13057 (
            .O(N__55177),
            .I(N__55164));
    LocalMux I__13056 (
            .O(N__55174),
            .I(N__55161));
    LocalMux I__13055 (
            .O(N__55171),
            .I(N__55157));
    InMux I__13054 (
            .O(N__55170),
            .I(N__55154));
    CascadeMux I__13053 (
            .O(N__55169),
            .I(N__55151));
    Span4Mux_v I__13052 (
            .O(N__55164),
            .I(N__55148));
    Span4Mux_v I__13051 (
            .O(N__55161),
            .I(N__55145));
    InMux I__13050 (
            .O(N__55160),
            .I(N__55142));
    Span4Mux_v I__13049 (
            .O(N__55157),
            .I(N__55139));
    LocalMux I__13048 (
            .O(N__55154),
            .I(N__55136));
    InMux I__13047 (
            .O(N__55151),
            .I(N__55133));
    Span4Mux_h I__13046 (
            .O(N__55148),
            .I(N__55129));
    Sp12to4 I__13045 (
            .O(N__55145),
            .I(N__55124));
    LocalMux I__13044 (
            .O(N__55142),
            .I(N__55124));
    Span4Mux_h I__13043 (
            .O(N__55139),
            .I(N__55117));
    Span4Mux_h I__13042 (
            .O(N__55136),
            .I(N__55117));
    LocalMux I__13041 (
            .O(N__55133),
            .I(N__55117));
    InMux I__13040 (
            .O(N__55132),
            .I(N__55114));
    Odrv4 I__13039 (
            .O(N__55129),
            .I(comm_rx_buf_5));
    Odrv12 I__13038 (
            .O(N__55124),
            .I(comm_rx_buf_5));
    Odrv4 I__13037 (
            .O(N__55117),
            .I(comm_rx_buf_5));
    LocalMux I__13036 (
            .O(N__55114),
            .I(comm_rx_buf_5));
    InMux I__13035 (
            .O(N__55105),
            .I(N__55102));
    LocalMux I__13034 (
            .O(N__55102),
            .I(N__55099));
    Span4Mux_h I__13033 (
            .O(N__55099),
            .I(N__55096));
    Odrv4 I__13032 (
            .O(N__55096),
            .I(buf_data_vac_13));
    InMux I__13031 (
            .O(N__55093),
            .I(N__55090));
    LocalMux I__13030 (
            .O(N__55090),
            .I(N__55087));
    Span4Mux_h I__13029 (
            .O(N__55087),
            .I(N__55084));
    Odrv4 I__13028 (
            .O(N__55084),
            .I(comm_buf_4_5));
    CascadeMux I__13027 (
            .O(N__55081),
            .I(N__55078));
    InMux I__13026 (
            .O(N__55078),
            .I(N__55073));
    InMux I__13025 (
            .O(N__55077),
            .I(N__55068));
    CascadeMux I__13024 (
            .O(N__55076),
            .I(N__55064));
    LocalMux I__13023 (
            .O(N__55073),
            .I(N__55061));
    InMux I__13022 (
            .O(N__55072),
            .I(N__55057));
    InMux I__13021 (
            .O(N__55071),
            .I(N__55054));
    LocalMux I__13020 (
            .O(N__55068),
            .I(N__55051));
    InMux I__13019 (
            .O(N__55067),
            .I(N__55048));
    InMux I__13018 (
            .O(N__55064),
            .I(N__55045));
    Span4Mux_v I__13017 (
            .O(N__55061),
            .I(N__55042));
    InMux I__13016 (
            .O(N__55060),
            .I(N__55039));
    LocalMux I__13015 (
            .O(N__55057),
            .I(N__55033));
    LocalMux I__13014 (
            .O(N__55054),
            .I(N__55033));
    Span4Mux_v I__13013 (
            .O(N__55051),
            .I(N__55028));
    LocalMux I__13012 (
            .O(N__55048),
            .I(N__55028));
    LocalMux I__13011 (
            .O(N__55045),
            .I(N__55025));
    Span4Mux_h I__13010 (
            .O(N__55042),
            .I(N__55020));
    LocalMux I__13009 (
            .O(N__55039),
            .I(N__55020));
    InMux I__13008 (
            .O(N__55038),
            .I(N__55017));
    Span12Mux_v I__13007 (
            .O(N__55033),
            .I(N__55013));
    Span4Mux_h I__13006 (
            .O(N__55028),
            .I(N__55010));
    Span12Mux_h I__13005 (
            .O(N__55025),
            .I(N__55003));
    Sp12to4 I__13004 (
            .O(N__55020),
            .I(N__55003));
    LocalMux I__13003 (
            .O(N__55017),
            .I(N__55003));
    InMux I__13002 (
            .O(N__55016),
            .I(N__55000));
    Odrv12 I__13001 (
            .O(N__55013),
            .I(comm_rx_buf_4));
    Odrv4 I__13000 (
            .O(N__55010),
            .I(comm_rx_buf_4));
    Odrv12 I__12999 (
            .O(N__55003),
            .I(comm_rx_buf_4));
    LocalMux I__12998 (
            .O(N__55000),
            .I(comm_rx_buf_4));
    InMux I__12997 (
            .O(N__54991),
            .I(N__54988));
    LocalMux I__12996 (
            .O(N__54988),
            .I(N__54985));
    Span12Mux_v I__12995 (
            .O(N__54985),
            .I(N__54982));
    Odrv12 I__12994 (
            .O(N__54982),
            .I(buf_data_vac_12));
    InMux I__12993 (
            .O(N__54979),
            .I(N__54976));
    LocalMux I__12992 (
            .O(N__54976),
            .I(N__54973));
    Span4Mux_v I__12991 (
            .O(N__54973),
            .I(N__54970));
    Span4Mux_h I__12990 (
            .O(N__54970),
            .I(N__54967));
    Odrv4 I__12989 (
            .O(N__54967),
            .I(comm_buf_4_4));
    InMux I__12988 (
            .O(N__54964),
            .I(N__54961));
    LocalMux I__12987 (
            .O(N__54961),
            .I(N__54958));
    Span4Mux_h I__12986 (
            .O(N__54958),
            .I(N__54955));
    Span4Mux_v I__12985 (
            .O(N__54955),
            .I(N__54952));
    Odrv4 I__12984 (
            .O(N__54952),
            .I(buf_data_vac_11));
    InMux I__12983 (
            .O(N__54949),
            .I(N__54946));
    LocalMux I__12982 (
            .O(N__54946),
            .I(N__54943));
    Odrv4 I__12981 (
            .O(N__54943),
            .I(comm_buf_4_3));
    InMux I__12980 (
            .O(N__54940),
            .I(N__54935));
    InMux I__12979 (
            .O(N__54939),
            .I(N__54932));
    InMux I__12978 (
            .O(N__54938),
            .I(N__54926));
    LocalMux I__12977 (
            .O(N__54935),
            .I(N__54920));
    LocalMux I__12976 (
            .O(N__54932),
            .I(N__54920));
    InMux I__12975 (
            .O(N__54931),
            .I(N__54917));
    InMux I__12974 (
            .O(N__54930),
            .I(N__54914));
    InMux I__12973 (
            .O(N__54929),
            .I(N__54911));
    LocalMux I__12972 (
            .O(N__54926),
            .I(N__54908));
    InMux I__12971 (
            .O(N__54925),
            .I(N__54905));
    Span4Mux_v I__12970 (
            .O(N__54920),
            .I(N__54900));
    LocalMux I__12969 (
            .O(N__54917),
            .I(N__54900));
    LocalMux I__12968 (
            .O(N__54914),
            .I(N__54897));
    LocalMux I__12967 (
            .O(N__54911),
            .I(N__54893));
    Span4Mux_v I__12966 (
            .O(N__54908),
            .I(N__54888));
    LocalMux I__12965 (
            .O(N__54905),
            .I(N__54888));
    Span4Mux_h I__12964 (
            .O(N__54900),
            .I(N__54885));
    Span4Mux_v I__12963 (
            .O(N__54897),
            .I(N__54882));
    InMux I__12962 (
            .O(N__54896),
            .I(N__54879));
    Span12Mux_v I__12961 (
            .O(N__54893),
            .I(N__54875));
    Span4Mux_h I__12960 (
            .O(N__54888),
            .I(N__54872));
    Span4Mux_v I__12959 (
            .O(N__54885),
            .I(N__54869));
    Span4Mux_h I__12958 (
            .O(N__54882),
            .I(N__54864));
    LocalMux I__12957 (
            .O(N__54879),
            .I(N__54864));
    InMux I__12956 (
            .O(N__54878),
            .I(N__54861));
    Odrv12 I__12955 (
            .O(N__54875),
            .I(comm_rx_buf_2));
    Odrv4 I__12954 (
            .O(N__54872),
            .I(comm_rx_buf_2));
    Odrv4 I__12953 (
            .O(N__54869),
            .I(comm_rx_buf_2));
    Odrv4 I__12952 (
            .O(N__54864),
            .I(comm_rx_buf_2));
    LocalMux I__12951 (
            .O(N__54861),
            .I(comm_rx_buf_2));
    InMux I__12950 (
            .O(N__54850),
            .I(N__54847));
    LocalMux I__12949 (
            .O(N__54847),
            .I(N__54844));
    Span12Mux_v I__12948 (
            .O(N__54844),
            .I(N__54841));
    Odrv12 I__12947 (
            .O(N__54841),
            .I(buf_data_vac_10));
    InMux I__12946 (
            .O(N__54838),
            .I(N__54835));
    LocalMux I__12945 (
            .O(N__54835),
            .I(N__54832));
    Span4Mux_h I__12944 (
            .O(N__54832),
            .I(N__54829));
    Span4Mux_h I__12943 (
            .O(N__54829),
            .I(N__54826));
    Odrv4 I__12942 (
            .O(N__54826),
            .I(comm_buf_4_2));
    CascadeMux I__12941 (
            .O(N__54823),
            .I(N__54820));
    InMux I__12940 (
            .O(N__54820),
            .I(N__54817));
    LocalMux I__12939 (
            .O(N__54817),
            .I(N__54813));
    InMux I__12938 (
            .O(N__54816),
            .I(N__54810));
    Span4Mux_v I__12937 (
            .O(N__54813),
            .I(N__54804));
    LocalMux I__12936 (
            .O(N__54810),
            .I(N__54804));
    InMux I__12935 (
            .O(N__54809),
            .I(N__54801));
    Span4Mux_v I__12934 (
            .O(N__54804),
            .I(N__54797));
    LocalMux I__12933 (
            .O(N__54801),
            .I(N__54793));
    InMux I__12932 (
            .O(N__54800),
            .I(N__54789));
    Span4Mux_h I__12931 (
            .O(N__54797),
            .I(N__54785));
    InMux I__12930 (
            .O(N__54796),
            .I(N__54782));
    Span4Mux_h I__12929 (
            .O(N__54793),
            .I(N__54779));
    InMux I__12928 (
            .O(N__54792),
            .I(N__54776));
    LocalMux I__12927 (
            .O(N__54789),
            .I(N__54773));
    InMux I__12926 (
            .O(N__54788),
            .I(N__54770));
    Span4Mux_h I__12925 (
            .O(N__54785),
            .I(N__54764));
    LocalMux I__12924 (
            .O(N__54782),
            .I(N__54764));
    Span4Mux_v I__12923 (
            .O(N__54779),
            .I(N__54759));
    LocalMux I__12922 (
            .O(N__54776),
            .I(N__54759));
    Span4Mux_v I__12921 (
            .O(N__54773),
            .I(N__54754));
    LocalMux I__12920 (
            .O(N__54770),
            .I(N__54754));
    InMux I__12919 (
            .O(N__54769),
            .I(N__54751));
    Span4Mux_v I__12918 (
            .O(N__54764),
            .I(N__54747));
    Span4Mux_h I__12917 (
            .O(N__54759),
            .I(N__54744));
    Span4Mux_h I__12916 (
            .O(N__54754),
            .I(N__54741));
    LocalMux I__12915 (
            .O(N__54751),
            .I(N__54738));
    InMux I__12914 (
            .O(N__54750),
            .I(N__54735));
    Odrv4 I__12913 (
            .O(N__54747),
            .I(comm_rx_buf_1));
    Odrv4 I__12912 (
            .O(N__54744),
            .I(comm_rx_buf_1));
    Odrv4 I__12911 (
            .O(N__54741),
            .I(comm_rx_buf_1));
    Odrv4 I__12910 (
            .O(N__54738),
            .I(comm_rx_buf_1));
    LocalMux I__12909 (
            .O(N__54735),
            .I(comm_rx_buf_1));
    InMux I__12908 (
            .O(N__54724),
            .I(N__54721));
    LocalMux I__12907 (
            .O(N__54721),
            .I(N__54718));
    Span4Mux_h I__12906 (
            .O(N__54718),
            .I(N__54715));
    Span4Mux_v I__12905 (
            .O(N__54715),
            .I(N__54712));
    Odrv4 I__12904 (
            .O(N__54712),
            .I(buf_data_vac_9));
    InMux I__12903 (
            .O(N__54709),
            .I(N__54706));
    LocalMux I__12902 (
            .O(N__54706),
            .I(N__54703));
    Span4Mux_h I__12901 (
            .O(N__54703),
            .I(N__54700));
    Span4Mux_v I__12900 (
            .O(N__54700),
            .I(N__54697));
    Odrv4 I__12899 (
            .O(N__54697),
            .I(comm_buf_4_1));
    CEMux I__12898 (
            .O(N__54694),
            .I(N__54691));
    LocalMux I__12897 (
            .O(N__54691),
            .I(n12892));
    SRMux I__12896 (
            .O(N__54688),
            .I(N__54685));
    LocalMux I__12895 (
            .O(N__54685),
            .I(N__54682));
    Span4Mux_h I__12894 (
            .O(N__54682),
            .I(N__54679));
    Odrv4 I__12893 (
            .O(N__54679),
            .I(n15510));
    InMux I__12892 (
            .O(N__54676),
            .I(N__54673));
    LocalMux I__12891 (
            .O(N__54673),
            .I(N__54669));
    InMux I__12890 (
            .O(N__54672),
            .I(N__54666));
    Span4Mux_h I__12889 (
            .O(N__54669),
            .I(N__54663));
    LocalMux I__12888 (
            .O(N__54666),
            .I(data_idxvec_7));
    Odrv4 I__12887 (
            .O(N__54663),
            .I(data_idxvec_7));
    InMux I__12886 (
            .O(N__54658),
            .I(N__54654));
    InMux I__12885 (
            .O(N__54657),
            .I(N__54651));
    LocalMux I__12884 (
            .O(N__54654),
            .I(N__54647));
    LocalMux I__12883 (
            .O(N__54651),
            .I(N__54644));
    InMux I__12882 (
            .O(N__54650),
            .I(N__54641));
    Span4Mux_h I__12881 (
            .O(N__54647),
            .I(N__54638));
    Span4Mux_h I__12880 (
            .O(N__54644),
            .I(N__54635));
    LocalMux I__12879 (
            .O(N__54641),
            .I(data_cntvec_7));
    Odrv4 I__12878 (
            .O(N__54638),
            .I(data_cntvec_7));
    Odrv4 I__12877 (
            .O(N__54635),
            .I(data_cntvec_7));
    InMux I__12876 (
            .O(N__54628),
            .I(N__54625));
    LocalMux I__12875 (
            .O(N__54625),
            .I(N__54622));
    Odrv12 I__12874 (
            .O(N__54622),
            .I(buf_data_iac_15));
    CascadeMux I__12873 (
            .O(N__54619),
            .I(n26_adj_1716_cascade_));
    CascadeMux I__12872 (
            .O(N__54616),
            .I(n22263_cascade_));
    InMux I__12871 (
            .O(N__54613),
            .I(N__54603));
    InMux I__12870 (
            .O(N__54612),
            .I(N__54603));
    InMux I__12869 (
            .O(N__54611),
            .I(N__54596));
    InMux I__12868 (
            .O(N__54610),
            .I(N__54593));
    InMux I__12867 (
            .O(N__54609),
            .I(N__54590));
    InMux I__12866 (
            .O(N__54608),
            .I(N__54581));
    LocalMux I__12865 (
            .O(N__54603),
            .I(N__54578));
    InMux I__12864 (
            .O(N__54602),
            .I(N__54573));
    InMux I__12863 (
            .O(N__54601),
            .I(N__54573));
    InMux I__12862 (
            .O(N__54600),
            .I(N__54567));
    InMux I__12861 (
            .O(N__54599),
            .I(N__54567));
    LocalMux I__12860 (
            .O(N__54596),
            .I(N__54562));
    LocalMux I__12859 (
            .O(N__54593),
            .I(N__54562));
    LocalMux I__12858 (
            .O(N__54590),
            .I(N__54559));
    InMux I__12857 (
            .O(N__54589),
            .I(N__54550));
    InMux I__12856 (
            .O(N__54588),
            .I(N__54550));
    InMux I__12855 (
            .O(N__54587),
            .I(N__54550));
    InMux I__12854 (
            .O(N__54586),
            .I(N__54550));
    InMux I__12853 (
            .O(N__54585),
            .I(N__54547));
    InMux I__12852 (
            .O(N__54584),
            .I(N__54543));
    LocalMux I__12851 (
            .O(N__54581),
            .I(N__54534));
    Span4Mux_h I__12850 (
            .O(N__54578),
            .I(N__54529));
    LocalMux I__12849 (
            .O(N__54573),
            .I(N__54529));
    InMux I__12848 (
            .O(N__54572),
            .I(N__54522));
    LocalMux I__12847 (
            .O(N__54567),
            .I(N__54513));
    Span4Mux_v I__12846 (
            .O(N__54562),
            .I(N__54513));
    Span4Mux_v I__12845 (
            .O(N__54559),
            .I(N__54513));
    LocalMux I__12844 (
            .O(N__54550),
            .I(N__54513));
    LocalMux I__12843 (
            .O(N__54547),
            .I(N__54510));
    InMux I__12842 (
            .O(N__54546),
            .I(N__54507));
    LocalMux I__12841 (
            .O(N__54543),
            .I(N__54504));
    InMux I__12840 (
            .O(N__54542),
            .I(N__54495));
    InMux I__12839 (
            .O(N__54541),
            .I(N__54495));
    InMux I__12838 (
            .O(N__54540),
            .I(N__54495));
    InMux I__12837 (
            .O(N__54539),
            .I(N__54495));
    InMux I__12836 (
            .O(N__54538),
            .I(N__54490));
    InMux I__12835 (
            .O(N__54537),
            .I(N__54490));
    Span4Mux_h I__12834 (
            .O(N__54534),
            .I(N__54487));
    Span4Mux_h I__12833 (
            .O(N__54529),
            .I(N__54484));
    InMux I__12832 (
            .O(N__54528),
            .I(N__54475));
    InMux I__12831 (
            .O(N__54527),
            .I(N__54475));
    InMux I__12830 (
            .O(N__54526),
            .I(N__54475));
    InMux I__12829 (
            .O(N__54525),
            .I(N__54475));
    LocalMux I__12828 (
            .O(N__54522),
            .I(N__54468));
    Span4Mux_h I__12827 (
            .O(N__54513),
            .I(N__54468));
    Span4Mux_v I__12826 (
            .O(N__54510),
            .I(N__54468));
    LocalMux I__12825 (
            .O(N__54507),
            .I(N__54465));
    Span4Mux_h I__12824 (
            .O(N__54504),
            .I(N__54458));
    LocalMux I__12823 (
            .O(N__54495),
            .I(N__54458));
    LocalMux I__12822 (
            .O(N__54490),
            .I(N__54458));
    Odrv4 I__12821 (
            .O(N__54487),
            .I(comm_index_2));
    Odrv4 I__12820 (
            .O(N__54484),
            .I(comm_index_2));
    LocalMux I__12819 (
            .O(N__54475),
            .I(comm_index_2));
    Odrv4 I__12818 (
            .O(N__54468),
            .I(comm_index_2));
    Odrv4 I__12817 (
            .O(N__54465),
            .I(comm_index_2));
    Odrv4 I__12816 (
            .O(N__54458),
            .I(comm_index_2));
    CascadeMux I__12815 (
            .O(N__54445),
            .I(N__54441));
    InMux I__12814 (
            .O(N__54444),
            .I(N__54438));
    InMux I__12813 (
            .O(N__54441),
            .I(N__54435));
    LocalMux I__12812 (
            .O(N__54438),
            .I(n21956));
    LocalMux I__12811 (
            .O(N__54435),
            .I(n21956));
    InMux I__12810 (
            .O(N__54430),
            .I(N__54427));
    LocalMux I__12809 (
            .O(N__54427),
            .I(n21862));
    CascadeMux I__12808 (
            .O(N__54424),
            .I(N__54410));
    InMux I__12807 (
            .O(N__54423),
            .I(N__54402));
    InMux I__12806 (
            .O(N__54422),
            .I(N__54391));
    InMux I__12805 (
            .O(N__54421),
            .I(N__54391));
    InMux I__12804 (
            .O(N__54420),
            .I(N__54391));
    InMux I__12803 (
            .O(N__54419),
            .I(N__54388));
    CascadeMux I__12802 (
            .O(N__54418),
            .I(N__54385));
    CascadeMux I__12801 (
            .O(N__54417),
            .I(N__54382));
    InMux I__12800 (
            .O(N__54416),
            .I(N__54373));
    InMux I__12799 (
            .O(N__54415),
            .I(N__54373));
    InMux I__12798 (
            .O(N__54414),
            .I(N__54373));
    InMux I__12797 (
            .O(N__54413),
            .I(N__54373));
    InMux I__12796 (
            .O(N__54410),
            .I(N__54367));
    InMux I__12795 (
            .O(N__54409),
            .I(N__54364));
    InMux I__12794 (
            .O(N__54408),
            .I(N__54353));
    InMux I__12793 (
            .O(N__54407),
            .I(N__54353));
    InMux I__12792 (
            .O(N__54406),
            .I(N__54353));
    InMux I__12791 (
            .O(N__54405),
            .I(N__54353));
    LocalMux I__12790 (
            .O(N__54402),
            .I(N__54350));
    InMux I__12789 (
            .O(N__54401),
            .I(N__54341));
    InMux I__12788 (
            .O(N__54400),
            .I(N__54341));
    InMux I__12787 (
            .O(N__54399),
            .I(N__54341));
    InMux I__12786 (
            .O(N__54398),
            .I(N__54341));
    LocalMux I__12785 (
            .O(N__54391),
            .I(N__54338));
    LocalMux I__12784 (
            .O(N__54388),
            .I(N__54335));
    InMux I__12783 (
            .O(N__54385),
            .I(N__54332));
    InMux I__12782 (
            .O(N__54382),
            .I(N__54327));
    LocalMux I__12781 (
            .O(N__54373),
            .I(N__54323));
    InMux I__12780 (
            .O(N__54372),
            .I(N__54316));
    InMux I__12779 (
            .O(N__54371),
            .I(N__54316));
    InMux I__12778 (
            .O(N__54370),
            .I(N__54316));
    LocalMux I__12777 (
            .O(N__54367),
            .I(N__54313));
    LocalMux I__12776 (
            .O(N__54364),
            .I(N__54303));
    InMux I__12775 (
            .O(N__54363),
            .I(N__54298));
    InMux I__12774 (
            .O(N__54362),
            .I(N__54298));
    LocalMux I__12773 (
            .O(N__54353),
            .I(N__54293));
    Span4Mux_v I__12772 (
            .O(N__54350),
            .I(N__54293));
    LocalMux I__12771 (
            .O(N__54341),
            .I(N__54290));
    Span4Mux_v I__12770 (
            .O(N__54338),
            .I(N__54287));
    Span4Mux_h I__12769 (
            .O(N__54335),
            .I(N__54282));
    LocalMux I__12768 (
            .O(N__54332),
            .I(N__54282));
    InMux I__12767 (
            .O(N__54331),
            .I(N__54277));
    InMux I__12766 (
            .O(N__54330),
            .I(N__54277));
    LocalMux I__12765 (
            .O(N__54327),
            .I(N__54274));
    InMux I__12764 (
            .O(N__54326),
            .I(N__54271));
    Span4Mux_v I__12763 (
            .O(N__54323),
            .I(N__54264));
    LocalMux I__12762 (
            .O(N__54316),
            .I(N__54264));
    Span4Mux_h I__12761 (
            .O(N__54313),
            .I(N__54264));
    InMux I__12760 (
            .O(N__54312),
            .I(N__54259));
    InMux I__12759 (
            .O(N__54311),
            .I(N__54259));
    InMux I__12758 (
            .O(N__54310),
            .I(N__54254));
    InMux I__12757 (
            .O(N__54309),
            .I(N__54254));
    InMux I__12756 (
            .O(N__54308),
            .I(N__54251));
    InMux I__12755 (
            .O(N__54307),
            .I(N__54246));
    InMux I__12754 (
            .O(N__54306),
            .I(N__54246));
    Span4Mux_h I__12753 (
            .O(N__54303),
            .I(N__54243));
    LocalMux I__12752 (
            .O(N__54298),
            .I(N__54234));
    Span4Mux_h I__12751 (
            .O(N__54293),
            .I(N__54234));
    Span4Mux_v I__12750 (
            .O(N__54290),
            .I(N__54234));
    Span4Mux_h I__12749 (
            .O(N__54287),
            .I(N__54234));
    Span4Mux_h I__12748 (
            .O(N__54282),
            .I(N__54231));
    LocalMux I__12747 (
            .O(N__54277),
            .I(N__54220));
    Span4Mux_h I__12746 (
            .O(N__54274),
            .I(N__54220));
    LocalMux I__12745 (
            .O(N__54271),
            .I(N__54220));
    Span4Mux_h I__12744 (
            .O(N__54264),
            .I(N__54220));
    LocalMux I__12743 (
            .O(N__54259),
            .I(N__54220));
    LocalMux I__12742 (
            .O(N__54254),
            .I(comm_index_0));
    LocalMux I__12741 (
            .O(N__54251),
            .I(comm_index_0));
    LocalMux I__12740 (
            .O(N__54246),
            .I(comm_index_0));
    Odrv4 I__12739 (
            .O(N__54243),
            .I(comm_index_0));
    Odrv4 I__12738 (
            .O(N__54234),
            .I(comm_index_0));
    Odrv4 I__12737 (
            .O(N__54231),
            .I(comm_index_0));
    Odrv4 I__12736 (
            .O(N__54220),
            .I(comm_index_0));
    CascadeMux I__12735 (
            .O(N__54205),
            .I(n21862_cascade_));
    InMux I__12734 (
            .O(N__54202),
            .I(N__54199));
    LocalMux I__12733 (
            .O(N__54199),
            .I(N__54195));
    InMux I__12732 (
            .O(N__54198),
            .I(N__54192));
    Span4Mux_h I__12731 (
            .O(N__54195),
            .I(N__54189));
    LocalMux I__12730 (
            .O(N__54192),
            .I(n30_adj_1720));
    Odrv4 I__12729 (
            .O(N__54189),
            .I(n30_adj_1720));
    CascadeMux I__12728 (
            .O(N__54184),
            .I(N__54179));
    CascadeMux I__12727 (
            .O(N__54183),
            .I(N__54176));
    InMux I__12726 (
            .O(N__54182),
            .I(N__54172));
    InMux I__12725 (
            .O(N__54179),
            .I(N__54168));
    InMux I__12724 (
            .O(N__54176),
            .I(N__54165));
    InMux I__12723 (
            .O(N__54175),
            .I(N__54162));
    LocalMux I__12722 (
            .O(N__54172),
            .I(N__54156));
    InMux I__12721 (
            .O(N__54171),
            .I(N__54153));
    LocalMux I__12720 (
            .O(N__54168),
            .I(N__54150));
    LocalMux I__12719 (
            .O(N__54165),
            .I(N__54145));
    LocalMux I__12718 (
            .O(N__54162),
            .I(N__54145));
    CascadeMux I__12717 (
            .O(N__54161),
            .I(N__54142));
    InMux I__12716 (
            .O(N__54160),
            .I(N__54137));
    InMux I__12715 (
            .O(N__54159),
            .I(N__54137));
    Span4Mux_h I__12714 (
            .O(N__54156),
            .I(N__54131));
    LocalMux I__12713 (
            .O(N__54153),
            .I(N__54131));
    Span4Mux_v I__12712 (
            .O(N__54150),
            .I(N__54128));
    Span4Mux_h I__12711 (
            .O(N__54145),
            .I(N__54125));
    InMux I__12710 (
            .O(N__54142),
            .I(N__54122));
    LocalMux I__12709 (
            .O(N__54137),
            .I(N__54119));
    InMux I__12708 (
            .O(N__54136),
            .I(N__54116));
    Span4Mux_h I__12707 (
            .O(N__54131),
            .I(N__54113));
    Span4Mux_h I__12706 (
            .O(N__54128),
            .I(N__54110));
    Span4Mux_v I__12705 (
            .O(N__54125),
            .I(N__54101));
    LocalMux I__12704 (
            .O(N__54122),
            .I(N__54101));
    Span4Mux_h I__12703 (
            .O(N__54119),
            .I(N__54101));
    LocalMux I__12702 (
            .O(N__54116),
            .I(N__54101));
    Span4Mux_v I__12701 (
            .O(N__54113),
            .I(N__54098));
    Odrv4 I__12700 (
            .O(N__54110),
            .I(n21968));
    Odrv4 I__12699 (
            .O(N__54101),
            .I(n21968));
    Odrv4 I__12698 (
            .O(N__54098),
            .I(n21968));
    CascadeMux I__12697 (
            .O(N__54091),
            .I(n22_adj_1725_cascade_));
    CascadeMux I__12696 (
            .O(N__54088),
            .I(n12677_cascade_));
    InMux I__12695 (
            .O(N__54085),
            .I(N__54082));
    LocalMux I__12694 (
            .O(N__54082),
            .I(N__54078));
    InMux I__12693 (
            .O(N__54081),
            .I(N__54075));
    Span4Mux_h I__12692 (
            .O(N__54078),
            .I(N__54072));
    LocalMux I__12691 (
            .O(N__54075),
            .I(N__54069));
    Sp12to4 I__12690 (
            .O(N__54072),
            .I(N__54060));
    Sp12to4 I__12689 (
            .O(N__54069),
            .I(N__54060));
    InMux I__12688 (
            .O(N__54068),
            .I(N__54057));
    InMux I__12687 (
            .O(N__54067),
            .I(N__54052));
    InMux I__12686 (
            .O(N__54066),
            .I(N__54052));
    InMux I__12685 (
            .O(N__54065),
            .I(N__54049));
    Span12Mux_v I__12684 (
            .O(N__54060),
            .I(N__54044));
    LocalMux I__12683 (
            .O(N__54057),
            .I(N__54044));
    LocalMux I__12682 (
            .O(N__54052),
            .I(n21895));
    LocalMux I__12681 (
            .O(N__54049),
            .I(n21895));
    Odrv12 I__12680 (
            .O(N__54044),
            .I(n21895));
    InMux I__12679 (
            .O(N__54037),
            .I(N__54034));
    LocalMux I__12678 (
            .O(N__54034),
            .I(N__54031));
    Span12Mux_v I__12677 (
            .O(N__54031),
            .I(N__54028));
    Odrv12 I__12676 (
            .O(N__54028),
            .I(buf_data_vac_8));
    InMux I__12675 (
            .O(N__54025),
            .I(N__54017));
    InMux I__12674 (
            .O(N__54024),
            .I(N__54012));
    InMux I__12673 (
            .O(N__54023),
            .I(N__54009));
    InMux I__12672 (
            .O(N__54022),
            .I(N__54006));
    InMux I__12671 (
            .O(N__54021),
            .I(N__54003));
    InMux I__12670 (
            .O(N__54020),
            .I(N__54000));
    LocalMux I__12669 (
            .O(N__54017),
            .I(N__53997));
    InMux I__12668 (
            .O(N__54016),
            .I(N__53994));
    InMux I__12667 (
            .O(N__54015),
            .I(N__53991));
    LocalMux I__12666 (
            .O(N__54012),
            .I(N__53987));
    LocalMux I__12665 (
            .O(N__54009),
            .I(N__53984));
    LocalMux I__12664 (
            .O(N__54006),
            .I(N__53979));
    LocalMux I__12663 (
            .O(N__54003),
            .I(N__53979));
    LocalMux I__12662 (
            .O(N__54000),
            .I(N__53970));
    Span4Mux_h I__12661 (
            .O(N__53997),
            .I(N__53970));
    LocalMux I__12660 (
            .O(N__53994),
            .I(N__53970));
    LocalMux I__12659 (
            .O(N__53991),
            .I(N__53970));
    InMux I__12658 (
            .O(N__53990),
            .I(N__53967));
    Span4Mux_v I__12657 (
            .O(N__53987),
            .I(N__53964));
    Span4Mux_v I__12656 (
            .O(N__53984),
            .I(N__53961));
    Span4Mux_v I__12655 (
            .O(N__53979),
            .I(N__53958));
    Span4Mux_v I__12654 (
            .O(N__53970),
            .I(N__53953));
    LocalMux I__12653 (
            .O(N__53967),
            .I(N__53953));
    Span4Mux_h I__12652 (
            .O(N__53964),
            .I(N__53948));
    Span4Mux_v I__12651 (
            .O(N__53961),
            .I(N__53948));
    Span4Mux_v I__12650 (
            .O(N__53958),
            .I(N__53943));
    Span4Mux_v I__12649 (
            .O(N__53953),
            .I(N__53943));
    Odrv4 I__12648 (
            .O(N__53948),
            .I(comm_rx_buf_0));
    Odrv4 I__12647 (
            .O(N__53943),
            .I(comm_rx_buf_0));
    InMux I__12646 (
            .O(N__53938),
            .I(N__53935));
    LocalMux I__12645 (
            .O(N__53935),
            .I(N__53932));
    Span4Mux_v I__12644 (
            .O(N__53932),
            .I(N__53929));
    Span4Mux_h I__12643 (
            .O(N__53929),
            .I(N__53926));
    Span4Mux_v I__12642 (
            .O(N__53926),
            .I(N__53923));
    Odrv4 I__12641 (
            .O(N__53923),
            .I(comm_buf_4_0));
    InMux I__12640 (
            .O(N__53920),
            .I(N__53917));
    LocalMux I__12639 (
            .O(N__53917),
            .I(N__53914));
    Span4Mux_v I__12638 (
            .O(N__53914),
            .I(N__53911));
    Odrv4 I__12637 (
            .O(N__53911),
            .I(buf_data_vac_15));
    InMux I__12636 (
            .O(N__53908),
            .I(N__53905));
    LocalMux I__12635 (
            .O(N__53905),
            .I(N__53902));
    Span12Mux_v I__12634 (
            .O(N__53902),
            .I(N__53899));
    Odrv12 I__12633 (
            .O(N__53899),
            .I(comm_buf_4_7));
    InMux I__12632 (
            .O(N__53896),
            .I(N__53890));
    InMux I__12631 (
            .O(N__53895),
            .I(N__53887));
    CascadeMux I__12630 (
            .O(N__53894),
            .I(N__53884));
    CascadeMux I__12629 (
            .O(N__53893),
            .I(N__53880));
    LocalMux I__12628 (
            .O(N__53890),
            .I(N__53874));
    LocalMux I__12627 (
            .O(N__53887),
            .I(N__53874));
    InMux I__12626 (
            .O(N__53884),
            .I(N__53871));
    InMux I__12625 (
            .O(N__53883),
            .I(N__53868));
    InMux I__12624 (
            .O(N__53880),
            .I(N__53865));
    InMux I__12623 (
            .O(N__53879),
            .I(N__53862));
    Span4Mux_v I__12622 (
            .O(N__53874),
            .I(N__53857));
    LocalMux I__12621 (
            .O(N__53871),
            .I(N__53857));
    LocalMux I__12620 (
            .O(N__53868),
            .I(N__53852));
    LocalMux I__12619 (
            .O(N__53865),
            .I(N__53847));
    LocalMux I__12618 (
            .O(N__53862),
            .I(N__53847));
    Span4Mux_h I__12617 (
            .O(N__53857),
            .I(N__53844));
    InMux I__12616 (
            .O(N__53856),
            .I(N__53841));
    InMux I__12615 (
            .O(N__53855),
            .I(N__53838));
    Span4Mux_v I__12614 (
            .O(N__53852),
            .I(N__53834));
    Span12Mux_v I__12613 (
            .O(N__53847),
            .I(N__53827));
    Sp12to4 I__12612 (
            .O(N__53844),
            .I(N__53827));
    LocalMux I__12611 (
            .O(N__53841),
            .I(N__53827));
    LocalMux I__12610 (
            .O(N__53838),
            .I(N__53824));
    InMux I__12609 (
            .O(N__53837),
            .I(N__53821));
    Odrv4 I__12608 (
            .O(N__53834),
            .I(comm_rx_buf_6));
    Odrv12 I__12607 (
            .O(N__53827),
            .I(comm_rx_buf_6));
    Odrv12 I__12606 (
            .O(N__53824),
            .I(comm_rx_buf_6));
    LocalMux I__12605 (
            .O(N__53821),
            .I(comm_rx_buf_6));
    InMux I__12604 (
            .O(N__53812),
            .I(N__53809));
    LocalMux I__12603 (
            .O(N__53809),
            .I(N__53806));
    Span4Mux_h I__12602 (
            .O(N__53806),
            .I(N__53803));
    Odrv4 I__12601 (
            .O(N__53803),
            .I(buf_data_vac_14));
    InMux I__12600 (
            .O(N__53800),
            .I(N__53797));
    LocalMux I__12599 (
            .O(N__53797),
            .I(N__53794));
    Span4Mux_v I__12598 (
            .O(N__53794),
            .I(N__53791));
    Sp12to4 I__12597 (
            .O(N__53791),
            .I(N__53788));
    Odrv12 I__12596 (
            .O(N__53788),
            .I(comm_buf_4_6));
    InMux I__12595 (
            .O(N__53785),
            .I(N__53782));
    LocalMux I__12594 (
            .O(N__53782),
            .I(N__53772));
    InMux I__12593 (
            .O(N__53781),
            .I(N__53756));
    InMux I__12592 (
            .O(N__53780),
            .I(N__53756));
    InMux I__12591 (
            .O(N__53779),
            .I(N__53756));
    InMux I__12590 (
            .O(N__53778),
            .I(N__53756));
    InMux I__12589 (
            .O(N__53777),
            .I(N__53756));
    InMux I__12588 (
            .O(N__53776),
            .I(N__53756));
    InMux I__12587 (
            .O(N__53775),
            .I(N__53756));
    Span4Mux_v I__12586 (
            .O(N__53772),
            .I(N__53753));
    InMux I__12585 (
            .O(N__53771),
            .I(N__53750));
    LocalMux I__12584 (
            .O(N__53756),
            .I(N__53747));
    Odrv4 I__12583 (
            .O(N__53753),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__12582 (
            .O(N__53750),
            .I(\comm_spi.bit_cnt_3 ));
    Odrv12 I__12581 (
            .O(N__53747),
            .I(\comm_spi.bit_cnt_3 ));
    InMux I__12580 (
            .O(N__53740),
            .I(N__53730));
    InMux I__12579 (
            .O(N__53739),
            .I(N__53715));
    InMux I__12578 (
            .O(N__53738),
            .I(N__53715));
    InMux I__12577 (
            .O(N__53737),
            .I(N__53715));
    InMux I__12576 (
            .O(N__53736),
            .I(N__53715));
    InMux I__12575 (
            .O(N__53735),
            .I(N__53715));
    InMux I__12574 (
            .O(N__53734),
            .I(N__53715));
    InMux I__12573 (
            .O(N__53733),
            .I(N__53715));
    LocalMux I__12572 (
            .O(N__53730),
            .I(\comm_spi.n18536 ));
    LocalMux I__12571 (
            .O(N__53715),
            .I(\comm_spi.n18536 ));
    ClkMux I__12570 (
            .O(N__53710),
            .I(N__53707));
    LocalMux I__12569 (
            .O(N__53707),
            .I(N__53703));
    ClkMux I__12568 (
            .O(N__53706),
            .I(N__53700));
    Span4Mux_h I__12567 (
            .O(N__53703),
            .I(N__53692));
    LocalMux I__12566 (
            .O(N__53700),
            .I(N__53692));
    ClkMux I__12565 (
            .O(N__53699),
            .I(N__53685));
    ClkMux I__12564 (
            .O(N__53698),
            .I(N__53682));
    ClkMux I__12563 (
            .O(N__53697),
            .I(N__53679));
    Span4Mux_v I__12562 (
            .O(N__53692),
            .I(N__53674));
    ClkMux I__12561 (
            .O(N__53691),
            .I(N__53671));
    ClkMux I__12560 (
            .O(N__53690),
            .I(N__53667));
    ClkMux I__12559 (
            .O(N__53689),
            .I(N__53662));
    ClkMux I__12558 (
            .O(N__53688),
            .I(N__53659));
    LocalMux I__12557 (
            .O(N__53685),
            .I(N__53656));
    LocalMux I__12556 (
            .O(N__53682),
            .I(N__53653));
    LocalMux I__12555 (
            .O(N__53679),
            .I(N__53650));
    ClkMux I__12554 (
            .O(N__53678),
            .I(N__53647));
    ClkMux I__12553 (
            .O(N__53677),
            .I(N__53644));
    Span4Mux_h I__12552 (
            .O(N__53674),
            .I(N__53639));
    LocalMux I__12551 (
            .O(N__53671),
            .I(N__53639));
    ClkMux I__12550 (
            .O(N__53670),
            .I(N__53635));
    LocalMux I__12549 (
            .O(N__53667),
            .I(N__53631));
    ClkMux I__12548 (
            .O(N__53666),
            .I(N__53628));
    ClkMux I__12547 (
            .O(N__53665),
            .I(N__53624));
    LocalMux I__12546 (
            .O(N__53662),
            .I(N__53621));
    LocalMux I__12545 (
            .O(N__53659),
            .I(N__53618));
    Span4Mux_v I__12544 (
            .O(N__53656),
            .I(N__53614));
    Span4Mux_v I__12543 (
            .O(N__53653),
            .I(N__53609));
    Span4Mux_v I__12542 (
            .O(N__53650),
            .I(N__53609));
    LocalMux I__12541 (
            .O(N__53647),
            .I(N__53606));
    LocalMux I__12540 (
            .O(N__53644),
            .I(N__53603));
    Span4Mux_v I__12539 (
            .O(N__53639),
            .I(N__53598));
    ClkMux I__12538 (
            .O(N__53638),
            .I(N__53595));
    LocalMux I__12537 (
            .O(N__53635),
            .I(N__53592));
    ClkMux I__12536 (
            .O(N__53634),
            .I(N__53589));
    Span4Mux_h I__12535 (
            .O(N__53631),
            .I(N__53583));
    LocalMux I__12534 (
            .O(N__53628),
            .I(N__53583));
    ClkMux I__12533 (
            .O(N__53627),
            .I(N__53580));
    LocalMux I__12532 (
            .O(N__53624),
            .I(N__53577));
    Span4Mux_h I__12531 (
            .O(N__53621),
            .I(N__53572));
    Span4Mux_h I__12530 (
            .O(N__53618),
            .I(N__53572));
    ClkMux I__12529 (
            .O(N__53617),
            .I(N__53569));
    Span4Mux_h I__12528 (
            .O(N__53614),
            .I(N__53561));
    Span4Mux_v I__12527 (
            .O(N__53609),
            .I(N__53561));
    Span4Mux_v I__12526 (
            .O(N__53606),
            .I(N__53561));
    Span4Mux_v I__12525 (
            .O(N__53603),
            .I(N__53558));
    ClkMux I__12524 (
            .O(N__53602),
            .I(N__53555));
    ClkMux I__12523 (
            .O(N__53601),
            .I(N__53552));
    Span4Mux_v I__12522 (
            .O(N__53598),
            .I(N__53547));
    LocalMux I__12521 (
            .O(N__53595),
            .I(N__53547));
    Span4Mux_v I__12520 (
            .O(N__53592),
            .I(N__53542));
    LocalMux I__12519 (
            .O(N__53589),
            .I(N__53542));
    ClkMux I__12518 (
            .O(N__53588),
            .I(N__53539));
    Span4Mux_v I__12517 (
            .O(N__53583),
            .I(N__53534));
    LocalMux I__12516 (
            .O(N__53580),
            .I(N__53534));
    Span4Mux_h I__12515 (
            .O(N__53577),
            .I(N__53531));
    Span4Mux_h I__12514 (
            .O(N__53572),
            .I(N__53526));
    LocalMux I__12513 (
            .O(N__53569),
            .I(N__53526));
    ClkMux I__12512 (
            .O(N__53568),
            .I(N__53523));
    Span4Mux_h I__12511 (
            .O(N__53561),
            .I(N__53520));
    Span4Mux_v I__12510 (
            .O(N__53558),
            .I(N__53517));
    LocalMux I__12509 (
            .O(N__53555),
            .I(N__53514));
    LocalMux I__12508 (
            .O(N__53552),
            .I(N__53511));
    Span4Mux_v I__12507 (
            .O(N__53547),
            .I(N__53504));
    Span4Mux_h I__12506 (
            .O(N__53542),
            .I(N__53504));
    LocalMux I__12505 (
            .O(N__53539),
            .I(N__53504));
    Span4Mux_h I__12504 (
            .O(N__53534),
            .I(N__53501));
    Span4Mux_h I__12503 (
            .O(N__53531),
            .I(N__53496));
    Span4Mux_v I__12502 (
            .O(N__53526),
            .I(N__53496));
    LocalMux I__12501 (
            .O(N__53523),
            .I(N__53493));
    Span4Mux_v I__12500 (
            .O(N__53520),
            .I(N__53490));
    Span4Mux_h I__12499 (
            .O(N__53517),
            .I(N__53485));
    Span4Mux_v I__12498 (
            .O(N__53514),
            .I(N__53485));
    Span4Mux_v I__12497 (
            .O(N__53511),
            .I(N__53480));
    Span4Mux_h I__12496 (
            .O(N__53504),
            .I(N__53480));
    Sp12to4 I__12495 (
            .O(N__53501),
            .I(N__53473));
    Sp12to4 I__12494 (
            .O(N__53496),
            .I(N__53473));
    Sp12to4 I__12493 (
            .O(N__53493),
            .I(N__53473));
    Odrv4 I__12492 (
            .O(N__53490),
            .I(\comm_spi.iclk ));
    Odrv4 I__12491 (
            .O(N__53485),
            .I(\comm_spi.iclk ));
    Odrv4 I__12490 (
            .O(N__53480),
            .I(\comm_spi.iclk ));
    Odrv12 I__12489 (
            .O(N__53473),
            .I(\comm_spi.iclk ));
    InMux I__12488 (
            .O(N__53464),
            .I(N__53461));
    LocalMux I__12487 (
            .O(N__53461),
            .I(N__53458));
    Odrv4 I__12486 (
            .O(N__53458),
            .I(n22330));
    CascadeMux I__12485 (
            .O(N__53455),
            .I(N__53452));
    InMux I__12484 (
            .O(N__53452),
            .I(N__53449));
    LocalMux I__12483 (
            .O(N__53449),
            .I(n22329));
    InMux I__12482 (
            .O(N__53446),
            .I(N__53443));
    LocalMux I__12481 (
            .O(N__53443),
            .I(N__53440));
    Span4Mux_v I__12480 (
            .O(N__53440),
            .I(N__53435));
    InMux I__12479 (
            .O(N__53439),
            .I(N__53432));
    InMux I__12478 (
            .O(N__53438),
            .I(N__53429));
    Span4Mux_h I__12477 (
            .O(N__53435),
            .I(N__53426));
    LocalMux I__12476 (
            .O(N__53432),
            .I(n15261));
    LocalMux I__12475 (
            .O(N__53429),
            .I(n15261));
    Odrv4 I__12474 (
            .O(N__53426),
            .I(n15261));
    CascadeMux I__12473 (
            .O(N__53419),
            .I(n22321_cascade_));
    CascadeMux I__12472 (
            .O(N__53416),
            .I(N__53413));
    InMux I__12471 (
            .O(N__53413),
            .I(N__53410));
    LocalMux I__12470 (
            .O(N__53410),
            .I(N__53406));
    InMux I__12469 (
            .O(N__53409),
            .I(N__53403));
    Odrv4 I__12468 (
            .O(N__53406),
            .I(n14851));
    LocalMux I__12467 (
            .O(N__53403),
            .I(n14851));
    InMux I__12466 (
            .O(N__53398),
            .I(N__53395));
    LocalMux I__12465 (
            .O(N__53395),
            .I(n22352));
    InMux I__12464 (
            .O(N__53392),
            .I(N__53388));
    InMux I__12463 (
            .O(N__53391),
            .I(N__53385));
    LocalMux I__12462 (
            .O(N__53388),
            .I(dds0_mclkcnt_6));
    LocalMux I__12461 (
            .O(N__53385),
            .I(dds0_mclkcnt_6));
    IoInMux I__12460 (
            .O(N__53380),
            .I(N__53377));
    LocalMux I__12459 (
            .O(N__53377),
            .I(N__53374));
    Span4Mux_s3_v I__12458 (
            .O(N__53374),
            .I(N__53371));
    Span4Mux_v I__12457 (
            .O(N__53371),
            .I(N__53368));
    Sp12to4 I__12456 (
            .O(N__53368),
            .I(N__53365));
    Span12Mux_v I__12455 (
            .O(N__53365),
            .I(N__53361));
    InMux I__12454 (
            .O(N__53364),
            .I(N__53358));
    Odrv12 I__12453 (
            .O(N__53361),
            .I(DDS_MCLK));
    LocalMux I__12452 (
            .O(N__53358),
            .I(DDS_MCLK));
    CascadeMux I__12451 (
            .O(N__53353),
            .I(n6888_cascade_));
    InMux I__12450 (
            .O(N__53350),
            .I(N__53346));
    InMux I__12449 (
            .O(N__53349),
            .I(N__53343));
    LocalMux I__12448 (
            .O(N__53346),
            .I(n21865));
    LocalMux I__12447 (
            .O(N__53343),
            .I(n21865));
    CascadeMux I__12446 (
            .O(N__53338),
            .I(N__53335));
    InMux I__12445 (
            .O(N__53335),
            .I(N__53332));
    LocalMux I__12444 (
            .O(N__53332),
            .I(N__53329));
    Odrv4 I__12443 (
            .O(N__53329),
            .I(n21981));
    InMux I__12442 (
            .O(N__53326),
            .I(N__53323));
    LocalMux I__12441 (
            .O(N__53323),
            .I(n22027));
    InMux I__12440 (
            .O(N__53320),
            .I(N__53317));
    LocalMux I__12439 (
            .O(N__53317),
            .I(n22018));
    InMux I__12438 (
            .O(N__53314),
            .I(N__53310));
    InMux I__12437 (
            .O(N__53313),
            .I(N__53307));
    LocalMux I__12436 (
            .O(N__53310),
            .I(dds0_mclkcnt_3));
    LocalMux I__12435 (
            .O(N__53307),
            .I(dds0_mclkcnt_3));
    InMux I__12434 (
            .O(N__53302),
            .I(N__53298));
    InMux I__12433 (
            .O(N__53301),
            .I(N__53295));
    LocalMux I__12432 (
            .O(N__53298),
            .I(dds0_mclkcnt_5));
    LocalMux I__12431 (
            .O(N__53295),
            .I(dds0_mclkcnt_5));
    CascadeMux I__12430 (
            .O(N__53290),
            .I(N__53287));
    InMux I__12429 (
            .O(N__53287),
            .I(N__53283));
    InMux I__12428 (
            .O(N__53286),
            .I(N__53280));
    LocalMux I__12427 (
            .O(N__53283),
            .I(N__53277));
    LocalMux I__12426 (
            .O(N__53280),
            .I(dds0_mclkcnt_1));
    Odrv4 I__12425 (
            .O(N__53277),
            .I(dds0_mclkcnt_1));
    InMux I__12424 (
            .O(N__53272),
            .I(N__53268));
    InMux I__12423 (
            .O(N__53271),
            .I(N__53265));
    LocalMux I__12422 (
            .O(N__53268),
            .I(dds0_mclkcnt_4));
    LocalMux I__12421 (
            .O(N__53265),
            .I(dds0_mclkcnt_4));
    InMux I__12420 (
            .O(N__53260),
            .I(N__53256));
    InMux I__12419 (
            .O(N__53259),
            .I(N__53253));
    LocalMux I__12418 (
            .O(N__53256),
            .I(N__53250));
    LocalMux I__12417 (
            .O(N__53253),
            .I(dds0_mclkcnt_7));
    Odrv4 I__12416 (
            .O(N__53250),
            .I(dds0_mclkcnt_7));
    InMux I__12415 (
            .O(N__53245),
            .I(N__53241));
    InMux I__12414 (
            .O(N__53244),
            .I(N__53238));
    LocalMux I__12413 (
            .O(N__53241),
            .I(dds0_mclkcnt_0));
    LocalMux I__12412 (
            .O(N__53238),
            .I(dds0_mclkcnt_0));
    CascadeMux I__12411 (
            .O(N__53233),
            .I(n12_adj_1685_cascade_));
    InMux I__12410 (
            .O(N__53230),
            .I(N__53226));
    InMux I__12409 (
            .O(N__53229),
            .I(N__53223));
    LocalMux I__12408 (
            .O(N__53226),
            .I(dds0_mclkcnt_2));
    LocalMux I__12407 (
            .O(N__53223),
            .I(dds0_mclkcnt_2));
    InMux I__12406 (
            .O(N__53218),
            .I(N__53212));
    InMux I__12405 (
            .O(N__53217),
            .I(N__53212));
    LocalMux I__12404 (
            .O(N__53212),
            .I(n21857));
    InMux I__12403 (
            .O(N__53209),
            .I(bfn_19_7_0_));
    InMux I__12402 (
            .O(N__53206),
            .I(n20819));
    InMux I__12401 (
            .O(N__53203),
            .I(n20820));
    InMux I__12400 (
            .O(N__53200),
            .I(n20821));
    InMux I__12399 (
            .O(N__53197),
            .I(n20822));
    InMux I__12398 (
            .O(N__53194),
            .I(n20823));
    InMux I__12397 (
            .O(N__53191),
            .I(n20824));
    InMux I__12396 (
            .O(N__53188),
            .I(n20825));
    InMux I__12395 (
            .O(N__53185),
            .I(N__53182));
    LocalMux I__12394 (
            .O(N__53182),
            .I(n10));
    InMux I__12393 (
            .O(N__53179),
            .I(\ADC_VDC.genclk.n20757 ));
    InMux I__12392 (
            .O(N__53176),
            .I(bfn_19_6_0_));
    InMux I__12391 (
            .O(N__53173),
            .I(\ADC_VDC.genclk.n20759 ));
    InMux I__12390 (
            .O(N__53170),
            .I(\ADC_VDC.genclk.n20760 ));
    InMux I__12389 (
            .O(N__53167),
            .I(\ADC_VDC.genclk.n20761 ));
    InMux I__12388 (
            .O(N__53164),
            .I(\ADC_VDC.genclk.n20762 ));
    InMux I__12387 (
            .O(N__53161),
            .I(\ADC_VDC.genclk.n20763 ));
    InMux I__12386 (
            .O(N__53158),
            .I(\ADC_VDC.genclk.n20764 ));
    InMux I__12385 (
            .O(N__53155),
            .I(\ADC_VDC.genclk.n20765 ));
    InMux I__12384 (
            .O(N__53152),
            .I(N__53148));
    InMux I__12383 (
            .O(N__53151),
            .I(N__53145));
    LocalMux I__12382 (
            .O(N__53148),
            .I(N__53142));
    LocalMux I__12381 (
            .O(N__53145),
            .I(N__53139));
    Span4Mux_v I__12380 (
            .O(N__53142),
            .I(N__53136));
    Span4Mux_h I__12379 (
            .O(N__53139),
            .I(N__53133));
    Span4Mux_h I__12378 (
            .O(N__53136),
            .I(N__53130));
    Span4Mux_v I__12377 (
            .O(N__53133),
            .I(N__53127));
    Odrv4 I__12376 (
            .O(N__53130),
            .I(n7));
    Odrv4 I__12375 (
            .O(N__53127),
            .I(n7));
    CascadeMux I__12374 (
            .O(N__53122),
            .I(N__53119));
    CascadeBuf I__12373 (
            .O(N__53119),
            .I(N__53116));
    CascadeMux I__12372 (
            .O(N__53116),
            .I(N__53113));
    CascadeBuf I__12371 (
            .O(N__53113),
            .I(N__53110));
    CascadeMux I__12370 (
            .O(N__53110),
            .I(N__53107));
    CascadeBuf I__12369 (
            .O(N__53107),
            .I(N__53104));
    CascadeMux I__12368 (
            .O(N__53104),
            .I(N__53101));
    CascadeBuf I__12367 (
            .O(N__53101),
            .I(N__53098));
    CascadeMux I__12366 (
            .O(N__53098),
            .I(N__53095));
    CascadeBuf I__12365 (
            .O(N__53095),
            .I(N__53092));
    CascadeMux I__12364 (
            .O(N__53092),
            .I(N__53089));
    CascadeBuf I__12363 (
            .O(N__53089),
            .I(N__53086));
    CascadeMux I__12362 (
            .O(N__53086),
            .I(N__53083));
    CascadeBuf I__12361 (
            .O(N__53083),
            .I(N__53079));
    CascadeMux I__12360 (
            .O(N__53082),
            .I(N__53076));
    CascadeMux I__12359 (
            .O(N__53079),
            .I(N__53073));
    CascadeBuf I__12358 (
            .O(N__53076),
            .I(N__53070));
    CascadeBuf I__12357 (
            .O(N__53073),
            .I(N__53067));
    CascadeMux I__12356 (
            .O(N__53070),
            .I(N__53064));
    CascadeMux I__12355 (
            .O(N__53067),
            .I(N__53061));
    InMux I__12354 (
            .O(N__53064),
            .I(N__53058));
    CascadeBuf I__12353 (
            .O(N__53061),
            .I(N__53055));
    LocalMux I__12352 (
            .O(N__53058),
            .I(N__53052));
    CascadeMux I__12351 (
            .O(N__53055),
            .I(N__53049));
    Span12Mux_h I__12350 (
            .O(N__53052),
            .I(N__53046));
    InMux I__12349 (
            .O(N__53049),
            .I(N__53043));
    Span12Mux_v I__12348 (
            .O(N__53046),
            .I(N__53038));
    LocalMux I__12347 (
            .O(N__53043),
            .I(N__53038));
    Odrv12 I__12346 (
            .O(N__53038),
            .I(data_index_9_N_236_0));
    InMux I__12345 (
            .O(N__53035),
            .I(N__53032));
    LocalMux I__12344 (
            .O(N__53032),
            .I(N__53029));
    Odrv4 I__12343 (
            .O(N__53029),
            .I(buf_data_iac_20));
    InMux I__12342 (
            .O(N__53026),
            .I(N__53023));
    LocalMux I__12341 (
            .O(N__53023),
            .I(N__53020));
    Span12Mux_v I__12340 (
            .O(N__53020),
            .I(N__53017));
    Odrv12 I__12339 (
            .O(N__53017),
            .I(n22500));
    InMux I__12338 (
            .O(N__53014),
            .I(bfn_19_5_0_));
    InMux I__12337 (
            .O(N__53011),
            .I(\ADC_VDC.genclk.n20751 ));
    InMux I__12336 (
            .O(N__53008),
            .I(\ADC_VDC.genclk.n20752 ));
    InMux I__12335 (
            .O(N__53005),
            .I(\ADC_VDC.genclk.n20753 ));
    InMux I__12334 (
            .O(N__53002),
            .I(\ADC_VDC.genclk.n20754 ));
    InMux I__12333 (
            .O(N__52999),
            .I(\ADC_VDC.genclk.n20755 ));
    InMux I__12332 (
            .O(N__52996),
            .I(\ADC_VDC.genclk.n20756 ));
    CascadeMux I__12331 (
            .O(N__52993),
            .I(n22152_cascade_));
    InMux I__12330 (
            .O(N__52990),
            .I(N__52987));
    LocalMux I__12329 (
            .O(N__52987),
            .I(N__52984));
    Sp12to4 I__12328 (
            .O(N__52984),
            .I(N__52981));
    Span12Mux_v I__12327 (
            .O(N__52981),
            .I(N__52978));
    Span12Mux_h I__12326 (
            .O(N__52978),
            .I(N__52975));
    Odrv12 I__12325 (
            .O(N__52975),
            .I(n22149));
    CascadeMux I__12324 (
            .O(N__52972),
            .I(n23444_cascade_));
    InMux I__12323 (
            .O(N__52969),
            .I(N__52966));
    LocalMux I__12322 (
            .O(N__52966),
            .I(N__52963));
    Span4Mux_h I__12321 (
            .O(N__52963),
            .I(N__52960));
    Odrv4 I__12320 (
            .O(N__52960),
            .I(n22148));
    InMux I__12319 (
            .O(N__52957),
            .I(N__52954));
    LocalMux I__12318 (
            .O(N__52954),
            .I(N__52951));
    Span4Mux_h I__12317 (
            .O(N__52951),
            .I(N__52948));
    Span4Mux_h I__12316 (
            .O(N__52948),
            .I(N__52945));
    Odrv4 I__12315 (
            .O(N__52945),
            .I(n111_adj_1750));
    CascadeMux I__12314 (
            .O(N__52942),
            .I(n23447_cascade_));
    CascadeMux I__12313 (
            .O(N__52939),
            .I(comm_buf_1_7_N_559_2_cascade_));
    InMux I__12312 (
            .O(N__52936),
            .I(N__52931));
    CascadeMux I__12311 (
            .O(N__52935),
            .I(N__52928));
    InMux I__12310 (
            .O(N__52934),
            .I(N__52922));
    LocalMux I__12309 (
            .O(N__52931),
            .I(N__52919));
    InMux I__12308 (
            .O(N__52928),
            .I(N__52916));
    InMux I__12307 (
            .O(N__52927),
            .I(N__52913));
    InMux I__12306 (
            .O(N__52926),
            .I(N__52910));
    CascadeMux I__12305 (
            .O(N__52925),
            .I(N__52906));
    LocalMux I__12304 (
            .O(N__52922),
            .I(N__52901));
    Span4Mux_v I__12303 (
            .O(N__52919),
            .I(N__52901));
    LocalMux I__12302 (
            .O(N__52916),
            .I(N__52896));
    LocalMux I__12301 (
            .O(N__52913),
            .I(N__52896));
    LocalMux I__12300 (
            .O(N__52910),
            .I(N__52893));
    InMux I__12299 (
            .O(N__52909),
            .I(N__52890));
    InMux I__12298 (
            .O(N__52906),
            .I(N__52885));
    Span4Mux_v I__12297 (
            .O(N__52901),
            .I(N__52880));
    Span4Mux_v I__12296 (
            .O(N__52896),
            .I(N__52880));
    Span4Mux_v I__12295 (
            .O(N__52893),
            .I(N__52875));
    LocalMux I__12294 (
            .O(N__52890),
            .I(N__52875));
    InMux I__12293 (
            .O(N__52889),
            .I(N__52870));
    InMux I__12292 (
            .O(N__52888),
            .I(N__52870));
    LocalMux I__12291 (
            .O(N__52885),
            .I(N__52867));
    Span4Mux_h I__12290 (
            .O(N__52880),
            .I(N__52864));
    Span4Mux_v I__12289 (
            .O(N__52875),
            .I(N__52859));
    LocalMux I__12288 (
            .O(N__52870),
            .I(N__52859));
    Span4Mux_h I__12287 (
            .O(N__52867),
            .I(N__52856));
    Span4Mux_h I__12286 (
            .O(N__52864),
            .I(N__52853));
    Span4Mux_h I__12285 (
            .O(N__52859),
            .I(N__52850));
    Odrv4 I__12284 (
            .O(N__52856),
            .I(comm_buf_1_2));
    Odrv4 I__12283 (
            .O(N__52853),
            .I(comm_buf_1_2));
    Odrv4 I__12282 (
            .O(N__52850),
            .I(comm_buf_1_2));
    InMux I__12281 (
            .O(N__52843),
            .I(N__52839));
    CascadeMux I__12280 (
            .O(N__52842),
            .I(N__52836));
    LocalMux I__12279 (
            .O(N__52839),
            .I(N__52833));
    InMux I__12278 (
            .O(N__52836),
            .I(N__52829));
    Span4Mux_h I__12277 (
            .O(N__52833),
            .I(N__52826));
    InMux I__12276 (
            .O(N__52832),
            .I(N__52823));
    LocalMux I__12275 (
            .O(N__52829),
            .I(req_data_cnt_2));
    Odrv4 I__12274 (
            .O(N__52826),
            .I(req_data_cnt_2));
    LocalMux I__12273 (
            .O(N__52823),
            .I(req_data_cnt_2));
    CascadeMux I__12272 (
            .O(N__52816),
            .I(N__52813));
    InMux I__12271 (
            .O(N__52813),
            .I(N__52808));
    InMux I__12270 (
            .O(N__52812),
            .I(N__52805));
    CascadeMux I__12269 (
            .O(N__52811),
            .I(N__52802));
    LocalMux I__12268 (
            .O(N__52808),
            .I(N__52799));
    LocalMux I__12267 (
            .O(N__52805),
            .I(N__52796));
    InMux I__12266 (
            .O(N__52802),
            .I(N__52793));
    Odrv4 I__12265 (
            .O(N__52799),
            .I(acadc_skipCount_2));
    Odrv12 I__12264 (
            .O(N__52796),
            .I(acadc_skipCount_2));
    LocalMux I__12263 (
            .O(N__52793),
            .I(acadc_skipCount_2));
    InMux I__12262 (
            .O(N__52786),
            .I(N__52783));
    LocalMux I__12261 (
            .O(N__52783),
            .I(n22151));
    IoInMux I__12260 (
            .O(N__52780),
            .I(N__52776));
    InMux I__12259 (
            .O(N__52779),
            .I(N__52773));
    LocalMux I__12258 (
            .O(N__52776),
            .I(N__52770));
    LocalMux I__12257 (
            .O(N__52773),
            .I(N__52767));
    Span4Mux_s3_v I__12256 (
            .O(N__52770),
            .I(N__52764));
    Span4Mux_h I__12255 (
            .O(N__52767),
            .I(N__52760));
    Span4Mux_v I__12254 (
            .O(N__52764),
            .I(N__52757));
    InMux I__12253 (
            .O(N__52763),
            .I(N__52754));
    Span4Mux_h I__12252 (
            .O(N__52760),
            .I(N__52751));
    Odrv4 I__12251 (
            .O(N__52757),
            .I(SELIRNG1));
    LocalMux I__12250 (
            .O(N__52754),
            .I(SELIRNG1));
    Odrv4 I__12249 (
            .O(N__52751),
            .I(SELIRNG1));
    InMux I__12248 (
            .O(N__52744),
            .I(N__52739));
    CascadeMux I__12247 (
            .O(N__52743),
            .I(N__52736));
    InMux I__12246 (
            .O(N__52742),
            .I(N__52733));
    LocalMux I__12245 (
            .O(N__52739),
            .I(N__52730));
    InMux I__12244 (
            .O(N__52736),
            .I(N__52727));
    LocalMux I__12243 (
            .O(N__52733),
            .I(acadc_skipCount_11));
    Odrv12 I__12242 (
            .O(N__52730),
            .I(acadc_skipCount_11));
    LocalMux I__12241 (
            .O(N__52727),
            .I(acadc_skipCount_11));
    InMux I__12240 (
            .O(N__52720),
            .I(N__52717));
    LocalMux I__12239 (
            .O(N__52717),
            .I(N__52713));
    InMux I__12238 (
            .O(N__52716),
            .I(N__52710));
    Span4Mux_v I__12237 (
            .O(N__52713),
            .I(N__52705));
    LocalMux I__12236 (
            .O(N__52710),
            .I(N__52705));
    Span4Mux_h I__12235 (
            .O(N__52705),
            .I(N__52701));
    InMux I__12234 (
            .O(N__52704),
            .I(N__52698));
    Span4Mux_h I__12233 (
            .O(N__52701),
            .I(N__52695));
    LocalMux I__12232 (
            .O(N__52698),
            .I(buf_adcdata_iac_9));
    Odrv4 I__12231 (
            .O(N__52695),
            .I(buf_adcdata_iac_9));
    InMux I__12230 (
            .O(N__52690),
            .I(N__52687));
    LocalMux I__12229 (
            .O(N__52687),
            .I(N__52684));
    Odrv12 I__12228 (
            .O(N__52684),
            .I(n16_adj_1751));
    InMux I__12227 (
            .O(N__52681),
            .I(N__52678));
    LocalMux I__12226 (
            .O(N__52678),
            .I(N__52675));
    Span4Mux_v I__12225 (
            .O(N__52675),
            .I(N__52672));
    Odrv4 I__12224 (
            .O(N__52672),
            .I(n22136));
    InMux I__12223 (
            .O(N__52669),
            .I(N__52666));
    LocalMux I__12222 (
            .O(N__52666),
            .I(N__52663));
    Span12Mux_h I__12221 (
            .O(N__52663),
            .I(N__52660));
    Span12Mux_v I__12220 (
            .O(N__52660),
            .I(N__52655));
    InMux I__12219 (
            .O(N__52659),
            .I(N__52652));
    InMux I__12218 (
            .O(N__52658),
            .I(N__52649));
    Odrv12 I__12217 (
            .O(N__52655),
            .I(wdtick_flag));
    LocalMux I__12216 (
            .O(N__52652),
            .I(wdtick_flag));
    LocalMux I__12215 (
            .O(N__52649),
            .I(wdtick_flag));
    CascadeMux I__12214 (
            .O(N__52642),
            .I(N__52639));
    InMux I__12213 (
            .O(N__52639),
            .I(N__52635));
    InMux I__12212 (
            .O(N__52638),
            .I(N__52632));
    LocalMux I__12211 (
            .O(N__52635),
            .I(N__52629));
    LocalMux I__12210 (
            .O(N__52632),
            .I(N__52626));
    Span4Mux_h I__12209 (
            .O(N__52629),
            .I(N__52622));
    Span4Mux_v I__12208 (
            .O(N__52626),
            .I(N__52619));
    InMux I__12207 (
            .O(N__52625),
            .I(N__52616));
    Span4Mux_h I__12206 (
            .O(N__52622),
            .I(N__52613));
    Odrv4 I__12205 (
            .O(N__52619),
            .I(buf_control_0));
    LocalMux I__12204 (
            .O(N__52616),
            .I(buf_control_0));
    Odrv4 I__12203 (
            .O(N__52613),
            .I(buf_control_0));
    IoInMux I__12202 (
            .O(N__52606),
            .I(N__52603));
    LocalMux I__12201 (
            .O(N__52603),
            .I(N__52600));
    Span4Mux_s1_v I__12200 (
            .O(N__52600),
            .I(N__52597));
    Span4Mux_h I__12199 (
            .O(N__52597),
            .I(N__52594));
    Span4Mux_v I__12198 (
            .O(N__52594),
            .I(N__52591));
    Odrv4 I__12197 (
            .O(N__52591),
            .I(CONT_SD));
    InMux I__12196 (
            .O(N__52588),
            .I(N__52584));
    InMux I__12195 (
            .O(N__52587),
            .I(N__52581));
    LocalMux I__12194 (
            .O(N__52584),
            .I(N__52578));
    LocalMux I__12193 (
            .O(N__52581),
            .I(N__52575));
    Span4Mux_h I__12192 (
            .O(N__52578),
            .I(N__52572));
    Odrv4 I__12191 (
            .O(N__52575),
            .I(n8_adj_1605));
    Odrv4 I__12190 (
            .O(N__52572),
            .I(n8_adj_1605));
    InMux I__12189 (
            .O(N__52567),
            .I(N__52564));
    LocalMux I__12188 (
            .O(N__52564),
            .I(N__52560));
    InMux I__12187 (
            .O(N__52563),
            .I(N__52557));
    Span4Mux_h I__12186 (
            .O(N__52560),
            .I(N__52554));
    LocalMux I__12185 (
            .O(N__52557),
            .I(data_idxvec_4));
    Odrv4 I__12184 (
            .O(N__52554),
            .I(data_idxvec_4));
    InMux I__12183 (
            .O(N__52549),
            .I(N__52546));
    LocalMux I__12182 (
            .O(N__52546),
            .I(N__52542));
    InMux I__12181 (
            .O(N__52545),
            .I(N__52538));
    Span4Mux_h I__12180 (
            .O(N__52542),
            .I(N__52535));
    InMux I__12179 (
            .O(N__52541),
            .I(N__52532));
    LocalMux I__12178 (
            .O(N__52538),
            .I(data_cntvec_4));
    Odrv4 I__12177 (
            .O(N__52535),
            .I(data_cntvec_4));
    LocalMux I__12176 (
            .O(N__52532),
            .I(data_cntvec_4));
    InMux I__12175 (
            .O(N__52525),
            .I(N__52522));
    LocalMux I__12174 (
            .O(N__52522),
            .I(N__52519));
    Odrv12 I__12173 (
            .O(N__52519),
            .I(n22301));
    CascadeMux I__12172 (
            .O(N__52516),
            .I(n26_adj_1735_cascade_));
    CascadeMux I__12171 (
            .O(N__52513),
            .I(N__52509));
    InMux I__12170 (
            .O(N__52512),
            .I(N__52506));
    InMux I__12169 (
            .O(N__52509),
            .I(N__52502));
    LocalMux I__12168 (
            .O(N__52506),
            .I(N__52499));
    InMux I__12167 (
            .O(N__52505),
            .I(N__52496));
    LocalMux I__12166 (
            .O(N__52502),
            .I(acadc_skipCount_4));
    Odrv4 I__12165 (
            .O(N__52499),
            .I(acadc_skipCount_4));
    LocalMux I__12164 (
            .O(N__52496),
            .I(acadc_skipCount_4));
    CascadeMux I__12163 (
            .O(N__52489),
            .I(n23318_cascade_));
    InMux I__12162 (
            .O(N__52486),
            .I(N__52483));
    LocalMux I__12161 (
            .O(N__52483),
            .I(N__52478));
    InMux I__12160 (
            .O(N__52482),
            .I(N__52475));
    InMux I__12159 (
            .O(N__52481),
            .I(N__52472));
    Span4Mux_v I__12158 (
            .O(N__52478),
            .I(N__52467));
    LocalMux I__12157 (
            .O(N__52475),
            .I(N__52467));
    LocalMux I__12156 (
            .O(N__52472),
            .I(req_data_cnt_4));
    Odrv4 I__12155 (
            .O(N__52467),
            .I(req_data_cnt_4));
    InMux I__12154 (
            .O(N__52462),
            .I(N__52459));
    LocalMux I__12153 (
            .O(N__52459),
            .I(N__52456));
    Span4Mux_h I__12152 (
            .O(N__52456),
            .I(N__52453));
    Span4Mux_h I__12151 (
            .O(N__52453),
            .I(N__52450));
    Odrv4 I__12150 (
            .O(N__52450),
            .I(n23441));
    CascadeMux I__12149 (
            .O(N__52447),
            .I(n23321_cascade_));
    InMux I__12148 (
            .O(N__52444),
            .I(N__52441));
    LocalMux I__12147 (
            .O(N__52441),
            .I(N__52438));
    Span4Mux_v I__12146 (
            .O(N__52438),
            .I(N__52435));
    Span4Mux_h I__12145 (
            .O(N__52435),
            .I(N__52432));
    Span4Mux_h I__12144 (
            .O(N__52432),
            .I(N__52429));
    Odrv4 I__12143 (
            .O(N__52429),
            .I(n111_adj_1737));
    CascadeMux I__12142 (
            .O(N__52426),
            .I(n30_adj_1736_cascade_));
    CascadeMux I__12141 (
            .O(N__52423),
            .I(comm_buf_1_7_N_559_4_cascade_));
    InMux I__12140 (
            .O(N__52420),
            .I(N__52416));
    InMux I__12139 (
            .O(N__52419),
            .I(N__52413));
    LocalMux I__12138 (
            .O(N__52416),
            .I(N__52408));
    LocalMux I__12137 (
            .O(N__52413),
            .I(N__52408));
    Odrv4 I__12136 (
            .O(N__52408),
            .I(data_idxvec_2));
    CascadeMux I__12135 (
            .O(N__52405),
            .I(N__52402));
    InMux I__12134 (
            .O(N__52402),
            .I(N__52399));
    LocalMux I__12133 (
            .O(N__52399),
            .I(N__52394));
    InMux I__12132 (
            .O(N__52398),
            .I(N__52391));
    InMux I__12131 (
            .O(N__52397),
            .I(N__52388));
    Span4Mux_h I__12130 (
            .O(N__52394),
            .I(N__52385));
    LocalMux I__12129 (
            .O(N__52391),
            .I(data_cntvec_2));
    LocalMux I__12128 (
            .O(N__52388),
            .I(data_cntvec_2));
    Odrv4 I__12127 (
            .O(N__52385),
            .I(data_cntvec_2));
    InMux I__12126 (
            .O(N__52378),
            .I(N__52375));
    LocalMux I__12125 (
            .O(N__52375),
            .I(N__52372));
    Span4Mux_v I__12124 (
            .O(N__52372),
            .I(N__52369));
    Odrv4 I__12123 (
            .O(N__52369),
            .I(buf_data_iac_10));
    CascadeMux I__12122 (
            .O(N__52366),
            .I(n26_adj_1748_cascade_));
    CascadeMux I__12121 (
            .O(N__52363),
            .I(comm_buf_1_7_N_559_5_cascade_));
    InMux I__12120 (
            .O(N__52360),
            .I(N__52357));
    LocalMux I__12119 (
            .O(N__52357),
            .I(N__52354));
    Span4Mux_v I__12118 (
            .O(N__52354),
            .I(N__52351));
    Span4Mux_h I__12117 (
            .O(N__52351),
            .I(N__52348));
    Span4Mux_h I__12116 (
            .O(N__52348),
            .I(N__52345));
    Odrv4 I__12115 (
            .O(N__52345),
            .I(n16_adj_1728));
    CascadeMux I__12114 (
            .O(N__52342),
            .I(N__52338));
    InMux I__12113 (
            .O(N__52341),
            .I(N__52335));
    InMux I__12112 (
            .O(N__52338),
            .I(N__52332));
    LocalMux I__12111 (
            .O(N__52335),
            .I(N__52329));
    LocalMux I__12110 (
            .O(N__52332),
            .I(N__52326));
    Span4Mux_v I__12109 (
            .O(N__52329),
            .I(N__52323));
    Span4Mux_v I__12108 (
            .O(N__52326),
            .I(N__52320));
    Sp12to4 I__12107 (
            .O(N__52323),
            .I(N__52316));
    Span4Mux_h I__12106 (
            .O(N__52320),
            .I(N__52313));
    InMux I__12105 (
            .O(N__52319),
            .I(N__52310));
    Span12Mux_h I__12104 (
            .O(N__52316),
            .I(N__52307));
    Span4Mux_h I__12103 (
            .O(N__52313),
            .I(N__52304));
    LocalMux I__12102 (
            .O(N__52310),
            .I(buf_adcdata_iac_13));
    Odrv12 I__12101 (
            .O(N__52307),
            .I(buf_adcdata_iac_13));
    Odrv4 I__12100 (
            .O(N__52304),
            .I(buf_adcdata_iac_13));
    InMux I__12099 (
            .O(N__52297),
            .I(N__52294));
    LocalMux I__12098 (
            .O(N__52294),
            .I(N__52291));
    Span4Mux_h I__12097 (
            .O(N__52291),
            .I(N__52288));
    Span4Mux_h I__12096 (
            .O(N__52288),
            .I(N__52285));
    Odrv4 I__12095 (
            .O(N__52285),
            .I(n23354));
    InMux I__12094 (
            .O(N__52282),
            .I(N__52279));
    LocalMux I__12093 (
            .O(N__52279),
            .I(n23357));
    InMux I__12092 (
            .O(N__52276),
            .I(N__52273));
    LocalMux I__12091 (
            .O(N__52273),
            .I(N__52269));
    InMux I__12090 (
            .O(N__52272),
            .I(N__52266));
    Span4Mux_h I__12089 (
            .O(N__52269),
            .I(N__52263));
    LocalMux I__12088 (
            .O(N__52266),
            .I(data_idxvec_1));
    Odrv4 I__12087 (
            .O(N__52263),
            .I(data_idxvec_1));
    InMux I__12086 (
            .O(N__52258),
            .I(N__52254));
    InMux I__12085 (
            .O(N__52257),
            .I(N__52251));
    LocalMux I__12084 (
            .O(N__52254),
            .I(N__52248));
    LocalMux I__12083 (
            .O(N__52251),
            .I(N__52242));
    Span4Mux_v I__12082 (
            .O(N__52248),
            .I(N__52242));
    InMux I__12081 (
            .O(N__52247),
            .I(N__52239));
    Odrv4 I__12080 (
            .O(N__52242),
            .I(data_cntvec_1));
    LocalMux I__12079 (
            .O(N__52239),
            .I(data_cntvec_1));
    InMux I__12078 (
            .O(N__52234),
            .I(N__52230));
    InMux I__12077 (
            .O(N__52233),
            .I(N__52226));
    LocalMux I__12076 (
            .O(N__52230),
            .I(N__52223));
    InMux I__12075 (
            .O(N__52229),
            .I(N__52220));
    LocalMux I__12074 (
            .O(N__52226),
            .I(N__52215));
    Span4Mux_h I__12073 (
            .O(N__52223),
            .I(N__52215));
    LocalMux I__12072 (
            .O(N__52220),
            .I(N__52212));
    Odrv4 I__12071 (
            .O(N__52215),
            .I(acadc_skipCount_1));
    Odrv4 I__12070 (
            .O(N__52212),
            .I(acadc_skipCount_1));
    InMux I__12069 (
            .O(N__52207),
            .I(N__52202));
    CascadeMux I__12068 (
            .O(N__52206),
            .I(N__52199));
    InMux I__12067 (
            .O(N__52205),
            .I(N__52196));
    LocalMux I__12066 (
            .O(N__52202),
            .I(N__52193));
    InMux I__12065 (
            .O(N__52199),
            .I(N__52190));
    LocalMux I__12064 (
            .O(N__52196),
            .I(req_data_cnt_1));
    Odrv4 I__12063 (
            .O(N__52193),
            .I(req_data_cnt_1));
    LocalMux I__12062 (
            .O(N__52190),
            .I(req_data_cnt_1));
    CascadeMux I__12061 (
            .O(N__52183),
            .I(n22142_cascade_));
    InMux I__12060 (
            .O(N__52180),
            .I(N__52177));
    LocalMux I__12059 (
            .O(N__52177),
            .I(N__52174));
    Span4Mux_v I__12058 (
            .O(N__52174),
            .I(N__52171));
    Sp12to4 I__12057 (
            .O(N__52171),
            .I(N__52168));
    Span12Mux_h I__12056 (
            .O(N__52168),
            .I(N__52165));
    Odrv12 I__12055 (
            .O(N__52165),
            .I(n22137));
    CascadeMux I__12054 (
            .O(N__52162),
            .I(n23408_cascade_));
    CascadeMux I__12053 (
            .O(N__52159),
            .I(n23411_cascade_));
    InMux I__12052 (
            .O(N__52156),
            .I(N__52153));
    LocalMux I__12051 (
            .O(N__52153),
            .I(N__52150));
    Odrv12 I__12050 (
            .O(N__52150),
            .I(n111_adj_1754));
    CascadeMux I__12049 (
            .O(N__52147),
            .I(comm_buf_1_7_N_559_1_cascade_));
    InMux I__12048 (
            .O(N__52144),
            .I(N__52139));
    InMux I__12047 (
            .O(N__52143),
            .I(N__52135));
    CascadeMux I__12046 (
            .O(N__52142),
            .I(N__52131));
    LocalMux I__12045 (
            .O(N__52139),
            .I(N__52128));
    InMux I__12044 (
            .O(N__52138),
            .I(N__52125));
    LocalMux I__12043 (
            .O(N__52135),
            .I(N__52122));
    CascadeMux I__12042 (
            .O(N__52134),
            .I(N__52118));
    InMux I__12041 (
            .O(N__52131),
            .I(N__52115));
    Span4Mux_v I__12040 (
            .O(N__52128),
            .I(N__52108));
    LocalMux I__12039 (
            .O(N__52125),
            .I(N__52108));
    Span4Mux_v I__12038 (
            .O(N__52122),
            .I(N__52108));
    InMux I__12037 (
            .O(N__52121),
            .I(N__52104));
    InMux I__12036 (
            .O(N__52118),
            .I(N__52101));
    LocalMux I__12035 (
            .O(N__52115),
            .I(N__52098));
    Span4Mux_v I__12034 (
            .O(N__52108),
            .I(N__52095));
    InMux I__12033 (
            .O(N__52107),
            .I(N__52092));
    LocalMux I__12032 (
            .O(N__52104),
            .I(N__52087));
    LocalMux I__12031 (
            .O(N__52101),
            .I(N__52084));
    Span4Mux_v I__12030 (
            .O(N__52098),
            .I(N__52077));
    Span4Mux_h I__12029 (
            .O(N__52095),
            .I(N__52077));
    LocalMux I__12028 (
            .O(N__52092),
            .I(N__52077));
    InMux I__12027 (
            .O(N__52091),
            .I(N__52072));
    InMux I__12026 (
            .O(N__52090),
            .I(N__52072));
    Span4Mux_v I__12025 (
            .O(N__52087),
            .I(N__52069));
    Sp12to4 I__12024 (
            .O(N__52084),
            .I(N__52066));
    Span4Mux_h I__12023 (
            .O(N__52077),
            .I(N__52063));
    LocalMux I__12022 (
            .O(N__52072),
            .I(N__52060));
    Span4Mux_h I__12021 (
            .O(N__52069),
            .I(N__52057));
    Span12Mux_v I__12020 (
            .O(N__52066),
            .I(N__52054));
    Span4Mux_h I__12019 (
            .O(N__52063),
            .I(N__52051));
    Span12Mux_h I__12018 (
            .O(N__52060),
            .I(N__52048));
    Odrv4 I__12017 (
            .O(N__52057),
            .I(comm_buf_1_1));
    Odrv12 I__12016 (
            .O(N__52054),
            .I(comm_buf_1_1));
    Odrv4 I__12015 (
            .O(N__52051),
            .I(comm_buf_1_1));
    Odrv12 I__12014 (
            .O(N__52048),
            .I(comm_buf_1_1));
    InMux I__12013 (
            .O(N__52039),
            .I(N__52036));
    LocalMux I__12012 (
            .O(N__52036),
            .I(N__52033));
    Span4Mux_h I__12011 (
            .O(N__52033),
            .I(N__52030));
    Span4Mux_v I__12010 (
            .O(N__52030),
            .I(N__52027));
    Odrv4 I__12009 (
            .O(N__52027),
            .I(buf_data_iac_9));
    CascadeMux I__12008 (
            .O(N__52024),
            .I(N__52021));
    InMux I__12007 (
            .O(N__52021),
            .I(N__52018));
    LocalMux I__12006 (
            .O(N__52018),
            .I(n26_adj_1753));
    InMux I__12005 (
            .O(N__52015),
            .I(N__52012));
    LocalMux I__12004 (
            .O(N__52012),
            .I(n22143));
    CascadeMux I__12003 (
            .O(N__52009),
            .I(n37_cascade_));
    CascadeMux I__12002 (
            .O(N__52006),
            .I(n12761_cascade_));
    InMux I__12001 (
            .O(N__52003),
            .I(N__52000));
    LocalMux I__12000 (
            .O(N__52000),
            .I(N__51996));
    InMux I__11999 (
            .O(N__51999),
            .I(N__51993));
    Span4Mux_v I__11998 (
            .O(N__51996),
            .I(N__51990));
    LocalMux I__11997 (
            .O(N__51993),
            .I(data_idxvec_5));
    Odrv4 I__11996 (
            .O(N__51990),
            .I(data_idxvec_5));
    InMux I__11995 (
            .O(N__51985),
            .I(N__51982));
    LocalMux I__11994 (
            .O(N__51982),
            .I(N__51977));
    InMux I__11993 (
            .O(N__51981),
            .I(N__51974));
    InMux I__11992 (
            .O(N__51980),
            .I(N__51971));
    Span4Mux_h I__11991 (
            .O(N__51977),
            .I(N__51968));
    LocalMux I__11990 (
            .O(N__51974),
            .I(N__51965));
    LocalMux I__11989 (
            .O(N__51971),
            .I(data_cntvec_5));
    Odrv4 I__11988 (
            .O(N__51968),
            .I(data_cntvec_5));
    Odrv4 I__11987 (
            .O(N__51965),
            .I(data_cntvec_5));
    CascadeMux I__11986 (
            .O(N__51958),
            .I(n26_adj_1730_cascade_));
    InMux I__11985 (
            .O(N__51955),
            .I(N__51952));
    LocalMux I__11984 (
            .O(N__51952),
            .I(N__51949));
    Span4Mux_v I__11983 (
            .O(N__51949),
            .I(N__51945));
    CascadeMux I__11982 (
            .O(N__51948),
            .I(N__51941));
    Span4Mux_h I__11981 (
            .O(N__51945),
            .I(N__51938));
    InMux I__11980 (
            .O(N__51944),
            .I(N__51933));
    InMux I__11979 (
            .O(N__51941),
            .I(N__51933));
    Odrv4 I__11978 (
            .O(N__51938),
            .I(req_data_cnt_5));
    LocalMux I__11977 (
            .O(N__51933),
            .I(req_data_cnt_5));
    CascadeMux I__11976 (
            .O(N__51928),
            .I(n23336_cascade_));
    CascadeMux I__11975 (
            .O(N__51925),
            .I(N__51921));
    InMux I__11974 (
            .O(N__51924),
            .I(N__51918));
    InMux I__11973 (
            .O(N__51921),
            .I(N__51914));
    LocalMux I__11972 (
            .O(N__51918),
            .I(N__51911));
    InMux I__11971 (
            .O(N__51917),
            .I(N__51908));
    LocalMux I__11970 (
            .O(N__51914),
            .I(acadc_skipCount_5));
    Odrv4 I__11969 (
            .O(N__51911),
            .I(acadc_skipCount_5));
    LocalMux I__11968 (
            .O(N__51908),
            .I(acadc_skipCount_5));
    CascadeMux I__11967 (
            .O(N__51901),
            .I(n23339_cascade_));
    CascadeMux I__11966 (
            .O(N__51898),
            .I(n30_adj_1731_cascade_));
    InMux I__11965 (
            .O(N__51895),
            .I(N__51892));
    LocalMux I__11964 (
            .O(N__51892),
            .I(N__51889));
    Span4Mux_v I__11963 (
            .O(N__51889),
            .I(N__51886));
    Span4Mux_h I__11962 (
            .O(N__51886),
            .I(N__51883));
    Span4Mux_h I__11961 (
            .O(N__51883),
            .I(N__51880));
    Odrv4 I__11960 (
            .O(N__51880),
            .I(n111_adj_1732));
    InMux I__11959 (
            .O(N__51877),
            .I(N__51874));
    LocalMux I__11958 (
            .O(N__51874),
            .I(N__51871));
    Span4Mux_h I__11957 (
            .O(N__51871),
            .I(N__51868));
    Odrv4 I__11956 (
            .O(N__51868),
            .I(n22354));
    CascadeMux I__11955 (
            .O(N__51865),
            .I(N__51862));
    InMux I__11954 (
            .O(N__51862),
            .I(N__51859));
    LocalMux I__11953 (
            .O(N__51859),
            .I(n22353));
    InMux I__11952 (
            .O(N__51856),
            .I(N__51853));
    LocalMux I__11951 (
            .O(N__51853),
            .I(N__51850));
    Span4Mux_h I__11950 (
            .O(N__51850),
            .I(N__51847));
    Odrv4 I__11949 (
            .O(N__51847),
            .I(comm_length_1));
    InMux I__11948 (
            .O(N__51844),
            .I(N__51841));
    LocalMux I__11947 (
            .O(N__51841),
            .I(n4_adj_1745));
    InMux I__11946 (
            .O(N__51838),
            .I(N__51834));
    InMux I__11945 (
            .O(N__51837),
            .I(N__51831));
    LocalMux I__11944 (
            .O(N__51834),
            .I(N__51824));
    LocalMux I__11943 (
            .O(N__51831),
            .I(N__51824));
    InMux I__11942 (
            .O(N__51830),
            .I(N__51818));
    InMux I__11941 (
            .O(N__51829),
            .I(N__51815));
    Span4Mux_v I__11940 (
            .O(N__51824),
            .I(N__51812));
    InMux I__11939 (
            .O(N__51823),
            .I(N__51809));
    InMux I__11938 (
            .O(N__51822),
            .I(N__51804));
    InMux I__11937 (
            .O(N__51821),
            .I(N__51801));
    LocalMux I__11936 (
            .O(N__51818),
            .I(N__51797));
    LocalMux I__11935 (
            .O(N__51815),
            .I(N__51792));
    Span4Mux_h I__11934 (
            .O(N__51812),
            .I(N__51792));
    LocalMux I__11933 (
            .O(N__51809),
            .I(N__51789));
    CascadeMux I__11932 (
            .O(N__51808),
            .I(N__51786));
    InMux I__11931 (
            .O(N__51807),
            .I(N__51781));
    LocalMux I__11930 (
            .O(N__51804),
            .I(N__51774));
    LocalMux I__11929 (
            .O(N__51801),
            .I(N__51774));
    InMux I__11928 (
            .O(N__51800),
            .I(N__51771));
    Span4Mux_h I__11927 (
            .O(N__51797),
            .I(N__51768));
    Span4Mux_v I__11926 (
            .O(N__51792),
            .I(N__51765));
    Span4Mux_h I__11925 (
            .O(N__51789),
            .I(N__51762));
    InMux I__11924 (
            .O(N__51786),
            .I(N__51755));
    InMux I__11923 (
            .O(N__51785),
            .I(N__51755));
    InMux I__11922 (
            .O(N__51784),
            .I(N__51755));
    LocalMux I__11921 (
            .O(N__51781),
            .I(N__51752));
    InMux I__11920 (
            .O(N__51780),
            .I(N__51747));
    InMux I__11919 (
            .O(N__51779),
            .I(N__51747));
    Odrv12 I__11918 (
            .O(N__51774),
            .I(comm_index_1));
    LocalMux I__11917 (
            .O(N__51771),
            .I(comm_index_1));
    Odrv4 I__11916 (
            .O(N__51768),
            .I(comm_index_1));
    Odrv4 I__11915 (
            .O(N__51765),
            .I(comm_index_1));
    Odrv4 I__11914 (
            .O(N__51762),
            .I(comm_index_1));
    LocalMux I__11913 (
            .O(N__51755),
            .I(comm_index_1));
    Odrv4 I__11912 (
            .O(N__51752),
            .I(comm_index_1));
    LocalMux I__11911 (
            .O(N__51747),
            .I(comm_index_1));
    InMux I__11910 (
            .O(N__51730),
            .I(N__51726));
    CascadeMux I__11909 (
            .O(N__51729),
            .I(N__51722));
    LocalMux I__11908 (
            .O(N__51726),
            .I(N__51719));
    InMux I__11907 (
            .O(N__51725),
            .I(N__51716));
    InMux I__11906 (
            .O(N__51722),
            .I(N__51713));
    Span4Mux_h I__11905 (
            .O(N__51719),
            .I(N__51708));
    LocalMux I__11904 (
            .O(N__51716),
            .I(N__51708));
    LocalMux I__11903 (
            .O(N__51713),
            .I(req_data_cnt_14));
    Odrv4 I__11902 (
            .O(N__51708),
            .I(req_data_cnt_14));
    InMux I__11901 (
            .O(N__51703),
            .I(N__51700));
    LocalMux I__11900 (
            .O(N__51700),
            .I(N__51696));
    InMux I__11899 (
            .O(N__51699),
            .I(N__51693));
    Span4Mux_v I__11898 (
            .O(N__51696),
            .I(N__51690));
    LocalMux I__11897 (
            .O(N__51693),
            .I(data_cntvec_14));
    Odrv4 I__11896 (
            .O(N__51690),
            .I(data_cntvec_14));
    InMux I__11895 (
            .O(N__51685),
            .I(N__51682));
    LocalMux I__11894 (
            .O(N__51682),
            .I(N__51679));
    Span4Mux_h I__11893 (
            .O(N__51679),
            .I(N__51676));
    Span4Mux_h I__11892 (
            .O(N__51676),
            .I(N__51673));
    Odrv4 I__11891 (
            .O(N__51673),
            .I(n23));
    InMux I__11890 (
            .O(N__51670),
            .I(N__51667));
    LocalMux I__11889 (
            .O(N__51667),
            .I(n111));
    InMux I__11888 (
            .O(N__51664),
            .I(N__51661));
    LocalMux I__11887 (
            .O(N__51661),
            .I(N__51658));
    Odrv4 I__11886 (
            .O(N__51658),
            .I(n30_adj_1579));
    InMux I__11885 (
            .O(N__51655),
            .I(N__51652));
    LocalMux I__11884 (
            .O(N__51652),
            .I(N__51649));
    Odrv4 I__11883 (
            .O(N__51649),
            .I(comm_buf_1_7_N_559_0));
    SRMux I__11882 (
            .O(N__51646),
            .I(N__51642));
    SRMux I__11881 (
            .O(N__51645),
            .I(N__51639));
    LocalMux I__11880 (
            .O(N__51642),
            .I(N__51636));
    LocalMux I__11879 (
            .O(N__51639),
            .I(N__51633));
    Span4Mux_v I__11878 (
            .O(N__51636),
            .I(N__51630));
    Odrv4 I__11877 (
            .O(N__51633),
            .I(n21271));
    Odrv4 I__11876 (
            .O(N__51630),
            .I(n21271));
    InMux I__11875 (
            .O(N__51625),
            .I(N__51620));
    InMux I__11874 (
            .O(N__51624),
            .I(N__51615));
    InMux I__11873 (
            .O(N__51623),
            .I(N__51615));
    LocalMux I__11872 (
            .O(N__51620),
            .I(N__51609));
    LocalMux I__11871 (
            .O(N__51615),
            .I(N__51609));
    InMux I__11870 (
            .O(N__51614),
            .I(N__51606));
    Odrv12 I__11869 (
            .O(N__51609),
            .I(n11258));
    LocalMux I__11868 (
            .O(N__51606),
            .I(n11258));
    CascadeMux I__11867 (
            .O(N__51601),
            .I(N__51598));
    InMux I__11866 (
            .O(N__51598),
            .I(N__51595));
    LocalMux I__11865 (
            .O(N__51595),
            .I(N__51592));
    Odrv4 I__11864 (
            .O(N__51592),
            .I(n22089));
    InMux I__11863 (
            .O(N__51589),
            .I(N__51586));
    LocalMux I__11862 (
            .O(N__51586),
            .I(N__51582));
    InMux I__11861 (
            .O(N__51585),
            .I(N__51579));
    Odrv4 I__11860 (
            .O(N__51582),
            .I(n20318));
    LocalMux I__11859 (
            .O(N__51579),
            .I(n20318));
    CascadeMux I__11858 (
            .O(N__51574),
            .I(n12_adj_1677_cascade_));
    CascadeMux I__11857 (
            .O(N__51571),
            .I(n12892_cascade_));
    InMux I__11856 (
            .O(N__51568),
            .I(N__51563));
    InMux I__11855 (
            .O(N__51567),
            .I(N__51560));
    InMux I__11854 (
            .O(N__51566),
            .I(N__51557));
    LocalMux I__11853 (
            .O(N__51563),
            .I(N__51554));
    LocalMux I__11852 (
            .O(N__51560),
            .I(n12951));
    LocalMux I__11851 (
            .O(N__51557),
            .I(n12951));
    Odrv4 I__11850 (
            .O(N__51554),
            .I(n12951));
    CascadeMux I__11849 (
            .O(N__51547),
            .I(N__51543));
    CascadeMux I__11848 (
            .O(N__51546),
            .I(N__51539));
    InMux I__11847 (
            .O(N__51543),
            .I(N__51536));
    InMux I__11846 (
            .O(N__51542),
            .I(N__51531));
    InMux I__11845 (
            .O(N__51539),
            .I(N__51531));
    LocalMux I__11844 (
            .O(N__51536),
            .I(N__51528));
    LocalMux I__11843 (
            .O(N__51531),
            .I(N__51525));
    Span12Mux_v I__11842 (
            .O(N__51528),
            .I(N__51522));
    Span12Mux_v I__11841 (
            .O(N__51525),
            .I(N__51519));
    Odrv12 I__11840 (
            .O(N__51522),
            .I(n9714));
    Odrv12 I__11839 (
            .O(N__51519),
            .I(n9714));
    InMux I__11838 (
            .O(N__51514),
            .I(N__51511));
    LocalMux I__11837 (
            .O(N__51511),
            .I(N__51508));
    Span4Mux_h I__11836 (
            .O(N__51508),
            .I(N__51505));
    Odrv4 I__11835 (
            .O(N__51505),
            .I(n11_adj_1585));
    InMux I__11834 (
            .O(N__51502),
            .I(N__51498));
    InMux I__11833 (
            .O(N__51501),
            .I(N__51495));
    LocalMux I__11832 (
            .O(N__51498),
            .I(N__51492));
    LocalMux I__11831 (
            .O(N__51495),
            .I(N__51489));
    Span4Mux_v I__11830 (
            .O(N__51492),
            .I(N__51486));
    Span4Mux_h I__11829 (
            .O(N__51489),
            .I(N__51483));
    Span4Mux_h I__11828 (
            .O(N__51486),
            .I(N__51478));
    Span4Mux_v I__11827 (
            .O(N__51483),
            .I(N__51478));
    Span4Mux_v I__11826 (
            .O(N__51478),
            .I(N__51475));
    Odrv4 I__11825 (
            .O(N__51475),
            .I(n14_adj_1652));
    InMux I__11824 (
            .O(N__51472),
            .I(N__51462));
    InMux I__11823 (
            .O(N__51471),
            .I(N__51462));
    InMux I__11822 (
            .O(N__51470),
            .I(N__51462));
    InMux I__11821 (
            .O(N__51469),
            .I(N__51459));
    LocalMux I__11820 (
            .O(N__51462),
            .I(N__51454));
    LocalMux I__11819 (
            .O(N__51459),
            .I(N__51454));
    Odrv4 I__11818 (
            .O(N__51454),
            .I(\comm_spi.bit_cnt_1 ));
    CascadeMux I__11817 (
            .O(N__51451),
            .I(N__51447));
    InMux I__11816 (
            .O(N__51450),
            .I(N__51441));
    InMux I__11815 (
            .O(N__51447),
            .I(N__51432));
    InMux I__11814 (
            .O(N__51446),
            .I(N__51432));
    InMux I__11813 (
            .O(N__51445),
            .I(N__51432));
    InMux I__11812 (
            .O(N__51444),
            .I(N__51432));
    LocalMux I__11811 (
            .O(N__51441),
            .I(N__51429));
    LocalMux I__11810 (
            .O(N__51432),
            .I(\comm_spi.bit_cnt_0 ));
    Odrv4 I__11809 (
            .O(N__51429),
            .I(\comm_spi.bit_cnt_0 ));
    InMux I__11808 (
            .O(N__51424),
            .I(N__51417));
    InMux I__11807 (
            .O(N__51423),
            .I(N__51417));
    InMux I__11806 (
            .O(N__51422),
            .I(N__51414));
    LocalMux I__11805 (
            .O(N__51417),
            .I(N__51409));
    LocalMux I__11804 (
            .O(N__51414),
            .I(N__51409));
    Odrv4 I__11803 (
            .O(N__51409),
            .I(\comm_spi.bit_cnt_2 ));
    InMux I__11802 (
            .O(N__51406),
            .I(N__51403));
    LocalMux I__11801 (
            .O(N__51403),
            .I(N__51400));
    Odrv4 I__11800 (
            .O(N__51400),
            .I(n22487));
    InMux I__11799 (
            .O(N__51397),
            .I(N__51393));
    InMux I__11798 (
            .O(N__51396),
            .I(N__51390));
    LocalMux I__11797 (
            .O(N__51393),
            .I(N__51387));
    LocalMux I__11796 (
            .O(N__51390),
            .I(N__51384));
    Span4Mux_h I__11795 (
            .O(N__51387),
            .I(N__51381));
    Span12Mux_h I__11794 (
            .O(N__51384),
            .I(N__51377));
    Span4Mux_h I__11793 (
            .O(N__51381),
            .I(N__51374));
    InMux I__11792 (
            .O(N__51380),
            .I(N__51371));
    Odrv12 I__11791 (
            .O(N__51377),
            .I(n21983));
    Odrv4 I__11790 (
            .O(N__51374),
            .I(n21983));
    LocalMux I__11789 (
            .O(N__51371),
            .I(n21983));
    InMux I__11788 (
            .O(N__51364),
            .I(N__51355));
    InMux I__11787 (
            .O(N__51363),
            .I(N__51355));
    InMux I__11786 (
            .O(N__51362),
            .I(N__51349));
    InMux I__11785 (
            .O(N__51361),
            .I(N__51343));
    InMux I__11784 (
            .O(N__51360),
            .I(N__51343));
    LocalMux I__11783 (
            .O(N__51355),
            .I(N__51340));
    InMux I__11782 (
            .O(N__51354),
            .I(N__51331));
    InMux I__11781 (
            .O(N__51353),
            .I(N__51331));
    InMux I__11780 (
            .O(N__51352),
            .I(N__51331));
    LocalMux I__11779 (
            .O(N__51349),
            .I(N__51328));
    InMux I__11778 (
            .O(N__51348),
            .I(N__51325));
    LocalMux I__11777 (
            .O(N__51343),
            .I(N__51320));
    Span4Mux_v I__11776 (
            .O(N__51340),
            .I(N__51317));
    InMux I__11775 (
            .O(N__51339),
            .I(N__51314));
    CascadeMux I__11774 (
            .O(N__51338),
            .I(N__51311));
    LocalMux I__11773 (
            .O(N__51331),
            .I(N__51307));
    Span4Mux_h I__11772 (
            .O(N__51328),
            .I(N__51302));
    LocalMux I__11771 (
            .O(N__51325),
            .I(N__51302));
    InMux I__11770 (
            .O(N__51324),
            .I(N__51299));
    InMux I__11769 (
            .O(N__51323),
            .I(N__51296));
    Span4Mux_v I__11768 (
            .O(N__51320),
            .I(N__51289));
    Span4Mux_h I__11767 (
            .O(N__51317),
            .I(N__51289));
    LocalMux I__11766 (
            .O(N__51314),
            .I(N__51289));
    InMux I__11765 (
            .O(N__51311),
            .I(N__51284));
    InMux I__11764 (
            .O(N__51310),
            .I(N__51284));
    Span4Mux_v I__11763 (
            .O(N__51307),
            .I(N__51280));
    Span4Mux_h I__11762 (
            .O(N__51302),
            .I(N__51277));
    LocalMux I__11761 (
            .O(N__51299),
            .I(N__51268));
    LocalMux I__11760 (
            .O(N__51296),
            .I(N__51268));
    Span4Mux_h I__11759 (
            .O(N__51289),
            .I(N__51268));
    LocalMux I__11758 (
            .O(N__51284),
            .I(N__51268));
    InMux I__11757 (
            .O(N__51283),
            .I(N__51265));
    Span4Mux_h I__11756 (
            .O(N__51280),
            .I(N__51262));
    Span4Mux_h I__11755 (
            .O(N__51277),
            .I(N__51259));
    Span4Mux_v I__11754 (
            .O(N__51268),
            .I(N__51256));
    LocalMux I__11753 (
            .O(N__51265),
            .I(n13171));
    Odrv4 I__11752 (
            .O(N__51262),
            .I(n13171));
    Odrv4 I__11751 (
            .O(N__51259),
            .I(n13171));
    Odrv4 I__11750 (
            .O(N__51256),
            .I(n13171));
    CascadeMux I__11749 (
            .O(N__51247),
            .I(n13171_cascade_));
    InMux I__11748 (
            .O(N__51244),
            .I(N__51241));
    LocalMux I__11747 (
            .O(N__51241),
            .I(n22033));
    CascadeMux I__11746 (
            .O(N__51238),
            .I(n12064_cascade_));
    CEMux I__11745 (
            .O(N__51235),
            .I(N__51232));
    LocalMux I__11744 (
            .O(N__51232),
            .I(n21885));
    CascadeMux I__11743 (
            .O(N__51229),
            .I(n22073_cascade_));
    SRMux I__11742 (
            .O(N__51226),
            .I(N__51220));
    SRMux I__11741 (
            .O(N__51225),
            .I(N__51216));
    SRMux I__11740 (
            .O(N__51224),
            .I(N__51213));
    SRMux I__11739 (
            .O(N__51223),
            .I(N__51210));
    LocalMux I__11738 (
            .O(N__51220),
            .I(N__51207));
    SRMux I__11737 (
            .O(N__51219),
            .I(N__51204));
    LocalMux I__11736 (
            .O(N__51216),
            .I(N__51197));
    LocalMux I__11735 (
            .O(N__51213),
            .I(N__51197));
    LocalMux I__11734 (
            .O(N__51210),
            .I(N__51197));
    Span4Mux_v I__11733 (
            .O(N__51207),
            .I(N__51192));
    LocalMux I__11732 (
            .O(N__51204),
            .I(N__51192));
    Span4Mux_v I__11731 (
            .O(N__51197),
            .I(N__51189));
    Odrv4 I__11730 (
            .O(N__51192),
            .I(flagcntwd));
    Odrv4 I__11729 (
            .O(N__51189),
            .I(flagcntwd));
    CEMux I__11728 (
            .O(N__51184),
            .I(N__51181));
    LocalMux I__11727 (
            .O(N__51181),
            .I(N__51178));
    Odrv4 I__11726 (
            .O(N__51178),
            .I(n12050));
    InMux I__11725 (
            .O(N__51175),
            .I(N__51172));
    LocalMux I__11724 (
            .O(N__51172),
            .I(n10_adj_1602));
    InMux I__11723 (
            .O(N__51169),
            .I(N__51161));
    InMux I__11722 (
            .O(N__51168),
            .I(N__51158));
    InMux I__11721 (
            .O(N__51167),
            .I(N__51153));
    InMux I__11720 (
            .O(N__51166),
            .I(N__51153));
    InMux I__11719 (
            .O(N__51165),
            .I(N__51148));
    InMux I__11718 (
            .O(N__51164),
            .I(N__51148));
    LocalMux I__11717 (
            .O(N__51161),
            .I(N__51141));
    LocalMux I__11716 (
            .O(N__51158),
            .I(N__51141));
    LocalMux I__11715 (
            .O(N__51153),
            .I(N__51141));
    LocalMux I__11714 (
            .O(N__51148),
            .I(N__51136));
    Span4Mux_v I__11713 (
            .O(N__51141),
            .I(N__51136));
    Odrv4 I__11712 (
            .O(N__51136),
            .I(comm_cmd_7));
    CascadeMux I__11711 (
            .O(N__51133),
            .I(N__51130));
    InMux I__11710 (
            .O(N__51130),
            .I(N__51127));
    LocalMux I__11709 (
            .O(N__51127),
            .I(n29));
    InMux I__11708 (
            .O(N__51124),
            .I(N__51121));
    LocalMux I__11707 (
            .O(N__51121),
            .I(N__51118));
    Span4Mux_v I__11706 (
            .O(N__51118),
            .I(N__51115));
    Span4Mux_h I__11705 (
            .O(N__51115),
            .I(N__51111));
    InMux I__11704 (
            .O(N__51114),
            .I(N__51108));
    Odrv4 I__11703 (
            .O(N__51111),
            .I(\comm_spi.n24034 ));
    LocalMux I__11702 (
            .O(N__51108),
            .I(\comm_spi.n24034 ));
    InMux I__11701 (
            .O(N__51103),
            .I(N__51100));
    LocalMux I__11700 (
            .O(N__51100),
            .I(N__51097));
    Span4Mux_h I__11699 (
            .O(N__51097),
            .I(N__51094));
    Span4Mux_h I__11698 (
            .O(N__51094),
            .I(N__51090));
    InMux I__11697 (
            .O(N__51093),
            .I(N__51087));
    Sp12to4 I__11696 (
            .O(N__51090),
            .I(N__51082));
    LocalMux I__11695 (
            .O(N__51087),
            .I(N__51082));
    Odrv12 I__11694 (
            .O(N__51082),
            .I(\comm_spi.n15352 ));
    InMux I__11693 (
            .O(N__51079),
            .I(N__51076));
    LocalMux I__11692 (
            .O(N__51076),
            .I(N__51072));
    InMux I__11691 (
            .O(N__51075),
            .I(N__51069));
    Span4Mux_h I__11690 (
            .O(N__51072),
            .I(N__51066));
    LocalMux I__11689 (
            .O(N__51069),
            .I(N__51063));
    Span4Mux_h I__11688 (
            .O(N__51066),
            .I(N__51060));
    Span4Mux_v I__11687 (
            .O(N__51063),
            .I(N__51057));
    Odrv4 I__11686 (
            .O(N__51060),
            .I(\comm_spi.n15353 ));
    Odrv4 I__11685 (
            .O(N__51057),
            .I(\comm_spi.n15353 ));
    InMux I__11684 (
            .O(N__51052),
            .I(N__51049));
    LocalMux I__11683 (
            .O(N__51049),
            .I(N__51046));
    Span4Mux_v I__11682 (
            .O(N__51046),
            .I(N__51042));
    InMux I__11681 (
            .O(N__51045),
            .I(N__51039));
    Span4Mux_v I__11680 (
            .O(N__51042),
            .I(N__51036));
    LocalMux I__11679 (
            .O(N__51039),
            .I(N__51033));
    Span4Mux_h I__11678 (
            .O(N__51036),
            .I(N__51028));
    Span4Mux_h I__11677 (
            .O(N__51033),
            .I(N__51028));
    Span4Mux_h I__11676 (
            .O(N__51028),
            .I(N__51025));
    Odrv4 I__11675 (
            .O(N__51025),
            .I(\comm_spi.n15357 ));
    SRMux I__11674 (
            .O(N__51022),
            .I(N__51019));
    LocalMux I__11673 (
            .O(N__51019),
            .I(N__51016));
    Span4Mux_v I__11672 (
            .O(N__51016),
            .I(N__51013));
    Span4Mux_h I__11671 (
            .O(N__51013),
            .I(N__51010));
    Span4Mux_v I__11670 (
            .O(N__51010),
            .I(N__51007));
    Odrv4 I__11669 (
            .O(N__51007),
            .I(\comm_spi.data_tx_7__N_874 ));
    CascadeMux I__11668 (
            .O(N__51004),
            .I(n22489_cascade_));
    CascadeMux I__11667 (
            .O(N__51001),
            .I(n20959_cascade_));
    CEMux I__11666 (
            .O(N__50998),
            .I(N__50995));
    LocalMux I__11665 (
            .O(N__50995),
            .I(n21883));
    InMux I__11664 (
            .O(N__50992),
            .I(N__50989));
    LocalMux I__11663 (
            .O(N__50989),
            .I(n19241));
    InMux I__11662 (
            .O(N__50986),
            .I(N__50983));
    LocalMux I__11661 (
            .O(N__50983),
            .I(N__50980));
    Odrv12 I__11660 (
            .O(N__50980),
            .I(n22177));
    InMux I__11659 (
            .O(N__50977),
            .I(N__50974));
    LocalMux I__11658 (
            .O(N__50974),
            .I(N__50971));
    Odrv12 I__11657 (
            .O(N__50971),
            .I(n22180));
    CascadeMux I__11656 (
            .O(N__50968),
            .I(n23462_cascade_));
    InMux I__11655 (
            .O(N__50965),
            .I(N__50962));
    LocalMux I__11654 (
            .O(N__50962),
            .I(N__50959));
    Span4Mux_h I__11653 (
            .O(N__50959),
            .I(N__50956));
    Odrv4 I__11652 (
            .O(N__50956),
            .I(n23465));
    CascadeMux I__11651 (
            .O(N__50953),
            .I(N__50950));
    InMux I__11650 (
            .O(N__50950),
            .I(N__50946));
    InMux I__11649 (
            .O(N__50949),
            .I(N__50943));
    LocalMux I__11648 (
            .O(N__50946),
            .I(data_idxvec_9));
    LocalMux I__11647 (
            .O(N__50943),
            .I(data_idxvec_9));
    InMux I__11646 (
            .O(N__50938),
            .I(N__50934));
    InMux I__11645 (
            .O(N__50937),
            .I(N__50930));
    LocalMux I__11644 (
            .O(N__50934),
            .I(N__50927));
    InMux I__11643 (
            .O(N__50933),
            .I(N__50924));
    LocalMux I__11642 (
            .O(N__50930),
            .I(data_cntvec_9));
    Odrv4 I__11641 (
            .O(N__50927),
            .I(data_cntvec_9));
    LocalMux I__11640 (
            .O(N__50924),
            .I(data_cntvec_9));
    InMux I__11639 (
            .O(N__50917),
            .I(N__50914));
    LocalMux I__11638 (
            .O(N__50914),
            .I(N__50911));
    Span4Mux_v I__11637 (
            .O(N__50911),
            .I(N__50908));
    Span4Mux_h I__11636 (
            .O(N__50908),
            .I(N__50905));
    Odrv4 I__11635 (
            .O(N__50905),
            .I(buf_data_iac_17));
    CascadeMux I__11634 (
            .O(N__50902),
            .I(n22184_cascade_));
    InMux I__11633 (
            .O(N__50899),
            .I(N__50896));
    LocalMux I__11632 (
            .O(N__50896),
            .I(n22186));
    InMux I__11631 (
            .O(N__50893),
            .I(N__50880));
    InMux I__11630 (
            .O(N__50892),
            .I(N__50880));
    InMux I__11629 (
            .O(N__50891),
            .I(N__50877));
    InMux I__11628 (
            .O(N__50890),
            .I(N__50872));
    InMux I__11627 (
            .O(N__50889),
            .I(N__50872));
    InMux I__11626 (
            .O(N__50888),
            .I(N__50865));
    InMux I__11625 (
            .O(N__50887),
            .I(N__50865));
    InMux I__11624 (
            .O(N__50886),
            .I(N__50865));
    CascadeMux I__11623 (
            .O(N__50885),
            .I(N__50862));
    LocalMux I__11622 (
            .O(N__50880),
            .I(N__50859));
    LocalMux I__11621 (
            .O(N__50877),
            .I(N__50853));
    LocalMux I__11620 (
            .O(N__50872),
            .I(N__50853));
    LocalMux I__11619 (
            .O(N__50865),
            .I(N__50850));
    InMux I__11618 (
            .O(N__50862),
            .I(N__50847));
    Span4Mux_h I__11617 (
            .O(N__50859),
            .I(N__50844));
    InMux I__11616 (
            .O(N__50858),
            .I(N__50841));
    Span4Mux_v I__11615 (
            .O(N__50853),
            .I(N__50836));
    Span4Mux_h I__11614 (
            .O(N__50850),
            .I(N__50836));
    LocalMux I__11613 (
            .O(N__50847),
            .I(N__50833));
    Span4Mux_h I__11612 (
            .O(N__50844),
            .I(N__50828));
    LocalMux I__11611 (
            .O(N__50841),
            .I(N__50828));
    Span4Mux_h I__11610 (
            .O(N__50836),
            .I(N__50825));
    Span12Mux_s11_h I__11609 (
            .O(N__50833),
            .I(N__50820));
    Sp12to4 I__11608 (
            .O(N__50828),
            .I(N__50820));
    Odrv4 I__11607 (
            .O(N__50825),
            .I(n21997));
    Odrv12 I__11606 (
            .O(N__50820),
            .I(n21997));
    InMux I__11605 (
            .O(N__50815),
            .I(N__50809));
    InMux I__11604 (
            .O(N__50814),
            .I(N__50809));
    LocalMux I__11603 (
            .O(N__50809),
            .I(N__50804));
    InMux I__11602 (
            .O(N__50808),
            .I(N__50801));
    InMux I__11601 (
            .O(N__50807),
            .I(N__50798));
    Span4Mux_v I__11600 (
            .O(N__50804),
            .I(N__50794));
    LocalMux I__11599 (
            .O(N__50801),
            .I(N__50791));
    LocalMux I__11598 (
            .O(N__50798),
            .I(N__50788));
    InMux I__11597 (
            .O(N__50797),
            .I(N__50785));
    Odrv4 I__11596 (
            .O(N__50794),
            .I(n14_adj_1656));
    Odrv12 I__11595 (
            .O(N__50791),
            .I(n14_adj_1656));
    Odrv4 I__11594 (
            .O(N__50788),
            .I(n14_adj_1656));
    LocalMux I__11593 (
            .O(N__50785),
            .I(n14_adj_1656));
    InMux I__11592 (
            .O(N__50776),
            .I(N__50772));
    InMux I__11591 (
            .O(N__50775),
            .I(N__50765));
    LocalMux I__11590 (
            .O(N__50772),
            .I(N__50760));
    InMux I__11589 (
            .O(N__50771),
            .I(N__50755));
    InMux I__11588 (
            .O(N__50770),
            .I(N__50755));
    InMux I__11587 (
            .O(N__50769),
            .I(N__50748));
    InMux I__11586 (
            .O(N__50768),
            .I(N__50748));
    LocalMux I__11585 (
            .O(N__50765),
            .I(N__50745));
    InMux I__11584 (
            .O(N__50764),
            .I(N__50742));
    InMux I__11583 (
            .O(N__50763),
            .I(N__50739));
    Span4Mux_v I__11582 (
            .O(N__50760),
            .I(N__50733));
    LocalMux I__11581 (
            .O(N__50755),
            .I(N__50730));
    InMux I__11580 (
            .O(N__50754),
            .I(N__50727));
    InMux I__11579 (
            .O(N__50753),
            .I(N__50724));
    LocalMux I__11578 (
            .O(N__50748),
            .I(N__50719));
    Span4Mux_v I__11577 (
            .O(N__50745),
            .I(N__50716));
    LocalMux I__11576 (
            .O(N__50742),
            .I(N__50711));
    LocalMux I__11575 (
            .O(N__50739),
            .I(N__50711));
    InMux I__11574 (
            .O(N__50738),
            .I(N__50704));
    InMux I__11573 (
            .O(N__50737),
            .I(N__50704));
    InMux I__11572 (
            .O(N__50736),
            .I(N__50704));
    Span4Mux_h I__11571 (
            .O(N__50733),
            .I(N__50697));
    Span4Mux_v I__11570 (
            .O(N__50730),
            .I(N__50697));
    LocalMux I__11569 (
            .O(N__50727),
            .I(N__50697));
    LocalMux I__11568 (
            .O(N__50724),
            .I(N__50694));
    InMux I__11567 (
            .O(N__50723),
            .I(N__50689));
    InMux I__11566 (
            .O(N__50722),
            .I(N__50689));
    Span4Mux_v I__11565 (
            .O(N__50719),
            .I(N__50685));
    Span4Mux_h I__11564 (
            .O(N__50716),
            .I(N__50682));
    Span4Mux_v I__11563 (
            .O(N__50711),
            .I(N__50679));
    LocalMux I__11562 (
            .O(N__50704),
            .I(N__50676));
    Span4Mux_v I__11561 (
            .O(N__50697),
            .I(N__50669));
    Span4Mux_h I__11560 (
            .O(N__50694),
            .I(N__50669));
    LocalMux I__11559 (
            .O(N__50689),
            .I(N__50669));
    InMux I__11558 (
            .O(N__50688),
            .I(N__50666));
    Span4Mux_h I__11557 (
            .O(N__50685),
            .I(N__50659));
    Span4Mux_v I__11556 (
            .O(N__50682),
            .I(N__50659));
    Span4Mux_h I__11555 (
            .O(N__50679),
            .I(N__50659));
    Span12Mux_v I__11554 (
            .O(N__50676),
            .I(N__50656));
    Span4Mux_v I__11553 (
            .O(N__50669),
            .I(N__50653));
    LocalMux I__11552 (
            .O(N__50666),
            .I(n13093));
    Odrv4 I__11551 (
            .O(N__50659),
            .I(n13093));
    Odrv12 I__11550 (
            .O(N__50656),
            .I(n13093));
    Odrv4 I__11549 (
            .O(N__50653),
            .I(n13093));
    CascadeMux I__11548 (
            .O(N__50644),
            .I(N__50641));
    InMux I__11547 (
            .O(N__50641),
            .I(N__50637));
    InMux I__11546 (
            .O(N__50640),
            .I(N__50634));
    LocalMux I__11545 (
            .O(N__50637),
            .I(N__50630));
    LocalMux I__11544 (
            .O(N__50634),
            .I(N__50627));
    InMux I__11543 (
            .O(N__50633),
            .I(N__50624));
    Span12Mux_h I__11542 (
            .O(N__50630),
            .I(N__50621));
    Odrv12 I__11541 (
            .O(N__50627),
            .I(buf_dds0_9));
    LocalMux I__11540 (
            .O(N__50624),
            .I(buf_dds0_9));
    Odrv12 I__11539 (
            .O(N__50621),
            .I(buf_dds0_9));
    InMux I__11538 (
            .O(N__50614),
            .I(N__50611));
    LocalMux I__11537 (
            .O(N__50611),
            .I(N__50605));
    InMux I__11536 (
            .O(N__50610),
            .I(N__50600));
    InMux I__11535 (
            .O(N__50609),
            .I(N__50600));
    InMux I__11534 (
            .O(N__50608),
            .I(N__50596));
    Span4Mux_h I__11533 (
            .O(N__50605),
            .I(N__50587));
    LocalMux I__11532 (
            .O(N__50600),
            .I(N__50587));
    InMux I__11531 (
            .O(N__50599),
            .I(N__50584));
    LocalMux I__11530 (
            .O(N__50596),
            .I(N__50581));
    InMux I__11529 (
            .O(N__50595),
            .I(N__50578));
    InMux I__11528 (
            .O(N__50594),
            .I(N__50573));
    InMux I__11527 (
            .O(N__50593),
            .I(N__50573));
    InMux I__11526 (
            .O(N__50592),
            .I(N__50570));
    Span4Mux_h I__11525 (
            .O(N__50587),
            .I(N__50567));
    LocalMux I__11524 (
            .O(N__50584),
            .I(dds_state_0));
    Odrv4 I__11523 (
            .O(N__50581),
            .I(dds_state_0));
    LocalMux I__11522 (
            .O(N__50578),
            .I(dds_state_0));
    LocalMux I__11521 (
            .O(N__50573),
            .I(dds_state_0));
    LocalMux I__11520 (
            .O(N__50570),
            .I(dds_state_0));
    Odrv4 I__11519 (
            .O(N__50567),
            .I(dds_state_0));
    InMux I__11518 (
            .O(N__50554),
            .I(N__50532));
    InMux I__11517 (
            .O(N__50553),
            .I(N__50521));
    InMux I__11516 (
            .O(N__50552),
            .I(N__50521));
    InMux I__11515 (
            .O(N__50551),
            .I(N__50521));
    InMux I__11514 (
            .O(N__50550),
            .I(N__50521));
    InMux I__11513 (
            .O(N__50549),
            .I(N__50521));
    InMux I__11512 (
            .O(N__50548),
            .I(N__50510));
    InMux I__11511 (
            .O(N__50547),
            .I(N__50510));
    InMux I__11510 (
            .O(N__50546),
            .I(N__50510));
    InMux I__11509 (
            .O(N__50545),
            .I(N__50510));
    InMux I__11508 (
            .O(N__50544),
            .I(N__50510));
    InMux I__11507 (
            .O(N__50543),
            .I(N__50507));
    InMux I__11506 (
            .O(N__50542),
            .I(N__50498));
    InMux I__11505 (
            .O(N__50541),
            .I(N__50498));
    InMux I__11504 (
            .O(N__50540),
            .I(N__50498));
    InMux I__11503 (
            .O(N__50539),
            .I(N__50498));
    InMux I__11502 (
            .O(N__50538),
            .I(N__50495));
    InMux I__11501 (
            .O(N__50537),
            .I(N__50492));
    InMux I__11500 (
            .O(N__50536),
            .I(N__50485));
    InMux I__11499 (
            .O(N__50535),
            .I(N__50485));
    LocalMux I__11498 (
            .O(N__50532),
            .I(N__50480));
    LocalMux I__11497 (
            .O(N__50521),
            .I(N__50480));
    LocalMux I__11496 (
            .O(N__50510),
            .I(N__50477));
    LocalMux I__11495 (
            .O(N__50507),
            .I(N__50474));
    LocalMux I__11494 (
            .O(N__50498),
            .I(N__50471));
    LocalMux I__11493 (
            .O(N__50495),
            .I(N__50466));
    LocalMux I__11492 (
            .O(N__50492),
            .I(N__50466));
    InMux I__11491 (
            .O(N__50491),
            .I(N__50461));
    InMux I__11490 (
            .O(N__50490),
            .I(N__50461));
    LocalMux I__11489 (
            .O(N__50485),
            .I(N__50456));
    Span4Mux_h I__11488 (
            .O(N__50480),
            .I(N__50452));
    Span12Mux_v I__11487 (
            .O(N__50477),
            .I(N__50449));
    Span4Mux_h I__11486 (
            .O(N__50474),
            .I(N__50440));
    Span4Mux_v I__11485 (
            .O(N__50471),
            .I(N__50440));
    Span4Mux_v I__11484 (
            .O(N__50466),
            .I(N__50440));
    LocalMux I__11483 (
            .O(N__50461),
            .I(N__50440));
    InMux I__11482 (
            .O(N__50460),
            .I(N__50435));
    InMux I__11481 (
            .O(N__50459),
            .I(N__50435));
    Span4Mux_h I__11480 (
            .O(N__50456),
            .I(N__50432));
    InMux I__11479 (
            .O(N__50455),
            .I(N__50429));
    Odrv4 I__11478 (
            .O(N__50452),
            .I(dds_state_2));
    Odrv12 I__11477 (
            .O(N__50449),
            .I(dds_state_2));
    Odrv4 I__11476 (
            .O(N__50440),
            .I(dds_state_2));
    LocalMux I__11475 (
            .O(N__50435),
            .I(dds_state_2));
    Odrv4 I__11474 (
            .O(N__50432),
            .I(dds_state_2));
    LocalMux I__11473 (
            .O(N__50429),
            .I(dds_state_2));
    InMux I__11472 (
            .O(N__50416),
            .I(N__50390));
    InMux I__11471 (
            .O(N__50415),
            .I(N__50390));
    InMux I__11470 (
            .O(N__50414),
            .I(N__50390));
    InMux I__11469 (
            .O(N__50413),
            .I(N__50390));
    InMux I__11468 (
            .O(N__50412),
            .I(N__50390));
    InMux I__11467 (
            .O(N__50411),
            .I(N__50390));
    InMux I__11466 (
            .O(N__50410),
            .I(N__50379));
    InMux I__11465 (
            .O(N__50409),
            .I(N__50379));
    InMux I__11464 (
            .O(N__50408),
            .I(N__50379));
    InMux I__11463 (
            .O(N__50407),
            .I(N__50379));
    InMux I__11462 (
            .O(N__50406),
            .I(N__50379));
    SRMux I__11461 (
            .O(N__50405),
            .I(N__50376));
    CEMux I__11460 (
            .O(N__50404),
            .I(N__50369));
    InMux I__11459 (
            .O(N__50403),
            .I(N__50365));
    LocalMux I__11458 (
            .O(N__50390),
            .I(N__50360));
    LocalMux I__11457 (
            .O(N__50379),
            .I(N__50357));
    LocalMux I__11456 (
            .O(N__50376),
            .I(N__50354));
    InMux I__11455 (
            .O(N__50375),
            .I(N__50345));
    InMux I__11454 (
            .O(N__50374),
            .I(N__50345));
    InMux I__11453 (
            .O(N__50373),
            .I(N__50345));
    InMux I__11452 (
            .O(N__50372),
            .I(N__50345));
    LocalMux I__11451 (
            .O(N__50369),
            .I(N__50342));
    InMux I__11450 (
            .O(N__50368),
            .I(N__50339));
    LocalMux I__11449 (
            .O(N__50365),
            .I(N__50336));
    InMux I__11448 (
            .O(N__50364),
            .I(N__50331));
    InMux I__11447 (
            .O(N__50363),
            .I(N__50331));
    Span4Mux_v I__11446 (
            .O(N__50360),
            .I(N__50326));
    Span4Mux_h I__11445 (
            .O(N__50357),
            .I(N__50319));
    Span4Mux_h I__11444 (
            .O(N__50354),
            .I(N__50319));
    LocalMux I__11443 (
            .O(N__50345),
            .I(N__50319));
    Span4Mux_v I__11442 (
            .O(N__50342),
            .I(N__50311));
    LocalMux I__11441 (
            .O(N__50339),
            .I(N__50304));
    Span4Mux_h I__11440 (
            .O(N__50336),
            .I(N__50304));
    LocalMux I__11439 (
            .O(N__50331),
            .I(N__50304));
    InMux I__11438 (
            .O(N__50330),
            .I(N__50301));
    InMux I__11437 (
            .O(N__50329),
            .I(N__50298));
    Span4Mux_h I__11436 (
            .O(N__50326),
            .I(N__50293));
    Span4Mux_h I__11435 (
            .O(N__50319),
            .I(N__50293));
    InMux I__11434 (
            .O(N__50318),
            .I(N__50288));
    InMux I__11433 (
            .O(N__50317),
            .I(N__50288));
    InMux I__11432 (
            .O(N__50316),
            .I(N__50281));
    InMux I__11431 (
            .O(N__50315),
            .I(N__50281));
    InMux I__11430 (
            .O(N__50314),
            .I(N__50281));
    Span4Mux_h I__11429 (
            .O(N__50311),
            .I(N__50276));
    Span4Mux_h I__11428 (
            .O(N__50304),
            .I(N__50276));
    LocalMux I__11427 (
            .O(N__50301),
            .I(dds_state_1));
    LocalMux I__11426 (
            .O(N__50298),
            .I(dds_state_1));
    Odrv4 I__11425 (
            .O(N__50293),
            .I(dds_state_1));
    LocalMux I__11424 (
            .O(N__50288),
            .I(dds_state_1));
    LocalMux I__11423 (
            .O(N__50281),
            .I(dds_state_1));
    Odrv4 I__11422 (
            .O(N__50276),
            .I(dds_state_1));
    IoInMux I__11421 (
            .O(N__50263),
            .I(N__50260));
    LocalMux I__11420 (
            .O(N__50260),
            .I(N__50257));
    IoSpan4Mux I__11419 (
            .O(N__50257),
            .I(N__50254));
    Sp12to4 I__11418 (
            .O(N__50254),
            .I(N__50251));
    Span12Mux_s6_v I__11417 (
            .O(N__50251),
            .I(N__50248));
    Odrv12 I__11416 (
            .O(N__50248),
            .I(DDS_CS));
    CEMux I__11415 (
            .O(N__50245),
            .I(N__50242));
    LocalMux I__11414 (
            .O(N__50242),
            .I(N__50239));
    Span4Mux_v I__11413 (
            .O(N__50239),
            .I(N__50236));
    Odrv4 I__11412 (
            .O(N__50236),
            .I(\SIG_DDS.n9_adj_1490 ));
    InMux I__11411 (
            .O(N__50233),
            .I(N__50230));
    LocalMux I__11410 (
            .O(N__50230),
            .I(N__50227));
    Span4Mux_v I__11409 (
            .O(N__50227),
            .I(N__50224));
    Odrv4 I__11408 (
            .O(N__50224),
            .I(buf_data_iac_23));
    CascadeMux I__11407 (
            .O(N__50221),
            .I(N__50218));
    InMux I__11406 (
            .O(N__50218),
            .I(N__50215));
    LocalMux I__11405 (
            .O(N__50215),
            .I(N__50212));
    Span4Mux_h I__11404 (
            .O(N__50212),
            .I(N__50209));
    Sp12to4 I__11403 (
            .O(N__50209),
            .I(N__50206));
    Span12Mux_v I__11402 (
            .O(N__50206),
            .I(N__50203));
    Odrv12 I__11401 (
            .O(N__50203),
            .I(n22595));
    InMux I__11400 (
            .O(N__50200),
            .I(N__50195));
    InMux I__11399 (
            .O(N__50199),
            .I(N__50192));
    InMux I__11398 (
            .O(N__50198),
            .I(N__50189));
    LocalMux I__11397 (
            .O(N__50195),
            .I(N__50185));
    LocalMux I__11396 (
            .O(N__50192),
            .I(N__50180));
    LocalMux I__11395 (
            .O(N__50189),
            .I(N__50180));
    InMux I__11394 (
            .O(N__50188),
            .I(N__50177));
    Span4Mux_v I__11393 (
            .O(N__50185),
            .I(N__50174));
    Span4Mux_v I__11392 (
            .O(N__50180),
            .I(N__50169));
    LocalMux I__11391 (
            .O(N__50177),
            .I(N__50169));
    Span4Mux_h I__11390 (
            .O(N__50174),
            .I(N__50165));
    Span4Mux_v I__11389 (
            .O(N__50169),
            .I(N__50162));
    InMux I__11388 (
            .O(N__50168),
            .I(N__50159));
    Span4Mux_v I__11387 (
            .O(N__50165),
            .I(N__50156));
    Span4Mux_v I__11386 (
            .O(N__50162),
            .I(N__50153));
    LocalMux I__11385 (
            .O(N__50159),
            .I(N__50150));
    Sp12to4 I__11384 (
            .O(N__50156),
            .I(N__50143));
    Sp12to4 I__11383 (
            .O(N__50153),
            .I(N__50143));
    Span12Mux_v I__11382 (
            .O(N__50150),
            .I(N__50143));
    Odrv12 I__11381 (
            .O(N__50143),
            .I(ICE_SPI_MOSI));
    SRMux I__11380 (
            .O(N__50140),
            .I(N__50137));
    LocalMux I__11379 (
            .O(N__50137),
            .I(N__50134));
    Odrv4 I__11378 (
            .O(N__50134),
            .I(\comm_spi.imosi_N_840 ));
    InMux I__11377 (
            .O(N__50131),
            .I(n20630));
    InMux I__11376 (
            .O(N__50128),
            .I(N__50124));
    CascadeMux I__11375 (
            .O(N__50127),
            .I(N__50121));
    LocalMux I__11374 (
            .O(N__50124),
            .I(N__50118));
    InMux I__11373 (
            .O(N__50121),
            .I(N__50114));
    Span4Mux_v I__11372 (
            .O(N__50118),
            .I(N__50111));
    InMux I__11371 (
            .O(N__50117),
            .I(N__50108));
    LocalMux I__11370 (
            .O(N__50114),
            .I(N__50105));
    Span4Mux_h I__11369 (
            .O(N__50111),
            .I(N__50102));
    LocalMux I__11368 (
            .O(N__50108),
            .I(N__50097));
    Span4Mux_h I__11367 (
            .O(N__50105),
            .I(N__50097));
    Odrv4 I__11366 (
            .O(N__50102),
            .I(data_cntvec_10));
    Odrv4 I__11365 (
            .O(N__50097),
            .I(data_cntvec_10));
    InMux I__11364 (
            .O(N__50092),
            .I(n20631));
    InMux I__11363 (
            .O(N__50089),
            .I(n20632));
    InMux I__11362 (
            .O(N__50086),
            .I(N__50083));
    LocalMux I__11361 (
            .O(N__50083),
            .I(N__50079));
    InMux I__11360 (
            .O(N__50082),
            .I(N__50076));
    Span4Mux_h I__11359 (
            .O(N__50079),
            .I(N__50073));
    LocalMux I__11358 (
            .O(N__50076),
            .I(data_cntvec_12));
    Odrv4 I__11357 (
            .O(N__50073),
            .I(data_cntvec_12));
    InMux I__11356 (
            .O(N__50068),
            .I(n20633));
    InMux I__11355 (
            .O(N__50065),
            .I(N__50062));
    LocalMux I__11354 (
            .O(N__50062),
            .I(N__50059));
    Span4Mux_h I__11353 (
            .O(N__50059),
            .I(N__50055));
    InMux I__11352 (
            .O(N__50058),
            .I(N__50052));
    Span4Mux_h I__11351 (
            .O(N__50055),
            .I(N__50049));
    LocalMux I__11350 (
            .O(N__50052),
            .I(data_cntvec_13));
    Odrv4 I__11349 (
            .O(N__50049),
            .I(data_cntvec_13));
    InMux I__11348 (
            .O(N__50044),
            .I(n20634));
    InMux I__11347 (
            .O(N__50041),
            .I(n20635));
    InMux I__11346 (
            .O(N__50038),
            .I(n20636));
    InMux I__11345 (
            .O(N__50035),
            .I(N__50031));
    InMux I__11344 (
            .O(N__50034),
            .I(N__50028));
    LocalMux I__11343 (
            .O(N__50031),
            .I(N__50025));
    LocalMux I__11342 (
            .O(N__50028),
            .I(data_cntvec_15));
    Odrv4 I__11341 (
            .O(N__50025),
            .I(data_cntvec_15));
    InMux I__11340 (
            .O(N__50020),
            .I(N__50014));
    CEMux I__11339 (
            .O(N__50019),
            .I(N__50010));
    CEMux I__11338 (
            .O(N__50018),
            .I(N__50007));
    CEMux I__11337 (
            .O(N__50017),
            .I(N__50004));
    LocalMux I__11336 (
            .O(N__50014),
            .I(N__50001));
    CEMux I__11335 (
            .O(N__50013),
            .I(N__49998));
    LocalMux I__11334 (
            .O(N__50010),
            .I(N__49995));
    LocalMux I__11333 (
            .O(N__50007),
            .I(N__49992));
    LocalMux I__11332 (
            .O(N__50004),
            .I(N__49989));
    Span4Mux_v I__11331 (
            .O(N__50001),
            .I(N__49986));
    LocalMux I__11330 (
            .O(N__49998),
            .I(N__49983));
    Span4Mux_h I__11329 (
            .O(N__49995),
            .I(N__49978));
    Span4Mux_h I__11328 (
            .O(N__49992),
            .I(N__49978));
    Span4Mux_v I__11327 (
            .O(N__49989),
            .I(N__49973));
    Span4Mux_v I__11326 (
            .O(N__49986),
            .I(N__49973));
    Span4Mux_h I__11325 (
            .O(N__49983),
            .I(N__49970));
    Sp12to4 I__11324 (
            .O(N__49978),
            .I(N__49967));
    Span4Mux_h I__11323 (
            .O(N__49973),
            .I(N__49964));
    Odrv4 I__11322 (
            .O(N__49970),
            .I(n12394));
    Odrv12 I__11321 (
            .O(N__49967),
            .I(n12394));
    Odrv4 I__11320 (
            .O(N__49964),
            .I(n12394));
    SRMux I__11319 (
            .O(N__49957),
            .I(N__49953));
    SRMux I__11318 (
            .O(N__49956),
            .I(N__49950));
    LocalMux I__11317 (
            .O(N__49953),
            .I(N__49947));
    LocalMux I__11316 (
            .O(N__49950),
            .I(N__49944));
    Span4Mux_v I__11315 (
            .O(N__49947),
            .I(N__49939));
    Span4Mux_v I__11314 (
            .O(N__49944),
            .I(N__49936));
    SRMux I__11313 (
            .O(N__49943),
            .I(N__49933));
    SRMux I__11312 (
            .O(N__49942),
            .I(N__49930));
    Span4Mux_h I__11311 (
            .O(N__49939),
            .I(N__49925));
    Span4Mux_h I__11310 (
            .O(N__49936),
            .I(N__49925));
    LocalMux I__11309 (
            .O(N__49933),
            .I(N__49922));
    LocalMux I__11308 (
            .O(N__49930),
            .I(N__49919));
    Span4Mux_h I__11307 (
            .O(N__49925),
            .I(N__49912));
    Span4Mux_v I__11306 (
            .O(N__49922),
            .I(N__49912));
    Span4Mux_v I__11305 (
            .O(N__49919),
            .I(N__49912));
    Odrv4 I__11304 (
            .O(N__49912),
            .I(n15431));
    InMux I__11303 (
            .O(N__49909),
            .I(N__49906));
    LocalMux I__11302 (
            .O(N__49906),
            .I(N__49903));
    Span4Mux_h I__11301 (
            .O(N__49903),
            .I(N__49900));
    Odrv4 I__11300 (
            .O(N__49900),
            .I(n23480));
    IoInMux I__11299 (
            .O(N__49897),
            .I(N__49894));
    LocalMux I__11298 (
            .O(N__49894),
            .I(N__49891));
    IoSpan4Mux I__11297 (
            .O(N__49891),
            .I(N__49888));
    IoSpan4Mux I__11296 (
            .O(N__49888),
            .I(N__49885));
    Span4Mux_s1_v I__11295 (
            .O(N__49885),
            .I(N__49881));
    CascadeMux I__11294 (
            .O(N__49884),
            .I(N__49878));
    Span4Mux_v I__11293 (
            .O(N__49881),
            .I(N__49875));
    InMux I__11292 (
            .O(N__49878),
            .I(N__49872));
    Span4Mux_v I__11291 (
            .O(N__49875),
            .I(N__49867));
    LocalMux I__11290 (
            .O(N__49872),
            .I(N__49867));
    Span4Mux_h I__11289 (
            .O(N__49867),
            .I(N__49863));
    InMux I__11288 (
            .O(N__49866),
            .I(N__49860));
    Span4Mux_v I__11287 (
            .O(N__49863),
            .I(N__49857));
    LocalMux I__11286 (
            .O(N__49860),
            .I(DDS_RNG_0));
    Odrv4 I__11285 (
            .O(N__49857),
            .I(DDS_RNG_0));
    InMux I__11284 (
            .O(N__49852),
            .I(N__49849));
    LocalMux I__11283 (
            .O(N__49849),
            .I(N__49845));
    InMux I__11282 (
            .O(N__49848),
            .I(N__49841));
    Span12Mux_h I__11281 (
            .O(N__49845),
            .I(N__49838));
    InMux I__11280 (
            .O(N__49844),
            .I(N__49835));
    LocalMux I__11279 (
            .O(N__49841),
            .I(acadc_skipCount_9));
    Odrv12 I__11278 (
            .O(N__49838),
            .I(acadc_skipCount_9));
    LocalMux I__11277 (
            .O(N__49835),
            .I(acadc_skipCount_9));
    CascadeMux I__11276 (
            .O(N__49828),
            .I(n22183_cascade_));
    InMux I__11275 (
            .O(N__49825),
            .I(n20622));
    InMux I__11274 (
            .O(N__49822),
            .I(n20623));
    InMux I__11273 (
            .O(N__49819),
            .I(N__49816));
    LocalMux I__11272 (
            .O(N__49816),
            .I(N__49812));
    InMux I__11271 (
            .O(N__49815),
            .I(N__49808));
    Span4Mux_h I__11270 (
            .O(N__49812),
            .I(N__49805));
    InMux I__11269 (
            .O(N__49811),
            .I(N__49802));
    LocalMux I__11268 (
            .O(N__49808),
            .I(data_cntvec_3));
    Odrv4 I__11267 (
            .O(N__49805),
            .I(data_cntvec_3));
    LocalMux I__11266 (
            .O(N__49802),
            .I(data_cntvec_3));
    InMux I__11265 (
            .O(N__49795),
            .I(n20624));
    InMux I__11264 (
            .O(N__49792),
            .I(n20625));
    InMux I__11263 (
            .O(N__49789),
            .I(n20626));
    InMux I__11262 (
            .O(N__49786),
            .I(N__49783));
    LocalMux I__11261 (
            .O(N__49783),
            .I(N__49779));
    InMux I__11260 (
            .O(N__49782),
            .I(N__49775));
    Span4Mux_h I__11259 (
            .O(N__49779),
            .I(N__49772));
    InMux I__11258 (
            .O(N__49778),
            .I(N__49769));
    LocalMux I__11257 (
            .O(N__49775),
            .I(data_cntvec_6));
    Odrv4 I__11256 (
            .O(N__49772),
            .I(data_cntvec_6));
    LocalMux I__11255 (
            .O(N__49769),
            .I(data_cntvec_6));
    InMux I__11254 (
            .O(N__49762),
            .I(n20627));
    InMux I__11253 (
            .O(N__49759),
            .I(n20628));
    InMux I__11252 (
            .O(N__49756),
            .I(N__49753));
    LocalMux I__11251 (
            .O(N__49753),
            .I(N__49750));
    Span4Mux_h I__11250 (
            .O(N__49750),
            .I(N__49747));
    Span4Mux_h I__11249 (
            .O(N__49747),
            .I(N__49743));
    InMux I__11248 (
            .O(N__49746),
            .I(N__49739));
    Span4Mux_h I__11247 (
            .O(N__49743),
            .I(N__49736));
    InMux I__11246 (
            .O(N__49742),
            .I(N__49733));
    LocalMux I__11245 (
            .O(N__49739),
            .I(data_cntvec_8));
    Odrv4 I__11244 (
            .O(N__49736),
            .I(data_cntvec_8));
    LocalMux I__11243 (
            .O(N__49733),
            .I(data_cntvec_8));
    InMux I__11242 (
            .O(N__49726),
            .I(bfn_17_16_0_));
    InMux I__11241 (
            .O(N__49723),
            .I(N__49720));
    LocalMux I__11240 (
            .O(N__49720),
            .I(N__49716));
    InMux I__11239 (
            .O(N__49719),
            .I(N__49713));
    Span4Mux_h I__11238 (
            .O(N__49716),
            .I(N__49710));
    LocalMux I__11237 (
            .O(N__49713),
            .I(data_idxvec_12));
    Odrv4 I__11236 (
            .O(N__49710),
            .I(data_idxvec_12));
    InMux I__11235 (
            .O(N__49705),
            .I(N__49702));
    LocalMux I__11234 (
            .O(N__49702),
            .I(N__49699));
    Span4Mux_v I__11233 (
            .O(N__49699),
            .I(N__49696));
    Sp12to4 I__11232 (
            .O(N__49696),
            .I(N__49693));
    Odrv12 I__11231 (
            .O(N__49693),
            .I(n22499));
    InMux I__11230 (
            .O(N__49690),
            .I(N__49687));
    LocalMux I__11229 (
            .O(N__49687),
            .I(N__49684));
    Span4Mux_h I__11228 (
            .O(N__49684),
            .I(N__49679));
    InMux I__11227 (
            .O(N__49683),
            .I(N__49674));
    InMux I__11226 (
            .O(N__49682),
            .I(N__49674));
    Odrv4 I__11225 (
            .O(N__49679),
            .I(acadc_skipCount_6));
    LocalMux I__11224 (
            .O(N__49674),
            .I(acadc_skipCount_6));
    CascadeMux I__11223 (
            .O(N__49669),
            .I(N__49666));
    InMux I__11222 (
            .O(N__49666),
            .I(N__49663));
    LocalMux I__11221 (
            .O(N__49663),
            .I(N__49660));
    Span4Mux_h I__11220 (
            .O(N__49660),
            .I(N__49657));
    Sp12to4 I__11219 (
            .O(N__49657),
            .I(N__49652));
    InMux I__11218 (
            .O(N__49656),
            .I(N__49647));
    InMux I__11217 (
            .O(N__49655),
            .I(N__49647));
    Odrv12 I__11216 (
            .O(N__49652),
            .I(req_data_cnt_6));
    LocalMux I__11215 (
            .O(N__49647),
            .I(req_data_cnt_6));
    CascadeMux I__11214 (
            .O(N__49642),
            .I(n23519_cascade_));
    InMux I__11213 (
            .O(N__49639),
            .I(N__49636));
    LocalMux I__11212 (
            .O(N__49636),
            .I(N__49633));
    Span4Mux_h I__11211 (
            .O(N__49633),
            .I(N__49630));
    Odrv4 I__11210 (
            .O(N__49630),
            .I(n23291));
    InMux I__11209 (
            .O(N__49627),
            .I(N__49624));
    LocalMux I__11208 (
            .O(N__49624),
            .I(N__49621));
    Odrv12 I__11207 (
            .O(N__49621),
            .I(n111_adj_1726));
    CascadeMux I__11206 (
            .O(N__49618),
            .I(n30_adj_1724_cascade_));
    InMux I__11205 (
            .O(N__49615),
            .I(N__49612));
    LocalMux I__11204 (
            .O(N__49612),
            .I(comm_buf_1_7_N_559_6));
    InMux I__11203 (
            .O(N__49609),
            .I(N__49606));
    LocalMux I__11202 (
            .O(N__49606),
            .I(N__49602));
    InMux I__11201 (
            .O(N__49605),
            .I(N__49599));
    Span4Mux_v I__11200 (
            .O(N__49602),
            .I(N__49596));
    LocalMux I__11199 (
            .O(N__49599),
            .I(data_idxvec_6));
    Odrv4 I__11198 (
            .O(N__49596),
            .I(data_idxvec_6));
    CascadeMux I__11197 (
            .O(N__49591),
            .I(n26_adj_1723_cascade_));
    InMux I__11196 (
            .O(N__49588),
            .I(N__49585));
    LocalMux I__11195 (
            .O(N__49585),
            .I(n23516));
    InMux I__11194 (
            .O(N__49582),
            .I(N__49579));
    LocalMux I__11193 (
            .O(N__49579),
            .I(n23303));
    InMux I__11192 (
            .O(N__49576),
            .I(N__49573));
    LocalMux I__11191 (
            .O(N__49573),
            .I(n23555));
    InMux I__11190 (
            .O(N__49570),
            .I(N__49564));
    InMux I__11189 (
            .O(N__49569),
            .I(N__49552));
    InMux I__11188 (
            .O(N__49568),
            .I(N__49552));
    InMux I__11187 (
            .O(N__49567),
            .I(N__49552));
    LocalMux I__11186 (
            .O(N__49564),
            .I(N__49549));
    InMux I__11185 (
            .O(N__49563),
            .I(N__49546));
    InMux I__11184 (
            .O(N__49562),
            .I(N__49543));
    InMux I__11183 (
            .O(N__49561),
            .I(N__49538));
    InMux I__11182 (
            .O(N__49560),
            .I(N__49538));
    InMux I__11181 (
            .O(N__49559),
            .I(N__49534));
    LocalMux I__11180 (
            .O(N__49552),
            .I(N__49531));
    Span4Mux_v I__11179 (
            .O(N__49549),
            .I(N__49522));
    LocalMux I__11178 (
            .O(N__49546),
            .I(N__49522));
    LocalMux I__11177 (
            .O(N__49543),
            .I(N__49522));
    LocalMux I__11176 (
            .O(N__49538),
            .I(N__49522));
    InMux I__11175 (
            .O(N__49537),
            .I(N__49519));
    LocalMux I__11174 (
            .O(N__49534),
            .I(N__49515));
    Span4Mux_v I__11173 (
            .O(N__49531),
            .I(N__49510));
    Span4Mux_v I__11172 (
            .O(N__49522),
            .I(N__49510));
    LocalMux I__11171 (
            .O(N__49519),
            .I(N__49507));
    InMux I__11170 (
            .O(N__49518),
            .I(N__49504));
    Span4Mux_h I__11169 (
            .O(N__49515),
            .I(N__49499));
    Span4Mux_h I__11168 (
            .O(N__49510),
            .I(N__49494));
    Span4Mux_v I__11167 (
            .O(N__49507),
            .I(N__49494));
    LocalMux I__11166 (
            .O(N__49504),
            .I(N__49491));
    InMux I__11165 (
            .O(N__49503),
            .I(N__49488));
    InMux I__11164 (
            .O(N__49502),
            .I(N__49485));
    Span4Mux_h I__11163 (
            .O(N__49499),
            .I(N__49482));
    Span4Mux_h I__11162 (
            .O(N__49494),
            .I(N__49479));
    Span12Mux_v I__11161 (
            .O(N__49491),
            .I(N__49474));
    LocalMux I__11160 (
            .O(N__49488),
            .I(N__49474));
    LocalMux I__11159 (
            .O(N__49485),
            .I(N__49471));
    Odrv4 I__11158 (
            .O(N__49482),
            .I(n18363));
    Odrv4 I__11157 (
            .O(N__49479),
            .I(n18363));
    Odrv12 I__11156 (
            .O(N__49474),
            .I(n18363));
    Odrv12 I__11155 (
            .O(N__49471),
            .I(n18363));
    InMux I__11154 (
            .O(N__49462),
            .I(N__49459));
    LocalMux I__11153 (
            .O(N__49459),
            .I(N__49454));
    InMux I__11152 (
            .O(N__49458),
            .I(N__49451));
    InMux I__11151 (
            .O(N__49457),
            .I(N__49448));
    Span12Mux_s10_h I__11150 (
            .O(N__49454),
            .I(N__49443));
    LocalMux I__11149 (
            .O(N__49451),
            .I(N__49443));
    LocalMux I__11148 (
            .O(N__49448),
            .I(buf_dds1_4));
    Odrv12 I__11147 (
            .O(N__49443),
            .I(buf_dds1_4));
    CascadeMux I__11146 (
            .O(N__49438),
            .I(N__49432));
    CascadeMux I__11145 (
            .O(N__49437),
            .I(N__49429));
    InMux I__11144 (
            .O(N__49436),
            .I(N__49424));
    InMux I__11143 (
            .O(N__49435),
            .I(N__49424));
    InMux I__11142 (
            .O(N__49432),
            .I(N__49421));
    InMux I__11141 (
            .O(N__49429),
            .I(N__49418));
    LocalMux I__11140 (
            .O(N__49424),
            .I(N__49413));
    LocalMux I__11139 (
            .O(N__49421),
            .I(N__49413));
    LocalMux I__11138 (
            .O(N__49418),
            .I(N__49409));
    Span12Mux_h I__11137 (
            .O(N__49413),
            .I(N__49406));
    InMux I__11136 (
            .O(N__49412),
            .I(N__49403));
    Odrv4 I__11135 (
            .O(N__49409),
            .I(iac_raw_buf_N_823));
    Odrv12 I__11134 (
            .O(N__49406),
            .I(iac_raw_buf_N_823));
    LocalMux I__11133 (
            .O(N__49403),
            .I(iac_raw_buf_N_823));
    InMux I__11132 (
            .O(N__49396),
            .I(N__49393));
    LocalMux I__11131 (
            .O(N__49393),
            .I(N__49389));
    InMux I__11130 (
            .O(N__49392),
            .I(N__49385));
    Span4Mux_h I__11129 (
            .O(N__49389),
            .I(N__49382));
    InMux I__11128 (
            .O(N__49388),
            .I(N__49379));
    LocalMux I__11127 (
            .O(N__49385),
            .I(data_cntvec_0));
    Odrv4 I__11126 (
            .O(N__49382),
            .I(data_cntvec_0));
    LocalMux I__11125 (
            .O(N__49379),
            .I(data_cntvec_0));
    InMux I__11124 (
            .O(N__49372),
            .I(N__49369));
    LocalMux I__11123 (
            .O(N__49369),
            .I(n22351));
    CascadeMux I__11122 (
            .O(N__49366),
            .I(n4_adj_1709_cascade_));
    CascadeMux I__11121 (
            .O(N__49363),
            .I(N__49359));
    CascadeMux I__11120 (
            .O(N__49362),
            .I(N__49356));
    InMux I__11119 (
            .O(N__49359),
            .I(N__49351));
    InMux I__11118 (
            .O(N__49356),
            .I(N__49351));
    LocalMux I__11117 (
            .O(N__49351),
            .I(n35));
    InMux I__11116 (
            .O(N__49348),
            .I(N__49345));
    LocalMux I__11115 (
            .O(N__49345),
            .I(n12_adj_1802));
    InMux I__11114 (
            .O(N__49342),
            .I(N__49339));
    LocalMux I__11113 (
            .O(N__49339),
            .I(N__49336));
    Span4Mux_h I__11112 (
            .O(N__49336),
            .I(N__49333));
    Odrv4 I__11111 (
            .O(N__49333),
            .I(comm_buf_1_7_N_559_3));
    InMux I__11110 (
            .O(N__49330),
            .I(N__49327));
    LocalMux I__11109 (
            .O(N__49327),
            .I(N__49323));
    InMux I__11108 (
            .O(N__49326),
            .I(N__49319));
    Span4Mux_h I__11107 (
            .O(N__49323),
            .I(N__49315));
    InMux I__11106 (
            .O(N__49322),
            .I(N__49312));
    LocalMux I__11105 (
            .O(N__49319),
            .I(N__49308));
    InMux I__11104 (
            .O(N__49318),
            .I(N__49305));
    Span4Mux_h I__11103 (
            .O(N__49315),
            .I(N__49300));
    LocalMux I__11102 (
            .O(N__49312),
            .I(N__49300));
    CascadeMux I__11101 (
            .O(N__49311),
            .I(N__49297));
    Span4Mux_h I__11100 (
            .O(N__49308),
            .I(N__49294));
    LocalMux I__11099 (
            .O(N__49305),
            .I(N__49289));
    Span4Mux_v I__11098 (
            .O(N__49300),
            .I(N__49286));
    InMux I__11097 (
            .O(N__49297),
            .I(N__49283));
    Span4Mux_v I__11096 (
            .O(N__49294),
            .I(N__49280));
    InMux I__11095 (
            .O(N__49293),
            .I(N__49277));
    CascadeMux I__11094 (
            .O(N__49292),
            .I(N__49274));
    Span4Mux_h I__11093 (
            .O(N__49289),
            .I(N__49268));
    Span4Mux_h I__11092 (
            .O(N__49286),
            .I(N__49268));
    LocalMux I__11091 (
            .O(N__49283),
            .I(N__49261));
    Sp12to4 I__11090 (
            .O(N__49280),
            .I(N__49261));
    LocalMux I__11089 (
            .O(N__49277),
            .I(N__49261));
    InMux I__11088 (
            .O(N__49274),
            .I(N__49258));
    InMux I__11087 (
            .O(N__49273),
            .I(N__49255));
    Sp12to4 I__11086 (
            .O(N__49268),
            .I(N__49250));
    Span12Mux_v I__11085 (
            .O(N__49261),
            .I(N__49250));
    LocalMux I__11084 (
            .O(N__49258),
            .I(comm_buf_1_3));
    LocalMux I__11083 (
            .O(N__49255),
            .I(comm_buf_1_3));
    Odrv12 I__11082 (
            .O(N__49250),
            .I(comm_buf_1_3));
    CascadeMux I__11081 (
            .O(N__49243),
            .I(N__49240));
    InMux I__11080 (
            .O(N__49240),
            .I(N__49236));
    InMux I__11079 (
            .O(N__49239),
            .I(N__49233));
    LocalMux I__11078 (
            .O(N__49236),
            .I(N__49225));
    LocalMux I__11077 (
            .O(N__49233),
            .I(N__49225));
    InMux I__11076 (
            .O(N__49232),
            .I(N__49222));
    InMux I__11075 (
            .O(N__49231),
            .I(N__49218));
    InMux I__11074 (
            .O(N__49230),
            .I(N__49215));
    Span4Mux_v I__11073 (
            .O(N__49225),
            .I(N__49211));
    LocalMux I__11072 (
            .O(N__49222),
            .I(N__49208));
    InMux I__11071 (
            .O(N__49221),
            .I(N__49205));
    LocalMux I__11070 (
            .O(N__49218),
            .I(N__49202));
    LocalMux I__11069 (
            .O(N__49215),
            .I(N__49199));
    InMux I__11068 (
            .O(N__49214),
            .I(N__49196));
    Span4Mux_v I__11067 (
            .O(N__49211),
            .I(N__49193));
    Span4Mux_v I__11066 (
            .O(N__49208),
            .I(N__49188));
    LocalMux I__11065 (
            .O(N__49205),
            .I(N__49188));
    Span4Mux_h I__11064 (
            .O(N__49202),
            .I(N__49185));
    Span4Mux_v I__11063 (
            .O(N__49199),
            .I(N__49182));
    LocalMux I__11062 (
            .O(N__49196),
            .I(N__49179));
    Sp12to4 I__11061 (
            .O(N__49193),
            .I(N__49176));
    Span4Mux_h I__11060 (
            .O(N__49188),
            .I(N__49173));
    Span4Mux_h I__11059 (
            .O(N__49185),
            .I(N__49170));
    Sp12to4 I__11058 (
            .O(N__49182),
            .I(N__49165));
    Span12Mux_h I__11057 (
            .O(N__49179),
            .I(N__49165));
    Span12Mux_h I__11056 (
            .O(N__49176),
            .I(N__49162));
    Span4Mux_v I__11055 (
            .O(N__49173),
            .I(N__49159));
    Odrv4 I__11054 (
            .O(N__49170),
            .I(comm_buf_1_6));
    Odrv12 I__11053 (
            .O(N__49165),
            .I(comm_buf_1_6));
    Odrv12 I__11052 (
            .O(N__49162),
            .I(comm_buf_1_6));
    Odrv4 I__11051 (
            .O(N__49159),
            .I(comm_buf_1_6));
    CascadeMux I__11050 (
            .O(N__49150),
            .I(N__49147));
    InMux I__11049 (
            .O(N__49147),
            .I(N__49143));
    InMux I__11048 (
            .O(N__49146),
            .I(N__49137));
    LocalMux I__11047 (
            .O(N__49143),
            .I(N__49134));
    CascadeMux I__11046 (
            .O(N__49142),
            .I(N__49130));
    CascadeMux I__11045 (
            .O(N__49141),
            .I(N__49126));
    CascadeMux I__11044 (
            .O(N__49140),
            .I(N__49123));
    LocalMux I__11043 (
            .O(N__49137),
            .I(N__49119));
    Span4Mux_v I__11042 (
            .O(N__49134),
            .I(N__49116));
    CascadeMux I__11041 (
            .O(N__49133),
            .I(N__49113));
    InMux I__11040 (
            .O(N__49130),
            .I(N__49110));
    InMux I__11039 (
            .O(N__49129),
            .I(N__49107));
    InMux I__11038 (
            .O(N__49126),
            .I(N__49103));
    InMux I__11037 (
            .O(N__49123),
            .I(N__49100));
    InMux I__11036 (
            .O(N__49122),
            .I(N__49097));
    Span4Mux_v I__11035 (
            .O(N__49119),
            .I(N__49094));
    Span4Mux_v I__11034 (
            .O(N__49116),
            .I(N__49091));
    InMux I__11033 (
            .O(N__49113),
            .I(N__49088));
    LocalMux I__11032 (
            .O(N__49110),
            .I(N__49082));
    LocalMux I__11031 (
            .O(N__49107),
            .I(N__49082));
    InMux I__11030 (
            .O(N__49106),
            .I(N__49079));
    LocalMux I__11029 (
            .O(N__49103),
            .I(N__49076));
    LocalMux I__11028 (
            .O(N__49100),
            .I(N__49073));
    LocalMux I__11027 (
            .O(N__49097),
            .I(N__49066));
    Span4Mux_v I__11026 (
            .O(N__49094),
            .I(N__49066));
    Span4Mux_h I__11025 (
            .O(N__49091),
            .I(N__49066));
    LocalMux I__11024 (
            .O(N__49088),
            .I(N__49063));
    InMux I__11023 (
            .O(N__49087),
            .I(N__49060));
    Span4Mux_v I__11022 (
            .O(N__49082),
            .I(N__49057));
    LocalMux I__11021 (
            .O(N__49079),
            .I(N__49052));
    Span12Mux_v I__11020 (
            .O(N__49076),
            .I(N__49052));
    Span4Mux_v I__11019 (
            .O(N__49073),
            .I(N__49047));
    Span4Mux_h I__11018 (
            .O(N__49066),
            .I(N__49047));
    Span12Mux_h I__11017 (
            .O(N__49063),
            .I(N__49042));
    LocalMux I__11016 (
            .O(N__49060),
            .I(N__49042));
    Span4Mux_h I__11015 (
            .O(N__49057),
            .I(N__49039));
    Odrv12 I__11014 (
            .O(N__49052),
            .I(comm_buf_1_0));
    Odrv4 I__11013 (
            .O(N__49047),
            .I(comm_buf_1_0));
    Odrv12 I__11012 (
            .O(N__49042),
            .I(comm_buf_1_0));
    Odrv4 I__11011 (
            .O(N__49039),
            .I(comm_buf_1_0));
    InMux I__11010 (
            .O(N__49030),
            .I(N__49027));
    LocalMux I__11009 (
            .O(N__49027),
            .I(N__49023));
    InMux I__11008 (
            .O(N__49026),
            .I(N__49020));
    Span4Mux_v I__11007 (
            .O(N__49023),
            .I(N__49017));
    LocalMux I__11006 (
            .O(N__49020),
            .I(data_idxvec_14));
    Odrv4 I__11005 (
            .O(N__49017),
            .I(data_idxvec_14));
    CascadeMux I__11004 (
            .O(N__49012),
            .I(N__49009));
    InMux I__11003 (
            .O(N__49009),
            .I(N__49006));
    LocalMux I__11002 (
            .O(N__49006),
            .I(N__49003));
    Span4Mux_h I__11001 (
            .O(N__49003),
            .I(N__49000));
    Odrv4 I__11000 (
            .O(N__49000),
            .I(n22296));
    CascadeMux I__10999 (
            .O(N__48997),
            .I(n46_cascade_));
    CascadeMux I__10998 (
            .O(N__48994),
            .I(N__48990));
    InMux I__10997 (
            .O(N__48993),
            .I(N__48987));
    InMux I__10996 (
            .O(N__48990),
            .I(N__48983));
    LocalMux I__10995 (
            .O(N__48987),
            .I(N__48980));
    InMux I__10994 (
            .O(N__48986),
            .I(N__48977));
    LocalMux I__10993 (
            .O(N__48983),
            .I(N__48974));
    Span4Mux_h I__10992 (
            .O(N__48980),
            .I(N__48971));
    LocalMux I__10991 (
            .O(N__48977),
            .I(comm_test_buf_24_0));
    Odrv12 I__10990 (
            .O(N__48974),
            .I(comm_test_buf_24_0));
    Odrv4 I__10989 (
            .O(N__48971),
            .I(comm_test_buf_24_0));
    InMux I__10988 (
            .O(N__48964),
            .I(N__48961));
    LocalMux I__10987 (
            .O(N__48961),
            .I(N__48958));
    Span4Mux_v I__10986 (
            .O(N__48958),
            .I(N__48954));
    InMux I__10985 (
            .O(N__48957),
            .I(N__48951));
    Span4Mux_h I__10984 (
            .O(N__48954),
            .I(N__48946));
    LocalMux I__10983 (
            .O(N__48951),
            .I(N__48946));
    Odrv4 I__10982 (
            .O(N__48946),
            .I(comm_test_buf_24_8));
    InMux I__10981 (
            .O(N__48943),
            .I(N__48938));
    InMux I__10980 (
            .O(N__48942),
            .I(N__48935));
    CascadeMux I__10979 (
            .O(N__48941),
            .I(N__48932));
    LocalMux I__10978 (
            .O(N__48938),
            .I(N__48929));
    LocalMux I__10977 (
            .O(N__48935),
            .I(N__48926));
    InMux I__10976 (
            .O(N__48932),
            .I(N__48923));
    Span4Mux_v I__10975 (
            .O(N__48929),
            .I(N__48920));
    Span4Mux_h I__10974 (
            .O(N__48926),
            .I(N__48917));
    LocalMux I__10973 (
            .O(N__48923),
            .I(N__48912));
    Span4Mux_h I__10972 (
            .O(N__48920),
            .I(N__48912));
    Span4Mux_v I__10971 (
            .O(N__48917),
            .I(N__48909));
    Span4Mux_h I__10970 (
            .O(N__48912),
            .I(N__48906));
    Odrv4 I__10969 (
            .O(N__48909),
            .I(n14_adj_1662));
    Odrv4 I__10968 (
            .O(N__48906),
            .I(n14_adj_1662));
    InMux I__10967 (
            .O(N__48901),
            .I(N__48897));
    InMux I__10966 (
            .O(N__48900),
            .I(N__48894));
    LocalMux I__10965 (
            .O(N__48897),
            .I(n4_adj_1749));
    LocalMux I__10964 (
            .O(N__48894),
            .I(n4_adj_1749));
    InMux I__10963 (
            .O(N__48889),
            .I(N__48886));
    LocalMux I__10962 (
            .O(N__48886),
            .I(N__48883));
    Odrv12 I__10961 (
            .O(N__48883),
            .I(n12_adj_1684));
    InMux I__10960 (
            .O(N__48880),
            .I(N__48876));
    InMux I__10959 (
            .O(N__48879),
            .I(N__48873));
    LocalMux I__10958 (
            .O(N__48876),
            .I(N__48867));
    LocalMux I__10957 (
            .O(N__48873),
            .I(N__48864));
    InMux I__10956 (
            .O(N__48872),
            .I(N__48861));
    InMux I__10955 (
            .O(N__48871),
            .I(N__48858));
    InMux I__10954 (
            .O(N__48870),
            .I(N__48854));
    Span4Mux_h I__10953 (
            .O(N__48867),
            .I(N__48849));
    Span4Mux_v I__10952 (
            .O(N__48864),
            .I(N__48849));
    LocalMux I__10951 (
            .O(N__48861),
            .I(N__48846));
    LocalMux I__10950 (
            .O(N__48858),
            .I(N__48843));
    InMux I__10949 (
            .O(N__48857),
            .I(N__48840));
    LocalMux I__10948 (
            .O(N__48854),
            .I(N__48833));
    Span4Mux_h I__10947 (
            .O(N__48849),
            .I(N__48833));
    Span4Mux_h I__10946 (
            .O(N__48846),
            .I(N__48833));
    Span4Mux_h I__10945 (
            .O(N__48843),
            .I(N__48830));
    LocalMux I__10944 (
            .O(N__48840),
            .I(N__48827));
    Span4Mux_v I__10943 (
            .O(N__48833),
            .I(N__48824));
    Span4Mux_v I__10942 (
            .O(N__48830),
            .I(N__48821));
    Odrv12 I__10941 (
            .O(N__48827),
            .I(n14_adj_1608));
    Odrv4 I__10940 (
            .O(N__48824),
            .I(n14_adj_1608));
    Odrv4 I__10939 (
            .O(N__48821),
            .I(n14_adj_1608));
    InMux I__10938 (
            .O(N__48814),
            .I(N__48811));
    LocalMux I__10937 (
            .O(N__48811),
            .I(N__48804));
    InMux I__10936 (
            .O(N__48810),
            .I(N__48801));
    InMux I__10935 (
            .O(N__48809),
            .I(N__48791));
    InMux I__10934 (
            .O(N__48808),
            .I(N__48791));
    InMux I__10933 (
            .O(N__48807),
            .I(N__48791));
    Span4Mux_v I__10932 (
            .O(N__48804),
            .I(N__48786));
    LocalMux I__10931 (
            .O(N__48801),
            .I(N__48786));
    InMux I__10930 (
            .O(N__48800),
            .I(N__48783));
    InMux I__10929 (
            .O(N__48799),
            .I(N__48780));
    InMux I__10928 (
            .O(N__48798),
            .I(N__48777));
    LocalMux I__10927 (
            .O(N__48791),
            .I(N__48774));
    Span4Mux_v I__10926 (
            .O(N__48786),
            .I(N__48771));
    LocalMux I__10925 (
            .O(N__48783),
            .I(N__48768));
    LocalMux I__10924 (
            .O(N__48780),
            .I(N__48765));
    LocalMux I__10923 (
            .O(N__48777),
            .I(N__48762));
    Span4Mux_v I__10922 (
            .O(N__48774),
            .I(N__48759));
    Span4Mux_v I__10921 (
            .O(N__48771),
            .I(N__48754));
    Span4Mux_v I__10920 (
            .O(N__48768),
            .I(N__48754));
    Span4Mux_h I__10919 (
            .O(N__48765),
            .I(N__48751));
    Span4Mux_v I__10918 (
            .O(N__48762),
            .I(N__48748));
    Sp12to4 I__10917 (
            .O(N__48759),
            .I(N__48745));
    Sp12to4 I__10916 (
            .O(N__48754),
            .I(N__48742));
    Sp12to4 I__10915 (
            .O(N__48751),
            .I(N__48739));
    Sp12to4 I__10914 (
            .O(N__48748),
            .I(N__48734));
    Span12Mux_h I__10913 (
            .O(N__48745),
            .I(N__48734));
    Span12Mux_h I__10912 (
            .O(N__48742),
            .I(N__48731));
    Odrv12 I__10911 (
            .O(N__48739),
            .I(n13129));
    Odrv12 I__10910 (
            .O(N__48734),
            .I(n13129));
    Odrv12 I__10909 (
            .O(N__48731),
            .I(n13129));
    CascadeMux I__10908 (
            .O(N__48724),
            .I(N__48721));
    InMux I__10907 (
            .O(N__48721),
            .I(N__48716));
    InMux I__10906 (
            .O(N__48720),
            .I(N__48713));
    InMux I__10905 (
            .O(N__48719),
            .I(N__48710));
    LocalMux I__10904 (
            .O(N__48716),
            .I(N__48707));
    LocalMux I__10903 (
            .O(N__48713),
            .I(N__48699));
    LocalMux I__10902 (
            .O(N__48710),
            .I(N__48699));
    Sp12to4 I__10901 (
            .O(N__48707),
            .I(N__48699));
    InMux I__10900 (
            .O(N__48706),
            .I(N__48696));
    Span12Mux_v I__10899 (
            .O(N__48699),
            .I(N__48693));
    LocalMux I__10898 (
            .O(N__48696),
            .I(N__48689));
    Span12Mux_h I__10897 (
            .O(N__48693),
            .I(N__48686));
    InMux I__10896 (
            .O(N__48692),
            .I(N__48683));
    Span4Mux_h I__10895 (
            .O(N__48689),
            .I(N__48680));
    Odrv12 I__10894 (
            .O(N__48686),
            .I(buf_cfgRTD_0));
    LocalMux I__10893 (
            .O(N__48683),
            .I(buf_cfgRTD_0));
    Odrv4 I__10892 (
            .O(N__48680),
            .I(buf_cfgRTD_0));
    CascadeMux I__10891 (
            .O(N__48673),
            .I(N__48670));
    InMux I__10890 (
            .O(N__48670),
            .I(N__48667));
    LocalMux I__10889 (
            .O(N__48667),
            .I(N__48664));
    Span4Mux_h I__10888 (
            .O(N__48664),
            .I(N__48661));
    Odrv4 I__10887 (
            .O(N__48661),
            .I(n22238));
    CascadeMux I__10886 (
            .O(N__48658),
            .I(n22240_cascade_));
    InMux I__10885 (
            .O(N__48655),
            .I(N__48652));
    LocalMux I__10884 (
            .O(N__48652),
            .I(n23053));
    CascadeMux I__10883 (
            .O(N__48649),
            .I(n11280_cascade_));
    CascadeMux I__10882 (
            .O(N__48646),
            .I(n12509_cascade_));
    InMux I__10881 (
            .O(N__48643),
            .I(N__48639));
    InMux I__10880 (
            .O(N__48642),
            .I(N__48636));
    LocalMux I__10879 (
            .O(N__48639),
            .I(N__48633));
    LocalMux I__10878 (
            .O(N__48636),
            .I(comm_length_2));
    Odrv4 I__10877 (
            .O(N__48633),
            .I(comm_length_2));
    CascadeMux I__10876 (
            .O(N__48628),
            .I(N__48625));
    InMux I__10875 (
            .O(N__48625),
            .I(N__48622));
    LocalMux I__10874 (
            .O(N__48622),
            .I(N__48619));
    Span4Mux_h I__10873 (
            .O(N__48619),
            .I(N__48616));
    Odrv4 I__10872 (
            .O(N__48616),
            .I(comm_length_0));
    InMux I__10871 (
            .O(N__48613),
            .I(N__48610));
    LocalMux I__10870 (
            .O(N__48610),
            .I(N__48606));
    InMux I__10869 (
            .O(N__48609),
            .I(N__48603));
    Span4Mux_h I__10868 (
            .O(N__48606),
            .I(N__48597));
    LocalMux I__10867 (
            .O(N__48603),
            .I(N__48597));
    InMux I__10866 (
            .O(N__48602),
            .I(N__48594));
    Span4Mux_h I__10865 (
            .O(N__48597),
            .I(N__48591));
    LocalMux I__10864 (
            .O(N__48594),
            .I(buf_adcdata_vac_17));
    Odrv4 I__10863 (
            .O(N__48591),
            .I(buf_adcdata_vac_17));
    InMux I__10862 (
            .O(N__48586),
            .I(N__48583));
    LocalMux I__10861 (
            .O(N__48583),
            .I(N__48580));
    Span4Mux_h I__10860 (
            .O(N__48580),
            .I(N__48577));
    Odrv4 I__10859 (
            .O(N__48577),
            .I(n23486));
    CascadeMux I__10858 (
            .O(N__48574),
            .I(N__48571));
    InMux I__10857 (
            .O(N__48571),
            .I(N__48568));
    LocalMux I__10856 (
            .O(N__48568),
            .I(N__48565));
    Span4Mux_v I__10855 (
            .O(N__48565),
            .I(N__48562));
    Span4Mux_h I__10854 (
            .O(N__48562),
            .I(N__48558));
    CascadeMux I__10853 (
            .O(N__48561),
            .I(N__48555));
    Span4Mux_h I__10852 (
            .O(N__48558),
            .I(N__48552));
    InMux I__10851 (
            .O(N__48555),
            .I(N__48549));
    Odrv4 I__10850 (
            .O(N__48552),
            .I(buf_adcdata_vdc_17));
    LocalMux I__10849 (
            .O(N__48549),
            .I(buf_adcdata_vdc_17));
    InMux I__10848 (
            .O(N__48544),
            .I(N__48523));
    InMux I__10847 (
            .O(N__48543),
            .I(N__48523));
    InMux I__10846 (
            .O(N__48542),
            .I(N__48523));
    InMux I__10845 (
            .O(N__48541),
            .I(N__48523));
    InMux I__10844 (
            .O(N__48540),
            .I(N__48514));
    InMux I__10843 (
            .O(N__48539),
            .I(N__48514));
    InMux I__10842 (
            .O(N__48538),
            .I(N__48514));
    InMux I__10841 (
            .O(N__48537),
            .I(N__48514));
    InMux I__10840 (
            .O(N__48536),
            .I(N__48493));
    InMux I__10839 (
            .O(N__48535),
            .I(N__48493));
    InMux I__10838 (
            .O(N__48534),
            .I(N__48493));
    InMux I__10837 (
            .O(N__48533),
            .I(N__48493));
    InMux I__10836 (
            .O(N__48532),
            .I(N__48490));
    LocalMux I__10835 (
            .O(N__48523),
            .I(N__48487));
    LocalMux I__10834 (
            .O(N__48514),
            .I(N__48484));
    InMux I__10833 (
            .O(N__48513),
            .I(N__48475));
    InMux I__10832 (
            .O(N__48512),
            .I(N__48475));
    InMux I__10831 (
            .O(N__48511),
            .I(N__48475));
    InMux I__10830 (
            .O(N__48510),
            .I(N__48475));
    InMux I__10829 (
            .O(N__48509),
            .I(N__48466));
    InMux I__10828 (
            .O(N__48508),
            .I(N__48466));
    InMux I__10827 (
            .O(N__48507),
            .I(N__48466));
    InMux I__10826 (
            .O(N__48506),
            .I(N__48466));
    InMux I__10825 (
            .O(N__48505),
            .I(N__48457));
    InMux I__10824 (
            .O(N__48504),
            .I(N__48457));
    InMux I__10823 (
            .O(N__48503),
            .I(N__48457));
    InMux I__10822 (
            .O(N__48502),
            .I(N__48457));
    LocalMux I__10821 (
            .O(N__48493),
            .I(N__48452));
    LocalMux I__10820 (
            .O(N__48490),
            .I(N__48452));
    Odrv4 I__10819 (
            .O(N__48487),
            .I(n49));
    Odrv4 I__10818 (
            .O(N__48484),
            .I(n49));
    LocalMux I__10817 (
            .O(N__48475),
            .I(n49));
    LocalMux I__10816 (
            .O(N__48466),
            .I(n49));
    LocalMux I__10815 (
            .O(N__48457),
            .I(n49));
    Odrv4 I__10814 (
            .O(N__48452),
            .I(n49));
    InMux I__10813 (
            .O(N__48439),
            .I(bfn_17_8_0_));
    InMux I__10812 (
            .O(N__48436),
            .I(N__48432));
    InMux I__10811 (
            .O(N__48435),
            .I(N__48429));
    LocalMux I__10810 (
            .O(N__48432),
            .I(N__48426));
    LocalMux I__10809 (
            .O(N__48429),
            .I(wdtick_cnt_24));
    Odrv4 I__10808 (
            .O(N__48426),
            .I(wdtick_cnt_24));
    InMux I__10807 (
            .O(N__48421),
            .I(N__48418));
    LocalMux I__10806 (
            .O(N__48418),
            .I(N__48397));
    ClkMux I__10805 (
            .O(N__48417),
            .I(N__48352));
    ClkMux I__10804 (
            .O(N__48416),
            .I(N__48352));
    ClkMux I__10803 (
            .O(N__48415),
            .I(N__48352));
    ClkMux I__10802 (
            .O(N__48414),
            .I(N__48352));
    ClkMux I__10801 (
            .O(N__48413),
            .I(N__48352));
    ClkMux I__10800 (
            .O(N__48412),
            .I(N__48352));
    ClkMux I__10799 (
            .O(N__48411),
            .I(N__48352));
    ClkMux I__10798 (
            .O(N__48410),
            .I(N__48352));
    ClkMux I__10797 (
            .O(N__48409),
            .I(N__48352));
    ClkMux I__10796 (
            .O(N__48408),
            .I(N__48352));
    ClkMux I__10795 (
            .O(N__48407),
            .I(N__48352));
    ClkMux I__10794 (
            .O(N__48406),
            .I(N__48352));
    ClkMux I__10793 (
            .O(N__48405),
            .I(N__48352));
    ClkMux I__10792 (
            .O(N__48404),
            .I(N__48352));
    ClkMux I__10791 (
            .O(N__48403),
            .I(N__48352));
    ClkMux I__10790 (
            .O(N__48402),
            .I(N__48352));
    ClkMux I__10789 (
            .O(N__48401),
            .I(N__48352));
    ClkMux I__10788 (
            .O(N__48400),
            .I(N__48352));
    Glb2LocalMux I__10787 (
            .O(N__48397),
            .I(N__48352));
    ClkMux I__10786 (
            .O(N__48396),
            .I(N__48352));
    ClkMux I__10785 (
            .O(N__48395),
            .I(N__48352));
    GlobalMux I__10784 (
            .O(N__48352),
            .I(DDS_MCLK1));
    CEMux I__10783 (
            .O(N__48349),
            .I(N__48346));
    LocalMux I__10782 (
            .O(N__48346),
            .I(N__48342));
    CEMux I__10781 (
            .O(N__48345),
            .I(N__48339));
    Span4Mux_v I__10780 (
            .O(N__48342),
            .I(N__48332));
    LocalMux I__10779 (
            .O(N__48339),
            .I(N__48332));
    CEMux I__10778 (
            .O(N__48338),
            .I(N__48329));
    CEMux I__10777 (
            .O(N__48337),
            .I(N__48326));
    Span4Mux_v I__10776 (
            .O(N__48332),
            .I(N__48323));
    LocalMux I__10775 (
            .O(N__48329),
            .I(N__48320));
    LocalMux I__10774 (
            .O(N__48326),
            .I(N__48317));
    Span4Mux_h I__10773 (
            .O(N__48323),
            .I(N__48314));
    Span4Mux_h I__10772 (
            .O(N__48320),
            .I(N__48311));
    Span4Mux_h I__10771 (
            .O(N__48317),
            .I(N__48308));
    Odrv4 I__10770 (
            .O(N__48314),
            .I(n12366));
    Odrv4 I__10769 (
            .O(N__48311),
            .I(n12366));
    Odrv4 I__10768 (
            .O(N__48308),
            .I(n12366));
    InMux I__10767 (
            .O(N__48301),
            .I(N__48298));
    LocalMux I__10766 (
            .O(N__48298),
            .I(n7_adj_1757));
    CascadeMux I__10765 (
            .O(N__48295),
            .I(n2562_cascade_));
    SRMux I__10764 (
            .O(N__48292),
            .I(N__48288));
    SRMux I__10763 (
            .O(N__48291),
            .I(N__48285));
    LocalMux I__10762 (
            .O(N__48288),
            .I(N__48282));
    LocalMux I__10761 (
            .O(N__48285),
            .I(N__48279));
    Span4Mux_v I__10760 (
            .O(N__48282),
            .I(N__48276));
    Odrv12 I__10759 (
            .O(N__48279),
            .I(n15378));
    Odrv4 I__10758 (
            .O(N__48276),
            .I(n15378));
    CascadeMux I__10757 (
            .O(N__48271),
            .I(N__48268));
    InMux I__10756 (
            .O(N__48268),
            .I(N__48265));
    LocalMux I__10755 (
            .O(N__48265),
            .I(n8_adj_1782));
    CEMux I__10754 (
            .O(N__48262),
            .I(N__48259));
    LocalMux I__10753 (
            .O(N__48259),
            .I(N__48256));
    Span4Mux_v I__10752 (
            .O(N__48256),
            .I(N__48253));
    Odrv4 I__10751 (
            .O(N__48253),
            .I(n12540));
    InMux I__10750 (
            .O(N__48250),
            .I(N__48247));
    LocalMux I__10749 (
            .O(N__48247),
            .I(N__48244));
    Span4Mux_h I__10748 (
            .O(N__48244),
            .I(N__48241));
    Span4Mux_v I__10747 (
            .O(N__48241),
            .I(N__48238));
    Odrv4 I__10746 (
            .O(N__48238),
            .I(n14_adj_1606));
    InMux I__10745 (
            .O(N__48235),
            .I(N__48231));
    InMux I__10744 (
            .O(N__48234),
            .I(N__48228));
    LocalMux I__10743 (
            .O(N__48231),
            .I(N__48225));
    LocalMux I__10742 (
            .O(N__48228),
            .I(wdtick_cnt_16));
    Odrv4 I__10741 (
            .O(N__48225),
            .I(wdtick_cnt_16));
    InMux I__10740 (
            .O(N__48220),
            .I(bfn_17_7_0_));
    InMux I__10739 (
            .O(N__48217),
            .I(N__48213));
    InMux I__10738 (
            .O(N__48216),
            .I(N__48210));
    LocalMux I__10737 (
            .O(N__48213),
            .I(wdtick_cnt_17));
    LocalMux I__10736 (
            .O(N__48210),
            .I(wdtick_cnt_17));
    InMux I__10735 (
            .O(N__48205),
            .I(n20782));
    InMux I__10734 (
            .O(N__48202),
            .I(N__48198));
    InMux I__10733 (
            .O(N__48201),
            .I(N__48195));
    LocalMux I__10732 (
            .O(N__48198),
            .I(N__48192));
    LocalMux I__10731 (
            .O(N__48195),
            .I(wdtick_cnt_18));
    Odrv4 I__10730 (
            .O(N__48192),
            .I(wdtick_cnt_18));
    InMux I__10729 (
            .O(N__48187),
            .I(n20783));
    CascadeMux I__10728 (
            .O(N__48184),
            .I(N__48180));
    InMux I__10727 (
            .O(N__48183),
            .I(N__48177));
    InMux I__10726 (
            .O(N__48180),
            .I(N__48174));
    LocalMux I__10725 (
            .O(N__48177),
            .I(wdtick_cnt_19));
    LocalMux I__10724 (
            .O(N__48174),
            .I(wdtick_cnt_19));
    InMux I__10723 (
            .O(N__48169),
            .I(n20784));
    InMux I__10722 (
            .O(N__48166),
            .I(N__48162));
    InMux I__10721 (
            .O(N__48165),
            .I(N__48159));
    LocalMux I__10720 (
            .O(N__48162),
            .I(wdtick_cnt_20));
    LocalMux I__10719 (
            .O(N__48159),
            .I(wdtick_cnt_20));
    InMux I__10718 (
            .O(N__48154),
            .I(n20785));
    InMux I__10717 (
            .O(N__48151),
            .I(N__48147));
    InMux I__10716 (
            .O(N__48150),
            .I(N__48144));
    LocalMux I__10715 (
            .O(N__48147),
            .I(wdtick_cnt_21));
    LocalMux I__10714 (
            .O(N__48144),
            .I(wdtick_cnt_21));
    InMux I__10713 (
            .O(N__48139),
            .I(n20786));
    InMux I__10712 (
            .O(N__48136),
            .I(N__48132));
    InMux I__10711 (
            .O(N__48135),
            .I(N__48129));
    LocalMux I__10710 (
            .O(N__48132),
            .I(wdtick_cnt_22));
    LocalMux I__10709 (
            .O(N__48129),
            .I(wdtick_cnt_22));
    InMux I__10708 (
            .O(N__48124),
            .I(n20787));
    InMux I__10707 (
            .O(N__48121),
            .I(N__48117));
    InMux I__10706 (
            .O(N__48120),
            .I(N__48114));
    LocalMux I__10705 (
            .O(N__48117),
            .I(wdtick_cnt_23));
    LocalMux I__10704 (
            .O(N__48114),
            .I(wdtick_cnt_23));
    InMux I__10703 (
            .O(N__48109),
            .I(n20788));
    CascadeMux I__10702 (
            .O(N__48106),
            .I(N__48103));
    InMux I__10701 (
            .O(N__48103),
            .I(N__48100));
    LocalMux I__10700 (
            .O(N__48100),
            .I(N__48096));
    InMux I__10699 (
            .O(N__48099),
            .I(N__48093));
    Odrv4 I__10698 (
            .O(N__48096),
            .I(wdtick_cnt_7));
    LocalMux I__10697 (
            .O(N__48093),
            .I(wdtick_cnt_7));
    InMux I__10696 (
            .O(N__48088),
            .I(n20772));
    InMux I__10695 (
            .O(N__48085),
            .I(N__48081));
    InMux I__10694 (
            .O(N__48084),
            .I(N__48078));
    LocalMux I__10693 (
            .O(N__48081),
            .I(N__48075));
    LocalMux I__10692 (
            .O(N__48078),
            .I(wdtick_cnt_8));
    Odrv4 I__10691 (
            .O(N__48075),
            .I(wdtick_cnt_8));
    InMux I__10690 (
            .O(N__48070),
            .I(bfn_17_6_0_));
    InMux I__10689 (
            .O(N__48067),
            .I(N__48063));
    InMux I__10688 (
            .O(N__48066),
            .I(N__48060));
    LocalMux I__10687 (
            .O(N__48063),
            .I(wdtick_cnt_9));
    LocalMux I__10686 (
            .O(N__48060),
            .I(wdtick_cnt_9));
    InMux I__10685 (
            .O(N__48055),
            .I(n20774));
    InMux I__10684 (
            .O(N__48052),
            .I(N__48048));
    InMux I__10683 (
            .O(N__48051),
            .I(N__48045));
    LocalMux I__10682 (
            .O(N__48048),
            .I(wdtick_cnt_10));
    LocalMux I__10681 (
            .O(N__48045),
            .I(wdtick_cnt_10));
    InMux I__10680 (
            .O(N__48040),
            .I(n20775));
    InMux I__10679 (
            .O(N__48037),
            .I(N__48033));
    InMux I__10678 (
            .O(N__48036),
            .I(N__48030));
    LocalMux I__10677 (
            .O(N__48033),
            .I(wdtick_cnt_11));
    LocalMux I__10676 (
            .O(N__48030),
            .I(wdtick_cnt_11));
    InMux I__10675 (
            .O(N__48025),
            .I(n20776));
    InMux I__10674 (
            .O(N__48022),
            .I(N__48018));
    InMux I__10673 (
            .O(N__48021),
            .I(N__48015));
    LocalMux I__10672 (
            .O(N__48018),
            .I(wdtick_cnt_12));
    LocalMux I__10671 (
            .O(N__48015),
            .I(wdtick_cnt_12));
    InMux I__10670 (
            .O(N__48010),
            .I(n20777));
    InMux I__10669 (
            .O(N__48007),
            .I(N__48003));
    InMux I__10668 (
            .O(N__48006),
            .I(N__48000));
    LocalMux I__10667 (
            .O(N__48003),
            .I(wdtick_cnt_13));
    LocalMux I__10666 (
            .O(N__48000),
            .I(wdtick_cnt_13));
    InMux I__10665 (
            .O(N__47995),
            .I(n20778));
    InMux I__10664 (
            .O(N__47992),
            .I(N__47988));
    InMux I__10663 (
            .O(N__47991),
            .I(N__47985));
    LocalMux I__10662 (
            .O(N__47988),
            .I(N__47980));
    LocalMux I__10661 (
            .O(N__47985),
            .I(N__47980));
    Odrv4 I__10660 (
            .O(N__47980),
            .I(wdtick_cnt_14));
    InMux I__10659 (
            .O(N__47977),
            .I(n20779));
    InMux I__10658 (
            .O(N__47974),
            .I(N__47970));
    InMux I__10657 (
            .O(N__47973),
            .I(N__47967));
    LocalMux I__10656 (
            .O(N__47970),
            .I(wdtick_cnt_15));
    LocalMux I__10655 (
            .O(N__47967),
            .I(wdtick_cnt_15));
    InMux I__10654 (
            .O(N__47962),
            .I(n20780));
    InMux I__10653 (
            .O(N__47959),
            .I(N__47955));
    InMux I__10652 (
            .O(N__47958),
            .I(N__47951));
    LocalMux I__10651 (
            .O(N__47955),
            .I(N__47948));
    InMux I__10650 (
            .O(N__47954),
            .I(N__47945));
    LocalMux I__10649 (
            .O(N__47951),
            .I(\comm_spi.n15330 ));
    Odrv4 I__10648 (
            .O(N__47948),
            .I(\comm_spi.n15330 ));
    LocalMux I__10647 (
            .O(N__47945),
            .I(\comm_spi.n15330 ));
    InMux I__10646 (
            .O(N__47938),
            .I(N__47934));
    InMux I__10645 (
            .O(N__47937),
            .I(N__47931));
    LocalMux I__10644 (
            .O(N__47934),
            .I(N__47926));
    LocalMux I__10643 (
            .O(N__47931),
            .I(N__47926));
    Odrv4 I__10642 (
            .O(N__47926),
            .I(wdtick_cnt_0));
    InMux I__10641 (
            .O(N__47923),
            .I(bfn_17_5_0_));
    InMux I__10640 (
            .O(N__47920),
            .I(N__47916));
    InMux I__10639 (
            .O(N__47919),
            .I(N__47913));
    LocalMux I__10638 (
            .O(N__47916),
            .I(wdtick_cnt_1));
    LocalMux I__10637 (
            .O(N__47913),
            .I(wdtick_cnt_1));
    InMux I__10636 (
            .O(N__47908),
            .I(n20766));
    InMux I__10635 (
            .O(N__47905),
            .I(N__47901));
    InMux I__10634 (
            .O(N__47904),
            .I(N__47898));
    LocalMux I__10633 (
            .O(N__47901),
            .I(wdtick_cnt_2));
    LocalMux I__10632 (
            .O(N__47898),
            .I(wdtick_cnt_2));
    InMux I__10631 (
            .O(N__47893),
            .I(n20767));
    CascadeMux I__10630 (
            .O(N__47890),
            .I(N__47887));
    InMux I__10629 (
            .O(N__47887),
            .I(N__47884));
    LocalMux I__10628 (
            .O(N__47884),
            .I(N__47880));
    InMux I__10627 (
            .O(N__47883),
            .I(N__47877));
    Odrv4 I__10626 (
            .O(N__47880),
            .I(wdtick_cnt_3));
    LocalMux I__10625 (
            .O(N__47877),
            .I(wdtick_cnt_3));
    InMux I__10624 (
            .O(N__47872),
            .I(n20768));
    InMux I__10623 (
            .O(N__47869),
            .I(N__47865));
    InMux I__10622 (
            .O(N__47868),
            .I(N__47862));
    LocalMux I__10621 (
            .O(N__47865),
            .I(wdtick_cnt_4));
    LocalMux I__10620 (
            .O(N__47862),
            .I(wdtick_cnt_4));
    InMux I__10619 (
            .O(N__47857),
            .I(n20769));
    CascadeMux I__10618 (
            .O(N__47854),
            .I(N__47851));
    InMux I__10617 (
            .O(N__47851),
            .I(N__47848));
    LocalMux I__10616 (
            .O(N__47848),
            .I(N__47844));
    InMux I__10615 (
            .O(N__47847),
            .I(N__47841));
    Odrv4 I__10614 (
            .O(N__47844),
            .I(wdtick_cnt_5));
    LocalMux I__10613 (
            .O(N__47841),
            .I(wdtick_cnt_5));
    InMux I__10612 (
            .O(N__47836),
            .I(n20770));
    CascadeMux I__10611 (
            .O(N__47833),
            .I(N__47829));
    InMux I__10610 (
            .O(N__47832),
            .I(N__47826));
    InMux I__10609 (
            .O(N__47829),
            .I(N__47823));
    LocalMux I__10608 (
            .O(N__47826),
            .I(wdtick_cnt_6));
    LocalMux I__10607 (
            .O(N__47823),
            .I(wdtick_cnt_6));
    InMux I__10606 (
            .O(N__47818),
            .I(n20771));
    InMux I__10605 (
            .O(N__47815),
            .I(N__47810));
    InMux I__10604 (
            .O(N__47814),
            .I(N__47807));
    InMux I__10603 (
            .O(N__47813),
            .I(N__47804));
    LocalMux I__10602 (
            .O(N__47810),
            .I(N__47799));
    LocalMux I__10601 (
            .O(N__47807),
            .I(N__47799));
    LocalMux I__10600 (
            .O(N__47804),
            .I(N__47796));
    Span4Mux_h I__10599 (
            .O(N__47799),
            .I(N__47793));
    Odrv4 I__10598 (
            .O(N__47796),
            .I(data_index_0));
    Odrv4 I__10597 (
            .O(N__47793),
            .I(data_index_0));
    InMux I__10596 (
            .O(N__47788),
            .I(N__47785));
    LocalMux I__10595 (
            .O(N__47785),
            .I(N__47780));
    CascadeMux I__10594 (
            .O(N__47784),
            .I(N__47777));
    CascadeMux I__10593 (
            .O(N__47783),
            .I(N__47766));
    Span4Mux_v I__10592 (
            .O(N__47780),
            .I(N__47763));
    InMux I__10591 (
            .O(N__47777),
            .I(N__47760));
    CascadeMux I__10590 (
            .O(N__47776),
            .I(N__47757));
    CascadeMux I__10589 (
            .O(N__47775),
            .I(N__47754));
    CascadeMux I__10588 (
            .O(N__47774),
            .I(N__47751));
    CascadeMux I__10587 (
            .O(N__47773),
            .I(N__47748));
    CascadeMux I__10586 (
            .O(N__47772),
            .I(N__47745));
    CascadeMux I__10585 (
            .O(N__47771),
            .I(N__47742));
    CascadeMux I__10584 (
            .O(N__47770),
            .I(N__47739));
    CascadeMux I__10583 (
            .O(N__47769),
            .I(N__47736));
    InMux I__10582 (
            .O(N__47766),
            .I(N__47733));
    Span4Mux_h I__10581 (
            .O(N__47763),
            .I(N__47728));
    LocalMux I__10580 (
            .O(N__47760),
            .I(N__47728));
    InMux I__10579 (
            .O(N__47757),
            .I(N__47719));
    InMux I__10578 (
            .O(N__47754),
            .I(N__47719));
    InMux I__10577 (
            .O(N__47751),
            .I(N__47719));
    InMux I__10576 (
            .O(N__47748),
            .I(N__47719));
    InMux I__10575 (
            .O(N__47745),
            .I(N__47710));
    InMux I__10574 (
            .O(N__47742),
            .I(N__47710));
    InMux I__10573 (
            .O(N__47739),
            .I(N__47710));
    InMux I__10572 (
            .O(N__47736),
            .I(N__47710));
    LocalMux I__10571 (
            .O(N__47733),
            .I(N__47707));
    Span4Mux_v I__10570 (
            .O(N__47728),
            .I(N__47704));
    LocalMux I__10569 (
            .O(N__47719),
            .I(N__47699));
    LocalMux I__10568 (
            .O(N__47710),
            .I(N__47699));
    Odrv12 I__10567 (
            .O(N__47707),
            .I(n11254));
    Odrv4 I__10566 (
            .O(N__47704),
            .I(n11254));
    Odrv4 I__10565 (
            .O(N__47699),
            .I(n11254));
    CEMux I__10564 (
            .O(N__47692),
            .I(N__47688));
    CEMux I__10563 (
            .O(N__47691),
            .I(N__47685));
    LocalMux I__10562 (
            .O(N__47688),
            .I(N__47682));
    LocalMux I__10561 (
            .O(N__47685),
            .I(N__47679));
    Odrv12 I__10560 (
            .O(N__47682),
            .I(n13052));
    Odrv4 I__10559 (
            .O(N__47679),
            .I(n13052));
    SRMux I__10558 (
            .O(N__47674),
            .I(N__47671));
    LocalMux I__10557 (
            .O(N__47671),
            .I(N__47668));
    Odrv4 I__10556 (
            .O(N__47668),
            .I(n15562));
    CascadeMux I__10555 (
            .O(N__47665),
            .I(n15562_cascade_));
    InMux I__10554 (
            .O(N__47662),
            .I(N__47656));
    InMux I__10553 (
            .O(N__47661),
            .I(N__47648));
    InMux I__10552 (
            .O(N__47660),
            .I(N__47648));
    InMux I__10551 (
            .O(N__47659),
            .I(N__47648));
    LocalMux I__10550 (
            .O(N__47656),
            .I(N__47645));
    InMux I__10549 (
            .O(N__47655),
            .I(N__47642));
    LocalMux I__10548 (
            .O(N__47648),
            .I(N__47637));
    Span4Mux_h I__10547 (
            .O(N__47645),
            .I(N__47637));
    LocalMux I__10546 (
            .O(N__47642),
            .I(bit_cnt_0));
    Odrv4 I__10545 (
            .O(N__47637),
            .I(bit_cnt_0));
    CEMux I__10544 (
            .O(N__47632),
            .I(N__47629));
    LocalMux I__10543 (
            .O(N__47629),
            .I(N__47626));
    Span4Mux_v I__10542 (
            .O(N__47626),
            .I(N__47622));
    CEMux I__10541 (
            .O(N__47625),
            .I(N__47619));
    Odrv4 I__10540 (
            .O(N__47622),
            .I(\SIG_DDS.n9 ));
    LocalMux I__10539 (
            .O(N__47619),
            .I(\SIG_DDS.n9 ));
    IoInMux I__10538 (
            .O(N__47614),
            .I(N__47611));
    LocalMux I__10537 (
            .O(N__47611),
            .I(N__47608));
    Span4Mux_s2_v I__10536 (
            .O(N__47608),
            .I(N__47605));
    Span4Mux_h I__10535 (
            .O(N__47605),
            .I(N__47602));
    Span4Mux_h I__10534 (
            .O(N__47602),
            .I(N__47598));
    CascadeMux I__10533 (
            .O(N__47601),
            .I(N__47595));
    Span4Mux_v I__10532 (
            .O(N__47598),
            .I(N__47592));
    InMux I__10531 (
            .O(N__47595),
            .I(N__47589));
    Odrv4 I__10530 (
            .O(N__47592),
            .I(DDS_SCK));
    LocalMux I__10529 (
            .O(N__47589),
            .I(DDS_SCK));
    CascadeMux I__10528 (
            .O(N__47584),
            .I(N__47579));
    CascadeMux I__10527 (
            .O(N__47583),
            .I(N__47576));
    CascadeMux I__10526 (
            .O(N__47582),
            .I(N__47572));
    InMux I__10525 (
            .O(N__47579),
            .I(N__47569));
    InMux I__10524 (
            .O(N__47576),
            .I(N__47566));
    InMux I__10523 (
            .O(N__47575),
            .I(N__47563));
    InMux I__10522 (
            .O(N__47572),
            .I(N__47560));
    LocalMux I__10521 (
            .O(N__47569),
            .I(N__47555));
    LocalMux I__10520 (
            .O(N__47566),
            .I(N__47555));
    LocalMux I__10519 (
            .O(N__47563),
            .I(N__47550));
    LocalMux I__10518 (
            .O(N__47560),
            .I(N__47550));
    Span12Mux_h I__10517 (
            .O(N__47555),
            .I(N__47547));
    Odrv12 I__10516 (
            .O(N__47550),
            .I(trig_dds0));
    Odrv12 I__10515 (
            .O(N__47547),
            .I(trig_dds0));
    InMux I__10514 (
            .O(N__47542),
            .I(N__47538));
    InMux I__10513 (
            .O(N__47541),
            .I(N__47535));
    LocalMux I__10512 (
            .O(N__47538),
            .I(\comm_spi.imosi ));
    LocalMux I__10511 (
            .O(N__47535),
            .I(\comm_spi.imosi ));
    SRMux I__10510 (
            .O(N__47530),
            .I(N__47527));
    LocalMux I__10509 (
            .O(N__47527),
            .I(N__47524));
    Odrv4 I__10508 (
            .O(N__47524),
            .I(\comm_spi.DOUT_7__N_834 ));
    InMux I__10507 (
            .O(N__47521),
            .I(N__47518));
    LocalMux I__10506 (
            .O(N__47518),
            .I(N__47512));
    InMux I__10505 (
            .O(N__47517),
            .I(N__47509));
    InMux I__10504 (
            .O(N__47516),
            .I(N__47506));
    InMux I__10503 (
            .O(N__47515),
            .I(N__47503));
    Span4Mux_h I__10502 (
            .O(N__47512),
            .I(N__47498));
    LocalMux I__10501 (
            .O(N__47509),
            .I(N__47498));
    LocalMux I__10500 (
            .O(N__47506),
            .I(N__47495));
    LocalMux I__10499 (
            .O(N__47503),
            .I(N__47492));
    Span4Mux_h I__10498 (
            .O(N__47498),
            .I(N__47489));
    Span4Mux_h I__10497 (
            .O(N__47495),
            .I(N__47486));
    Odrv12 I__10496 (
            .O(N__47492),
            .I(n14_adj_1609));
    Odrv4 I__10495 (
            .O(N__47489),
            .I(n14_adj_1609));
    Odrv4 I__10494 (
            .O(N__47486),
            .I(n14_adj_1609));
    InMux I__10493 (
            .O(N__47479),
            .I(n20667));
    InMux I__10492 (
            .O(N__47476),
            .I(N__47472));
    InMux I__10491 (
            .O(N__47475),
            .I(N__47469));
    LocalMux I__10490 (
            .O(N__47472),
            .I(N__47466));
    LocalMux I__10489 (
            .O(N__47469),
            .I(data_idxvec_8));
    Odrv4 I__10488 (
            .O(N__47466),
            .I(data_idxvec_8));
    InMux I__10487 (
            .O(N__47461),
            .I(bfn_16_17_0_));
    InMux I__10486 (
            .O(N__47458),
            .I(n20669));
    InMux I__10485 (
            .O(N__47455),
            .I(N__47446));
    InMux I__10484 (
            .O(N__47454),
            .I(N__47446));
    CascadeMux I__10483 (
            .O(N__47453),
            .I(N__47443));
    InMux I__10482 (
            .O(N__47452),
            .I(N__47440));
    InMux I__10481 (
            .O(N__47451),
            .I(N__47437));
    LocalMux I__10480 (
            .O(N__47446),
            .I(N__47434));
    InMux I__10479 (
            .O(N__47443),
            .I(N__47431));
    LocalMux I__10478 (
            .O(N__47440),
            .I(N__47428));
    LocalMux I__10477 (
            .O(N__47437),
            .I(N__47425));
    Span4Mux_h I__10476 (
            .O(N__47434),
            .I(N__47419));
    LocalMux I__10475 (
            .O(N__47431),
            .I(N__47419));
    Span4Mux_v I__10474 (
            .O(N__47428),
            .I(N__47416));
    Span4Mux_v I__10473 (
            .O(N__47425),
            .I(N__47413));
    InMux I__10472 (
            .O(N__47424),
            .I(N__47410));
    Span4Mux_v I__10471 (
            .O(N__47419),
            .I(N__47407));
    Span4Mux_h I__10470 (
            .O(N__47416),
            .I(N__47402));
    Span4Mux_v I__10469 (
            .O(N__47413),
            .I(N__47402));
    LocalMux I__10468 (
            .O(N__47410),
            .I(N__47397));
    Span4Mux_h I__10467 (
            .O(N__47407),
            .I(N__47397));
    Odrv4 I__10466 (
            .O(N__47402),
            .I(n14_adj_1655));
    Odrv4 I__10465 (
            .O(N__47397),
            .I(n14_adj_1655));
    InMux I__10464 (
            .O(N__47392),
            .I(N__47388));
    InMux I__10463 (
            .O(N__47391),
            .I(N__47385));
    LocalMux I__10462 (
            .O(N__47388),
            .I(data_idxvec_10));
    LocalMux I__10461 (
            .O(N__47385),
            .I(data_idxvec_10));
    InMux I__10460 (
            .O(N__47380),
            .I(n20670));
    InMux I__10459 (
            .O(N__47377),
            .I(n20671));
    InMux I__10458 (
            .O(N__47374),
            .I(N__47368));
    InMux I__10457 (
            .O(N__47373),
            .I(N__47368));
    LocalMux I__10456 (
            .O(N__47368),
            .I(N__47364));
    InMux I__10455 (
            .O(N__47367),
            .I(N__47360));
    Span4Mux_v I__10454 (
            .O(N__47364),
            .I(N__47357));
    InMux I__10453 (
            .O(N__47363),
            .I(N__47353));
    LocalMux I__10452 (
            .O(N__47360),
            .I(N__47349));
    Span4Mux_v I__10451 (
            .O(N__47357),
            .I(N__47346));
    InMux I__10450 (
            .O(N__47356),
            .I(N__47343));
    LocalMux I__10449 (
            .O(N__47353),
            .I(N__47340));
    InMux I__10448 (
            .O(N__47352),
            .I(N__47337));
    Span4Mux_h I__10447 (
            .O(N__47349),
            .I(N__47334));
    Sp12to4 I__10446 (
            .O(N__47346),
            .I(N__47329));
    LocalMux I__10445 (
            .O(N__47343),
            .I(N__47329));
    Span4Mux_h I__10444 (
            .O(N__47340),
            .I(N__47324));
    LocalMux I__10443 (
            .O(N__47337),
            .I(N__47324));
    Odrv4 I__10442 (
            .O(N__47334),
            .I(n14_adj_1653));
    Odrv12 I__10441 (
            .O(N__47329),
            .I(n14_adj_1653));
    Odrv4 I__10440 (
            .O(N__47324),
            .I(n14_adj_1653));
    InMux I__10439 (
            .O(N__47317),
            .I(n20672));
    InMux I__10438 (
            .O(N__47314),
            .I(n20673));
    InMux I__10437 (
            .O(N__47311),
            .I(n20674));
    InMux I__10436 (
            .O(N__47308),
            .I(N__47305));
    LocalMux I__10435 (
            .O(N__47305),
            .I(N__47302));
    Span4Mux_v I__10434 (
            .O(N__47302),
            .I(N__47299));
    Odrv4 I__10433 (
            .O(N__47299),
            .I(n14_adj_1607));
    InMux I__10432 (
            .O(N__47296),
            .I(n20675));
    InMux I__10431 (
            .O(N__47293),
            .I(N__47290));
    LocalMux I__10430 (
            .O(N__47290),
            .I(N__47286));
    CascadeMux I__10429 (
            .O(N__47289),
            .I(N__47283));
    Span4Mux_h I__10428 (
            .O(N__47286),
            .I(N__47280));
    InMux I__10427 (
            .O(N__47283),
            .I(N__47277));
    Span4Mux_h I__10426 (
            .O(N__47280),
            .I(N__47274));
    LocalMux I__10425 (
            .O(N__47277),
            .I(data_idxvec_15));
    Odrv4 I__10424 (
            .O(N__47274),
            .I(data_idxvec_15));
    InMux I__10423 (
            .O(N__47269),
            .I(N__47264));
    InMux I__10422 (
            .O(N__47268),
            .I(N__47261));
    CascadeMux I__10421 (
            .O(N__47267),
            .I(N__47258));
    LocalMux I__10420 (
            .O(N__47264),
            .I(N__47255));
    LocalMux I__10419 (
            .O(N__47261),
            .I(N__47252));
    InMux I__10418 (
            .O(N__47258),
            .I(N__47249));
    Span4Mux_h I__10417 (
            .O(N__47255),
            .I(N__47246));
    Span4Mux_h I__10416 (
            .O(N__47252),
            .I(N__47243));
    LocalMux I__10415 (
            .O(N__47249),
            .I(N__47236));
    Span4Mux_h I__10414 (
            .O(N__47246),
            .I(N__47236));
    Span4Mux_h I__10413 (
            .O(N__47243),
            .I(N__47236));
    Odrv4 I__10412 (
            .O(N__47236),
            .I(buf_dds0_4));
    InMux I__10411 (
            .O(N__47233),
            .I(N__47229));
    InMux I__10410 (
            .O(N__47232),
            .I(N__47226));
    LocalMux I__10409 (
            .O(N__47229),
            .I(N__47223));
    LocalMux I__10408 (
            .O(N__47226),
            .I(N__47220));
    Span4Mux_v I__10407 (
            .O(N__47223),
            .I(N__47214));
    Span4Mux_h I__10406 (
            .O(N__47220),
            .I(N__47214));
    InMux I__10405 (
            .O(N__47219),
            .I(N__47211));
    Span4Mux_h I__10404 (
            .O(N__47214),
            .I(N__47208));
    LocalMux I__10403 (
            .O(N__47211),
            .I(buf_dds0_0));
    Odrv4 I__10402 (
            .O(N__47208),
            .I(buf_dds0_0));
    InMux I__10401 (
            .O(N__47203),
            .I(N__47199));
    InMux I__10400 (
            .O(N__47202),
            .I(N__47196));
    LocalMux I__10399 (
            .O(N__47199),
            .I(N__47193));
    LocalMux I__10398 (
            .O(N__47196),
            .I(data_idxvec_0));
    Odrv4 I__10397 (
            .O(N__47193),
            .I(data_idxvec_0));
    InMux I__10396 (
            .O(N__47188),
            .I(bfn_16_16_0_));
    InMux I__10395 (
            .O(N__47185),
            .I(N__47182));
    LocalMux I__10394 (
            .O(N__47182),
            .I(N__47179));
    Span4Mux_v I__10393 (
            .O(N__47179),
            .I(N__47176));
    Span4Mux_v I__10392 (
            .O(N__47176),
            .I(N__47172));
    InMux I__10391 (
            .O(N__47175),
            .I(N__47169));
    Sp12to4 I__10390 (
            .O(N__47172),
            .I(N__47164));
    LocalMux I__10389 (
            .O(N__47169),
            .I(N__47164));
    Odrv12 I__10388 (
            .O(N__47164),
            .I(n14_adj_1613));
    InMux I__10387 (
            .O(N__47161),
            .I(n20661));
    InMux I__10386 (
            .O(N__47158),
            .I(N__47155));
    LocalMux I__10385 (
            .O(N__47155),
            .I(N__47151));
    InMux I__10384 (
            .O(N__47154),
            .I(N__47148));
    Span4Mux_v I__10383 (
            .O(N__47151),
            .I(N__47145));
    LocalMux I__10382 (
            .O(N__47148),
            .I(n14_adj_1612));
    Odrv4 I__10381 (
            .O(N__47145),
            .I(n14_adj_1612));
    InMux I__10380 (
            .O(N__47140),
            .I(n20662));
    CascadeMux I__10379 (
            .O(N__47137),
            .I(N__47134));
    InMux I__10378 (
            .O(N__47134),
            .I(N__47130));
    InMux I__10377 (
            .O(N__47133),
            .I(N__47127));
    LocalMux I__10376 (
            .O(N__47130),
            .I(N__47124));
    LocalMux I__10375 (
            .O(N__47127),
            .I(data_idxvec_3));
    Odrv4 I__10374 (
            .O(N__47124),
            .I(data_idxvec_3));
    InMux I__10373 (
            .O(N__47119),
            .I(n20663));
    InMux I__10372 (
            .O(N__47116),
            .I(n20664));
    CascadeMux I__10371 (
            .O(N__47113),
            .I(N__47109));
    InMux I__10370 (
            .O(N__47112),
            .I(N__47106));
    InMux I__10369 (
            .O(N__47109),
            .I(N__47103));
    LocalMux I__10368 (
            .O(N__47106),
            .I(N__47100));
    LocalMux I__10367 (
            .O(N__47103),
            .I(N__47094));
    Span4Mux_h I__10366 (
            .O(N__47100),
            .I(N__47094));
    InMux I__10365 (
            .O(N__47099),
            .I(N__47091));
    Span4Mux_h I__10364 (
            .O(N__47094),
            .I(N__47088));
    LocalMux I__10363 (
            .O(N__47091),
            .I(N__47085));
    Odrv4 I__10362 (
            .O(N__47088),
            .I(n14_adj_1661));
    Odrv12 I__10361 (
            .O(N__47085),
            .I(n14_adj_1661));
    InMux I__10360 (
            .O(N__47080),
            .I(n20665));
    InMux I__10359 (
            .O(N__47077),
            .I(N__47073));
    CascadeMux I__10358 (
            .O(N__47076),
            .I(N__47070));
    LocalMux I__10357 (
            .O(N__47073),
            .I(N__47066));
    InMux I__10356 (
            .O(N__47070),
            .I(N__47063));
    InMux I__10355 (
            .O(N__47069),
            .I(N__47060));
    Span4Mux_v I__10354 (
            .O(N__47066),
            .I(N__47057));
    LocalMux I__10353 (
            .O(N__47063),
            .I(N__47052));
    LocalMux I__10352 (
            .O(N__47060),
            .I(N__47052));
    Span4Mux_h I__10351 (
            .O(N__47057),
            .I(N__47047));
    Span4Mux_v I__10350 (
            .O(N__47052),
            .I(N__47047));
    Odrv4 I__10349 (
            .O(N__47047),
            .I(n14_adj_1610));
    InMux I__10348 (
            .O(N__47044),
            .I(n20666));
    CascadeMux I__10347 (
            .O(N__47041),
            .I(n26_adj_1580_cascade_));
    InMux I__10346 (
            .O(N__47038),
            .I(N__47035));
    LocalMux I__10345 (
            .O(N__47035),
            .I(N__47032));
    Span4Mux_h I__10344 (
            .O(N__47032),
            .I(N__47027));
    InMux I__10343 (
            .O(N__47031),
            .I(N__47022));
    InMux I__10342 (
            .O(N__47030),
            .I(N__47022));
    Odrv4 I__10341 (
            .O(N__47027),
            .I(acadc_skipCount_0));
    LocalMux I__10340 (
            .O(N__47022),
            .I(acadc_skipCount_0));
    CascadeMux I__10339 (
            .O(N__47017),
            .I(n23552_cascade_));
    InMux I__10338 (
            .O(N__47014),
            .I(N__47010));
    CascadeMux I__10337 (
            .O(N__47013),
            .I(N__47006));
    LocalMux I__10336 (
            .O(N__47010),
            .I(N__47003));
    InMux I__10335 (
            .O(N__47009),
            .I(N__47000));
    InMux I__10334 (
            .O(N__47006),
            .I(N__46997));
    Odrv4 I__10333 (
            .O(N__47003),
            .I(req_data_cnt_0));
    LocalMux I__10332 (
            .O(N__47000),
            .I(req_data_cnt_0));
    LocalMux I__10331 (
            .O(N__46997),
            .I(req_data_cnt_0));
    InMux I__10330 (
            .O(N__46990),
            .I(N__46987));
    LocalMux I__10329 (
            .O(N__46987),
            .I(N__46984));
    Span4Mux_h I__10328 (
            .O(N__46984),
            .I(N__46981));
    Span4Mux_h I__10327 (
            .O(N__46981),
            .I(N__46978));
    Odrv4 I__10326 (
            .O(N__46978),
            .I(n16));
    InMux I__10325 (
            .O(N__46975),
            .I(N__46972));
    LocalMux I__10324 (
            .O(N__46972),
            .I(N__46969));
    Span4Mux_v I__10323 (
            .O(N__46969),
            .I(N__46966));
    Sp12to4 I__10322 (
            .O(N__46966),
            .I(N__46963));
    Odrv12 I__10321 (
            .O(N__46963),
            .I(n23300));
    CascadeMux I__10320 (
            .O(N__46960),
            .I(N__46957));
    InMux I__10319 (
            .O(N__46957),
            .I(N__46953));
    InMux I__10318 (
            .O(N__46956),
            .I(N__46950));
    LocalMux I__10317 (
            .O(N__46953),
            .I(N__46947));
    LocalMux I__10316 (
            .O(N__46950),
            .I(N__46943));
    Span4Mux_h I__10315 (
            .O(N__46947),
            .I(N__46940));
    InMux I__10314 (
            .O(N__46946),
            .I(N__46937));
    Span12Mux_s9_v I__10313 (
            .O(N__46943),
            .I(N__46934));
    Span4Mux_h I__10312 (
            .O(N__46940),
            .I(N__46931));
    LocalMux I__10311 (
            .O(N__46937),
            .I(buf_adcdata_iac_8));
    Odrv12 I__10310 (
            .O(N__46934),
            .I(buf_adcdata_iac_8));
    Odrv4 I__10309 (
            .O(N__46931),
            .I(buf_adcdata_iac_8));
    InMux I__10308 (
            .O(N__46924),
            .I(N__46921));
    LocalMux I__10307 (
            .O(N__46921),
            .I(N__46917));
    InMux I__10306 (
            .O(N__46920),
            .I(N__46914));
    Span4Mux_h I__10305 (
            .O(N__46917),
            .I(N__46911));
    LocalMux I__10304 (
            .O(N__46914),
            .I(N__46907));
    Span4Mux_v I__10303 (
            .O(N__46911),
            .I(N__46904));
    CascadeMux I__10302 (
            .O(N__46910),
            .I(N__46901));
    Span4Mux_h I__10301 (
            .O(N__46907),
            .I(N__46898));
    Span4Mux_h I__10300 (
            .O(N__46904),
            .I(N__46895));
    InMux I__10299 (
            .O(N__46901),
            .I(N__46892));
    Span4Mux_h I__10298 (
            .O(N__46898),
            .I(N__46889));
    Span4Mux_h I__10297 (
            .O(N__46895),
            .I(N__46886));
    LocalMux I__10296 (
            .O(N__46892),
            .I(buf_adcdata_iac_15));
    Odrv4 I__10295 (
            .O(N__46889),
            .I(buf_adcdata_iac_15));
    Odrv4 I__10294 (
            .O(N__46886),
            .I(buf_adcdata_iac_15));
    InMux I__10293 (
            .O(N__46879),
            .I(N__46876));
    LocalMux I__10292 (
            .O(N__46876),
            .I(N__46873));
    Span4Mux_h I__10291 (
            .O(N__46873),
            .I(N__46870));
    Span4Mux_h I__10290 (
            .O(N__46870),
            .I(N__46867));
    Odrv4 I__10289 (
            .O(N__46867),
            .I(n16_adj_1713));
    InMux I__10288 (
            .O(N__46864),
            .I(N__46861));
    LocalMux I__10287 (
            .O(N__46861),
            .I(N__46858));
    Span4Mux_v I__10286 (
            .O(N__46858),
            .I(N__46855));
    Odrv4 I__10285 (
            .O(N__46855),
            .I(n22268));
    InMux I__10284 (
            .O(N__46852),
            .I(N__46839));
    InMux I__10283 (
            .O(N__46851),
            .I(N__46836));
    InMux I__10282 (
            .O(N__46850),
            .I(N__46831));
    InMux I__10281 (
            .O(N__46849),
            .I(N__46831));
    InMux I__10280 (
            .O(N__46848),
            .I(N__46826));
    InMux I__10279 (
            .O(N__46847),
            .I(N__46826));
    InMux I__10278 (
            .O(N__46846),
            .I(N__46821));
    InMux I__10277 (
            .O(N__46845),
            .I(N__46821));
    CascadeMux I__10276 (
            .O(N__46844),
            .I(N__46814));
    CascadeMux I__10275 (
            .O(N__46843),
            .I(N__46811));
    InMux I__10274 (
            .O(N__46842),
            .I(N__46807));
    LocalMux I__10273 (
            .O(N__46839),
            .I(N__46804));
    LocalMux I__10272 (
            .O(N__46836),
            .I(N__46799));
    LocalMux I__10271 (
            .O(N__46831),
            .I(N__46799));
    LocalMux I__10270 (
            .O(N__46826),
            .I(N__46794));
    LocalMux I__10269 (
            .O(N__46821),
            .I(N__46794));
    InMux I__10268 (
            .O(N__46820),
            .I(N__46791));
    InMux I__10267 (
            .O(N__46819),
            .I(N__46788));
    InMux I__10266 (
            .O(N__46818),
            .I(N__46785));
    InMux I__10265 (
            .O(N__46817),
            .I(N__46782));
    InMux I__10264 (
            .O(N__46814),
            .I(N__46775));
    InMux I__10263 (
            .O(N__46811),
            .I(N__46775));
    InMux I__10262 (
            .O(N__46810),
            .I(N__46775));
    LocalMux I__10261 (
            .O(N__46807),
            .I(N__46768));
    Span4Mux_v I__10260 (
            .O(N__46804),
            .I(N__46768));
    Span4Mux_v I__10259 (
            .O(N__46799),
            .I(N__46768));
    Span4Mux_h I__10258 (
            .O(N__46794),
            .I(N__46765));
    LocalMux I__10257 (
            .O(N__46791),
            .I(n13141));
    LocalMux I__10256 (
            .O(N__46788),
            .I(n13141));
    LocalMux I__10255 (
            .O(N__46785),
            .I(n13141));
    LocalMux I__10254 (
            .O(N__46782),
            .I(n13141));
    LocalMux I__10253 (
            .O(N__46775),
            .I(n13141));
    Odrv4 I__10252 (
            .O(N__46768),
            .I(n13141));
    Odrv4 I__10251 (
            .O(N__46765),
            .I(n13141));
    InMux I__10250 (
            .O(N__46750),
            .I(N__46745));
    InMux I__10249 (
            .O(N__46749),
            .I(N__46742));
    InMux I__10248 (
            .O(N__46748),
            .I(N__46739));
    LocalMux I__10247 (
            .O(N__46745),
            .I(N__46733));
    LocalMux I__10246 (
            .O(N__46742),
            .I(N__46730));
    LocalMux I__10245 (
            .O(N__46739),
            .I(N__46727));
    InMux I__10244 (
            .O(N__46738),
            .I(N__46720));
    InMux I__10243 (
            .O(N__46737),
            .I(N__46720));
    InMux I__10242 (
            .O(N__46736),
            .I(N__46720));
    Span4Mux_v I__10241 (
            .O(N__46733),
            .I(N__46717));
    Span4Mux_v I__10240 (
            .O(N__46730),
            .I(N__46712));
    Span4Mux_v I__10239 (
            .O(N__46727),
            .I(N__46712));
    LocalMux I__10238 (
            .O(N__46720),
            .I(N__46709));
    Span4Mux_v I__10237 (
            .O(N__46717),
            .I(N__46706));
    Span4Mux_h I__10236 (
            .O(N__46712),
            .I(N__46701));
    Span4Mux_v I__10235 (
            .O(N__46709),
            .I(N__46701));
    Span4Mux_v I__10234 (
            .O(N__46706),
            .I(N__46698));
    Sp12to4 I__10233 (
            .O(N__46701),
            .I(N__46695));
    Odrv4 I__10232 (
            .O(N__46698),
            .I(n12610));
    Odrv12 I__10231 (
            .O(N__46695),
            .I(n12610));
    CascadeMux I__10230 (
            .O(N__46690),
            .I(n12021_cascade_));
    CEMux I__10229 (
            .O(N__46687),
            .I(N__46684));
    LocalMux I__10228 (
            .O(N__46684),
            .I(n12614));
    CascadeMux I__10227 (
            .O(N__46681),
            .I(n25_cascade_));
    CEMux I__10226 (
            .O(N__46678),
            .I(N__46675));
    LocalMux I__10225 (
            .O(N__46675),
            .I(N__46672));
    Span4Mux_v I__10224 (
            .O(N__46672),
            .I(N__46669));
    Sp12to4 I__10223 (
            .O(N__46669),
            .I(N__46666));
    Odrv12 I__10222 (
            .O(N__46666),
            .I(n12548));
    CascadeMux I__10221 (
            .O(N__46663),
            .I(N__46659));
    CascadeMux I__10220 (
            .O(N__46662),
            .I(N__46655));
    InMux I__10219 (
            .O(N__46659),
            .I(N__46651));
    CascadeMux I__10218 (
            .O(N__46658),
            .I(N__46648));
    InMux I__10217 (
            .O(N__46655),
            .I(N__46643));
    CascadeMux I__10216 (
            .O(N__46654),
            .I(N__46639));
    LocalMux I__10215 (
            .O(N__46651),
            .I(N__46636));
    InMux I__10214 (
            .O(N__46648),
            .I(N__46633));
    InMux I__10213 (
            .O(N__46647),
            .I(N__46630));
    InMux I__10212 (
            .O(N__46646),
            .I(N__46626));
    LocalMux I__10211 (
            .O(N__46643),
            .I(N__46623));
    InMux I__10210 (
            .O(N__46642),
            .I(N__46617));
    InMux I__10209 (
            .O(N__46639),
            .I(N__46614));
    Span4Mux_v I__10208 (
            .O(N__46636),
            .I(N__46611));
    LocalMux I__10207 (
            .O(N__46633),
            .I(N__46608));
    LocalMux I__10206 (
            .O(N__46630),
            .I(N__46605));
    CascadeMux I__10205 (
            .O(N__46629),
            .I(N__46602));
    LocalMux I__10204 (
            .O(N__46626),
            .I(N__46599));
    Span4Mux_v I__10203 (
            .O(N__46623),
            .I(N__46596));
    InMux I__10202 (
            .O(N__46622),
            .I(N__46593));
    InMux I__10201 (
            .O(N__46621),
            .I(N__46588));
    InMux I__10200 (
            .O(N__46620),
            .I(N__46588));
    LocalMux I__10199 (
            .O(N__46617),
            .I(N__46585));
    LocalMux I__10198 (
            .O(N__46614),
            .I(N__46582));
    Span4Mux_h I__10197 (
            .O(N__46611),
            .I(N__46575));
    Span4Mux_h I__10196 (
            .O(N__46608),
            .I(N__46575));
    Span4Mux_v I__10195 (
            .O(N__46605),
            .I(N__46575));
    InMux I__10194 (
            .O(N__46602),
            .I(N__46572));
    Span4Mux_v I__10193 (
            .O(N__46599),
            .I(N__46569));
    Span4Mux_h I__10192 (
            .O(N__46596),
            .I(N__46564));
    LocalMux I__10191 (
            .O(N__46593),
            .I(N__46564));
    LocalMux I__10190 (
            .O(N__46588),
            .I(N__46561));
    Span4Mux_h I__10189 (
            .O(N__46585),
            .I(N__46558));
    Span12Mux_v I__10188 (
            .O(N__46582),
            .I(N__46555));
    Span4Mux_v I__10187 (
            .O(N__46575),
            .I(N__46552));
    LocalMux I__10186 (
            .O(N__46572),
            .I(N__46541));
    Span4Mux_v I__10185 (
            .O(N__46569),
            .I(N__46541));
    Span4Mux_h I__10184 (
            .O(N__46564),
            .I(N__46541));
    Span4Mux_h I__10183 (
            .O(N__46561),
            .I(N__46541));
    Span4Mux_h I__10182 (
            .O(N__46558),
            .I(N__46541));
    Odrv12 I__10181 (
            .O(N__46555),
            .I(comm_buf_0_7));
    Odrv4 I__10180 (
            .O(N__46552),
            .I(comm_buf_0_7));
    Odrv4 I__10179 (
            .O(N__46541),
            .I(comm_buf_0_7));
    CascadeMux I__10178 (
            .O(N__46534),
            .I(N__46531));
    InMux I__10177 (
            .O(N__46531),
            .I(N__46527));
    InMux I__10176 (
            .O(N__46530),
            .I(N__46524));
    LocalMux I__10175 (
            .O(N__46527),
            .I(N__46521));
    LocalMux I__10174 (
            .O(N__46524),
            .I(N__46517));
    Span4Mux_h I__10173 (
            .O(N__46521),
            .I(N__46514));
    InMux I__10172 (
            .O(N__46520),
            .I(N__46511));
    Odrv4 I__10171 (
            .O(N__46517),
            .I(n21964));
    Odrv4 I__10170 (
            .O(N__46514),
            .I(n21964));
    LocalMux I__10169 (
            .O(N__46511),
            .I(n21964));
    CascadeMux I__10168 (
            .O(N__46504),
            .I(N__46501));
    InMux I__10167 (
            .O(N__46501),
            .I(N__46498));
    LocalMux I__10166 (
            .O(N__46498),
            .I(N__46495));
    Span4Mux_v I__10165 (
            .O(N__46495),
            .I(N__46492));
    Span4Mux_v I__10164 (
            .O(N__46492),
            .I(N__46489));
    Odrv4 I__10163 (
            .O(N__46489),
            .I(n11379));
    InMux I__10162 (
            .O(N__46486),
            .I(N__46483));
    LocalMux I__10161 (
            .O(N__46483),
            .I(N__46478));
    InMux I__10160 (
            .O(N__46482),
            .I(N__46475));
    InMux I__10159 (
            .O(N__46481),
            .I(N__46471));
    Span4Mux_v I__10158 (
            .O(N__46478),
            .I(N__46468));
    LocalMux I__10157 (
            .O(N__46475),
            .I(N__46465));
    InMux I__10156 (
            .O(N__46474),
            .I(N__46462));
    LocalMux I__10155 (
            .O(N__46471),
            .I(n9));
    Odrv4 I__10154 (
            .O(N__46468),
            .I(n9));
    Odrv4 I__10153 (
            .O(N__46465),
            .I(n9));
    LocalMux I__10152 (
            .O(N__46462),
            .I(n9));
    InMux I__10151 (
            .O(N__46453),
            .I(N__46450));
    LocalMux I__10150 (
            .O(N__46450),
            .I(n22059));
    CascadeMux I__10149 (
            .O(N__46447),
            .I(N__46444));
    InMux I__10148 (
            .O(N__46444),
            .I(N__46441));
    LocalMux I__10147 (
            .O(N__46441),
            .I(N__46438));
    Odrv4 I__10146 (
            .O(N__46438),
            .I(n26_adj_1740));
    CascadeMux I__10145 (
            .O(N__46435),
            .I(n18850_cascade_));
    CEMux I__10144 (
            .O(N__46432),
            .I(N__46428));
    CEMux I__10143 (
            .O(N__46431),
            .I(N__46423));
    LocalMux I__10142 (
            .O(N__46428),
            .I(N__46420));
    CEMux I__10141 (
            .O(N__46427),
            .I(N__46416));
    CEMux I__10140 (
            .O(N__46426),
            .I(N__46413));
    LocalMux I__10139 (
            .O(N__46423),
            .I(N__46408));
    Span4Mux_h I__10138 (
            .O(N__46420),
            .I(N__46408));
    CEMux I__10137 (
            .O(N__46419),
            .I(N__46405));
    LocalMux I__10136 (
            .O(N__46416),
            .I(N__46399));
    LocalMux I__10135 (
            .O(N__46413),
            .I(N__46396));
    Span4Mux_v I__10134 (
            .O(N__46408),
            .I(N__46391));
    LocalMux I__10133 (
            .O(N__46405),
            .I(N__46391));
    CEMux I__10132 (
            .O(N__46404),
            .I(N__46387));
    CEMux I__10131 (
            .O(N__46403),
            .I(N__46384));
    CEMux I__10130 (
            .O(N__46402),
            .I(N__46381));
    Span4Mux_v I__10129 (
            .O(N__46399),
            .I(N__46378));
    Span12Mux_h I__10128 (
            .O(N__46396),
            .I(N__46375));
    Span4Mux_h I__10127 (
            .O(N__46391),
            .I(N__46372));
    InMux I__10126 (
            .O(N__46390),
            .I(N__46369));
    LocalMux I__10125 (
            .O(N__46387),
            .I(n13076));
    LocalMux I__10124 (
            .O(N__46384),
            .I(n13076));
    LocalMux I__10123 (
            .O(N__46381),
            .I(n13076));
    Odrv4 I__10122 (
            .O(N__46378),
            .I(n13076));
    Odrv12 I__10121 (
            .O(N__46375),
            .I(n13076));
    Odrv4 I__10120 (
            .O(N__46372),
            .I(n13076));
    LocalMux I__10119 (
            .O(N__46369),
            .I(n13076));
    SRMux I__10118 (
            .O(N__46354),
            .I(N__46345));
    SRMux I__10117 (
            .O(N__46353),
            .I(N__46342));
    SRMux I__10116 (
            .O(N__46352),
            .I(N__46338));
    SRMux I__10115 (
            .O(N__46351),
            .I(N__46335));
    SRMux I__10114 (
            .O(N__46350),
            .I(N__46332));
    SRMux I__10113 (
            .O(N__46349),
            .I(N__46329));
    SRMux I__10112 (
            .O(N__46348),
            .I(N__46326));
    LocalMux I__10111 (
            .O(N__46345),
            .I(N__46323));
    LocalMux I__10110 (
            .O(N__46342),
            .I(N__46320));
    SRMux I__10109 (
            .O(N__46341),
            .I(N__46317));
    LocalMux I__10108 (
            .O(N__46338),
            .I(N__46314));
    LocalMux I__10107 (
            .O(N__46335),
            .I(N__46311));
    LocalMux I__10106 (
            .O(N__46332),
            .I(N__46306));
    LocalMux I__10105 (
            .O(N__46329),
            .I(N__46306));
    LocalMux I__10104 (
            .O(N__46326),
            .I(N__46303));
    Span4Mux_h I__10103 (
            .O(N__46323),
            .I(N__46300));
    Span4Mux_v I__10102 (
            .O(N__46320),
            .I(N__46297));
    LocalMux I__10101 (
            .O(N__46317),
            .I(N__46290));
    Span4Mux_h I__10100 (
            .O(N__46314),
            .I(N__46290));
    Span4Mux_h I__10099 (
            .O(N__46311),
            .I(N__46290));
    Span4Mux_h I__10098 (
            .O(N__46306),
            .I(N__46285));
    Span4Mux_h I__10097 (
            .O(N__46303),
            .I(N__46285));
    Odrv4 I__10096 (
            .O(N__46300),
            .I(n15531));
    Odrv4 I__10095 (
            .O(N__46297),
            .I(n15531));
    Odrv4 I__10094 (
            .O(N__46290),
            .I(n15531));
    Odrv4 I__10093 (
            .O(N__46285),
            .I(n15531));
    InMux I__10092 (
            .O(N__46276),
            .I(N__46273));
    LocalMux I__10091 (
            .O(N__46273),
            .I(N__46270));
    Span4Mux_v I__10090 (
            .O(N__46270),
            .I(N__46267));
    Span4Mux_v I__10089 (
            .O(N__46267),
            .I(N__46264));
    Sp12to4 I__10088 (
            .O(N__46264),
            .I(N__46261));
    Odrv12 I__10087 (
            .O(N__46261),
            .I(comm_buf_3_3));
    InMux I__10086 (
            .O(N__46258),
            .I(N__46254));
    InMux I__10085 (
            .O(N__46257),
            .I(N__46251));
    LocalMux I__10084 (
            .O(N__46254),
            .I(N__46248));
    LocalMux I__10083 (
            .O(N__46251),
            .I(N__46245));
    Span4Mux_v I__10082 (
            .O(N__46248),
            .I(N__46242));
    Odrv4 I__10081 (
            .O(N__46245),
            .I(comm_buf_6_3));
    Odrv4 I__10080 (
            .O(N__46242),
            .I(comm_buf_6_3));
    InMux I__10079 (
            .O(N__46237),
            .I(N__46234));
    LocalMux I__10078 (
            .O(N__46234),
            .I(N__46231));
    Odrv4 I__10077 (
            .O(N__46231),
            .I(n18851));
    InMux I__10076 (
            .O(N__46228),
            .I(N__46225));
    LocalMux I__10075 (
            .O(N__46225),
            .I(N__46222));
    Odrv4 I__10074 (
            .O(N__46222),
            .I(comm_buf_5_3));
    InMux I__10073 (
            .O(N__46219),
            .I(N__46216));
    LocalMux I__10072 (
            .O(N__46216),
            .I(n22346));
    CascadeMux I__10071 (
            .O(N__46213),
            .I(n18853_cascade_));
    InMux I__10070 (
            .O(N__46210),
            .I(N__46207));
    LocalMux I__10069 (
            .O(N__46207),
            .I(n23378));
    InMux I__10068 (
            .O(N__46204),
            .I(N__46196));
    InMux I__10067 (
            .O(N__46203),
            .I(N__46192));
    InMux I__10066 (
            .O(N__46202),
            .I(N__46189));
    InMux I__10065 (
            .O(N__46201),
            .I(N__46186));
    InMux I__10064 (
            .O(N__46200),
            .I(N__46183));
    InMux I__10063 (
            .O(N__46199),
            .I(N__46180));
    LocalMux I__10062 (
            .O(N__46196),
            .I(N__46177));
    InMux I__10061 (
            .O(N__46195),
            .I(N__46174));
    LocalMux I__10060 (
            .O(N__46192),
            .I(N__46171));
    LocalMux I__10059 (
            .O(N__46189),
            .I(N__46168));
    LocalMux I__10058 (
            .O(N__46186),
            .I(N__46165));
    LocalMux I__10057 (
            .O(N__46183),
            .I(N__46160));
    LocalMux I__10056 (
            .O(N__46180),
            .I(N__46157));
    Span4Mux_h I__10055 (
            .O(N__46177),
            .I(N__46150));
    LocalMux I__10054 (
            .O(N__46174),
            .I(N__46150));
    Span4Mux_h I__10053 (
            .O(N__46171),
            .I(N__46150));
    Span4Mux_h I__10052 (
            .O(N__46168),
            .I(N__46145));
    Span4Mux_h I__10051 (
            .O(N__46165),
            .I(N__46145));
    InMux I__10050 (
            .O(N__46164),
            .I(N__46142));
    InMux I__10049 (
            .O(N__46163),
            .I(N__46139));
    Span4Mux_v I__10048 (
            .O(N__46160),
            .I(N__46132));
    Span4Mux_v I__10047 (
            .O(N__46157),
            .I(N__46132));
    Span4Mux_v I__10046 (
            .O(N__46150),
            .I(N__46132));
    Odrv4 I__10045 (
            .O(N__46145),
            .I(n6776));
    LocalMux I__10044 (
            .O(N__46142),
            .I(n6776));
    LocalMux I__10043 (
            .O(N__46139),
            .I(n6776));
    Odrv4 I__10042 (
            .O(N__46132),
            .I(n6776));
    CascadeMux I__10041 (
            .O(N__46123),
            .I(N__46120));
    InMux I__10040 (
            .O(N__46120),
            .I(N__46117));
    LocalMux I__10039 (
            .O(N__46117),
            .I(N__46113));
    CascadeMux I__10038 (
            .O(N__46116),
            .I(N__46110));
    Span4Mux_v I__10037 (
            .O(N__46113),
            .I(N__46106));
    InMux I__10036 (
            .O(N__46110),
            .I(N__46101));
    InMux I__10035 (
            .O(N__46109),
            .I(N__46101));
    Sp12to4 I__10034 (
            .O(N__46106),
            .I(N__46096));
    LocalMux I__10033 (
            .O(N__46101),
            .I(N__46096));
    Odrv12 I__10032 (
            .O(N__46096),
            .I(comm_buf_2_3));
    InMux I__10031 (
            .O(N__46093),
            .I(N__46090));
    LocalMux I__10030 (
            .O(N__46090),
            .I(N__46087));
    Span4Mux_h I__10029 (
            .O(N__46087),
            .I(N__46084));
    Span4Mux_h I__10028 (
            .O(N__46084),
            .I(N__46081));
    Odrv4 I__10027 (
            .O(N__46081),
            .I(n18858));
    InMux I__10026 (
            .O(N__46078),
            .I(N__46075));
    LocalMux I__10025 (
            .O(N__46075),
            .I(N__46072));
    Span4Mux_v I__10024 (
            .O(N__46072),
            .I(N__46068));
    InMux I__10023 (
            .O(N__46071),
            .I(N__46065));
    Span4Mux_h I__10022 (
            .O(N__46068),
            .I(N__46062));
    LocalMux I__10021 (
            .O(N__46065),
            .I(N__46059));
    Span4Mux_v I__10020 (
            .O(N__46062),
            .I(N__46053));
    Span4Mux_h I__10019 (
            .O(N__46059),
            .I(N__46053));
    InMux I__10018 (
            .O(N__46058),
            .I(N__46050));
    Odrv4 I__10017 (
            .O(N__46053),
            .I(comm_tx_buf_3));
    LocalMux I__10016 (
            .O(N__46050),
            .I(comm_tx_buf_3));
    InMux I__10015 (
            .O(N__46045),
            .I(N__46042));
    LocalMux I__10014 (
            .O(N__46042),
            .I(N__46039));
    Span4Mux_h I__10013 (
            .O(N__46039),
            .I(N__46036));
    Sp12to4 I__10012 (
            .O(N__46036),
            .I(N__46033));
    Span12Mux_v I__10011 (
            .O(N__46033),
            .I(N__46030));
    Span12Mux_h I__10010 (
            .O(N__46030),
            .I(N__46027));
    Odrv12 I__10009 (
            .O(N__46027),
            .I(THERMOSTAT));
    InMux I__10008 (
            .O(N__46024),
            .I(N__46021));
    LocalMux I__10007 (
            .O(N__46021),
            .I(N__46018));
    Span4Mux_h I__10006 (
            .O(N__46018),
            .I(N__46015));
    Odrv4 I__10005 (
            .O(N__46015),
            .I(buf_control_7));
    CascadeMux I__10004 (
            .O(N__46012),
            .I(N__46009));
    InMux I__10003 (
            .O(N__46009),
            .I(N__46002));
    InMux I__10002 (
            .O(N__46008),
            .I(N__46002));
    InMux I__10001 (
            .O(N__46007),
            .I(N__45999));
    LocalMux I__10000 (
            .O(N__46002),
            .I(N__45992));
    LocalMux I__9999 (
            .O(N__45999),
            .I(N__45989));
    InMux I__9998 (
            .O(N__45998),
            .I(N__45986));
    InMux I__9997 (
            .O(N__45997),
            .I(N__45981));
    InMux I__9996 (
            .O(N__45996),
            .I(N__45981));
    InMux I__9995 (
            .O(N__45995),
            .I(N__45978));
    Span4Mux_v I__9994 (
            .O(N__45992),
            .I(N__45968));
    Span4Mux_h I__9993 (
            .O(N__45989),
            .I(N__45968));
    LocalMux I__9992 (
            .O(N__45986),
            .I(N__45968));
    LocalMux I__9991 (
            .O(N__45981),
            .I(N__45968));
    LocalMux I__9990 (
            .O(N__45978),
            .I(N__45965));
    InMux I__9989 (
            .O(N__45977),
            .I(N__45962));
    Odrv4 I__9988 (
            .O(N__45968),
            .I(n12585));
    Odrv12 I__9987 (
            .O(N__45965),
            .I(n12585));
    LocalMux I__9986 (
            .O(N__45962),
            .I(n12585));
    CascadeMux I__9985 (
            .O(N__45955),
            .I(N__45950));
    CascadeMux I__9984 (
            .O(N__45954),
            .I(N__45946));
    CascadeMux I__9983 (
            .O(N__45953),
            .I(N__45943));
    InMux I__9982 (
            .O(N__45950),
            .I(N__45937));
    InMux I__9981 (
            .O(N__45949),
            .I(N__45934));
    InMux I__9980 (
            .O(N__45946),
            .I(N__45930));
    InMux I__9979 (
            .O(N__45943),
            .I(N__45925));
    InMux I__9978 (
            .O(N__45942),
            .I(N__45925));
    InMux I__9977 (
            .O(N__45941),
            .I(N__45920));
    InMux I__9976 (
            .O(N__45940),
            .I(N__45920));
    LocalMux I__9975 (
            .O(N__45937),
            .I(N__45917));
    LocalMux I__9974 (
            .O(N__45934),
            .I(N__45914));
    InMux I__9973 (
            .O(N__45933),
            .I(N__45911));
    LocalMux I__9972 (
            .O(N__45930),
            .I(N__45904));
    LocalMux I__9971 (
            .O(N__45925),
            .I(N__45904));
    LocalMux I__9970 (
            .O(N__45920),
            .I(N__45904));
    Span4Mux_h I__9969 (
            .O(N__45917),
            .I(N__45901));
    Span4Mux_h I__9968 (
            .O(N__45914),
            .I(N__45898));
    LocalMux I__9967 (
            .O(N__45911),
            .I(N__45891));
    Span4Mux_v I__9966 (
            .O(N__45904),
            .I(N__45891));
    Span4Mux_v I__9965 (
            .O(N__45901),
            .I(N__45891));
    Odrv4 I__9964 (
            .O(N__45898),
            .I(n15238));
    Odrv4 I__9963 (
            .O(N__45891),
            .I(n15238));
    CEMux I__9962 (
            .O(N__45886),
            .I(N__45882));
    InMux I__9961 (
            .O(N__45885),
            .I(N__45879));
    LocalMux I__9960 (
            .O(N__45882),
            .I(n12958));
    LocalMux I__9959 (
            .O(N__45879),
            .I(n12958));
    InMux I__9958 (
            .O(N__45874),
            .I(N__45871));
    LocalMux I__9957 (
            .O(N__45871),
            .I(N__45868));
    Odrv4 I__9956 (
            .O(N__45868),
            .I(n22397));
    InMux I__9955 (
            .O(N__45865),
            .I(N__45862));
    LocalMux I__9954 (
            .O(N__45862),
            .I(n29_adj_1688));
    CascadeMux I__9953 (
            .O(N__45859),
            .I(n11402_cascade_));
    InMux I__9952 (
            .O(N__45856),
            .I(N__45853));
    LocalMux I__9951 (
            .O(N__45853),
            .I(N__45850));
    Odrv12 I__9950 (
            .O(N__45850),
            .I(comm_state_3_N_500_2));
    CascadeMux I__9949 (
            .O(N__45847),
            .I(n22375_cascade_));
    InMux I__9948 (
            .O(N__45844),
            .I(N__45841));
    LocalMux I__9947 (
            .O(N__45841),
            .I(N__45838));
    Span4Mux_v I__9946 (
            .O(N__45838),
            .I(N__45835));
    Span4Mux_h I__9945 (
            .O(N__45835),
            .I(N__45832));
    Odrv4 I__9944 (
            .O(N__45832),
            .I(buf_data_iac_22));
    InMux I__9943 (
            .O(N__45829),
            .I(N__45826));
    LocalMux I__9942 (
            .O(N__45826),
            .I(N__45823));
    Span4Mux_h I__9941 (
            .O(N__45823),
            .I(N__45820));
    Odrv4 I__9940 (
            .O(N__45820),
            .I(n22297));
    InMux I__9939 (
            .O(N__45817),
            .I(N__45814));
    LocalMux I__9938 (
            .O(N__45814),
            .I(N__45811));
    Span4Mux_v I__9937 (
            .O(N__45811),
            .I(N__45806));
    InMux I__9936 (
            .O(N__45810),
            .I(N__45801));
    InMux I__9935 (
            .O(N__45809),
            .I(N__45801));
    Span4Mux_v I__9934 (
            .O(N__45806),
            .I(N__45794));
    LocalMux I__9933 (
            .O(N__45801),
            .I(N__45791));
    InMux I__9932 (
            .O(N__45800),
            .I(N__45784));
    InMux I__9931 (
            .O(N__45799),
            .I(N__45774));
    InMux I__9930 (
            .O(N__45798),
            .I(N__45774));
    InMux I__9929 (
            .O(N__45797),
            .I(N__45774));
    Span4Mux_h I__9928 (
            .O(N__45794),
            .I(N__45769));
    Span4Mux_h I__9927 (
            .O(N__45791),
            .I(N__45769));
    InMux I__9926 (
            .O(N__45790),
            .I(N__45760));
    InMux I__9925 (
            .O(N__45789),
            .I(N__45760));
    InMux I__9924 (
            .O(N__45788),
            .I(N__45760));
    InMux I__9923 (
            .O(N__45787),
            .I(N__45760));
    LocalMux I__9922 (
            .O(N__45784),
            .I(N__45757));
    InMux I__9921 (
            .O(N__45783),
            .I(N__45754));
    InMux I__9920 (
            .O(N__45782),
            .I(N__45749));
    InMux I__9919 (
            .O(N__45781),
            .I(N__45749));
    LocalMux I__9918 (
            .O(N__45774),
            .I(eis_state_1));
    Odrv4 I__9917 (
            .O(N__45769),
            .I(eis_state_1));
    LocalMux I__9916 (
            .O(N__45760),
            .I(eis_state_1));
    Odrv4 I__9915 (
            .O(N__45757),
            .I(eis_state_1));
    LocalMux I__9914 (
            .O(N__45754),
            .I(eis_state_1));
    LocalMux I__9913 (
            .O(N__45749),
            .I(eis_state_1));
    SRMux I__9912 (
            .O(N__45736),
            .I(N__45733));
    LocalMux I__9911 (
            .O(N__45733),
            .I(N__45730));
    Odrv12 I__9910 (
            .O(N__45730),
            .I(n15517));
    InMux I__9909 (
            .O(N__45727),
            .I(N__45724));
    LocalMux I__9908 (
            .O(N__45724),
            .I(N__45721));
    Span4Mux_h I__9907 (
            .O(N__45721),
            .I(N__45718));
    Odrv4 I__9906 (
            .O(N__45718),
            .I(comm_buf_3_5));
    CascadeMux I__9905 (
            .O(N__45715),
            .I(N__45711));
    InMux I__9904 (
            .O(N__45714),
            .I(N__45708));
    InMux I__9903 (
            .O(N__45711),
            .I(N__45705));
    LocalMux I__9902 (
            .O(N__45708),
            .I(comm_buf_6_5));
    LocalMux I__9901 (
            .O(N__45705),
            .I(comm_buf_6_5));
    InMux I__9900 (
            .O(N__45700),
            .I(N__45696));
    InMux I__9899 (
            .O(N__45699),
            .I(N__45692));
    LocalMux I__9898 (
            .O(N__45696),
            .I(N__45689));
    InMux I__9897 (
            .O(N__45695),
            .I(N__45686));
    LocalMux I__9896 (
            .O(N__45692),
            .I(N__45683));
    Span4Mux_v I__9895 (
            .O(N__45689),
            .I(N__45678));
    LocalMux I__9894 (
            .O(N__45686),
            .I(N__45678));
    Span4Mux_v I__9893 (
            .O(N__45683),
            .I(N__45675));
    Span4Mux_h I__9892 (
            .O(N__45678),
            .I(N__45672));
    Odrv4 I__9891 (
            .O(N__45675),
            .I(comm_buf_2_5));
    Odrv4 I__9890 (
            .O(N__45672),
            .I(comm_buf_2_5));
    InMux I__9889 (
            .O(N__45667),
            .I(N__45664));
    LocalMux I__9888 (
            .O(N__45664),
            .I(n18882));
    CascadeMux I__9887 (
            .O(N__45661),
            .I(n18883_cascade_));
    InMux I__9886 (
            .O(N__45658),
            .I(N__45654));
    InMux I__9885 (
            .O(N__45657),
            .I(N__45650));
    LocalMux I__9884 (
            .O(N__45654),
            .I(N__45647));
    InMux I__9883 (
            .O(N__45653),
            .I(N__45644));
    LocalMux I__9882 (
            .O(N__45650),
            .I(N__45641));
    Span4Mux_v I__9881 (
            .O(N__45647),
            .I(N__45636));
    LocalMux I__9880 (
            .O(N__45644),
            .I(N__45636));
    Span12Mux_v I__9879 (
            .O(N__45641),
            .I(N__45633));
    Span4Mux_h I__9878 (
            .O(N__45636),
            .I(N__45630));
    Odrv12 I__9877 (
            .O(N__45633),
            .I(comm_tx_buf_5));
    Odrv4 I__9876 (
            .O(N__45630),
            .I(comm_tx_buf_5));
    InMux I__9875 (
            .O(N__45625),
            .I(N__45622));
    LocalMux I__9874 (
            .O(N__45622),
            .I(N__45619));
    Odrv4 I__9873 (
            .O(N__45619),
            .I(comm_buf_5_5));
    InMux I__9872 (
            .O(N__45616),
            .I(N__45613));
    LocalMux I__9871 (
            .O(N__45613),
            .I(n22371));
    CascadeMux I__9870 (
            .O(N__45610),
            .I(n18885_cascade_));
    InMux I__9869 (
            .O(N__45607),
            .I(N__45604));
    LocalMux I__9868 (
            .O(N__45604),
            .I(n23414));
    InMux I__9867 (
            .O(N__45601),
            .I(N__45598));
    LocalMux I__9866 (
            .O(N__45598),
            .I(N__45595));
    Span4Mux_v I__9865 (
            .O(N__45595),
            .I(N__45592));
    Span4Mux_h I__9864 (
            .O(N__45592),
            .I(N__45589));
    Odrv4 I__9863 (
            .O(N__45589),
            .I(n22618));
    InMux I__9862 (
            .O(N__45586),
            .I(N__45583));
    LocalMux I__9861 (
            .O(N__45583),
            .I(N__45580));
    Span4Mux_h I__9860 (
            .O(N__45580),
            .I(N__45577));
    Span4Mux_h I__9859 (
            .O(N__45577),
            .I(N__45574));
    Odrv4 I__9858 (
            .O(N__45574),
            .I(n8_adj_1755));
    CascadeMux I__9857 (
            .O(N__45571),
            .I(N__45566));
    InMux I__9856 (
            .O(N__45570),
            .I(N__45563));
    InMux I__9855 (
            .O(N__45569),
            .I(N__45559));
    InMux I__9854 (
            .O(N__45566),
            .I(N__45553));
    LocalMux I__9853 (
            .O(N__45563),
            .I(N__45550));
    InMux I__9852 (
            .O(N__45562),
            .I(N__45547));
    LocalMux I__9851 (
            .O(N__45559),
            .I(N__45544));
    InMux I__9850 (
            .O(N__45558),
            .I(N__45537));
    InMux I__9849 (
            .O(N__45557),
            .I(N__45537));
    InMux I__9848 (
            .O(N__45556),
            .I(N__45537));
    LocalMux I__9847 (
            .O(N__45553),
            .I(N__45532));
    Span4Mux_h I__9846 (
            .O(N__45550),
            .I(N__45532));
    LocalMux I__9845 (
            .O(N__45547),
            .I(N__45527));
    Span4Mux_v I__9844 (
            .O(N__45544),
            .I(N__45527));
    LocalMux I__9843 (
            .O(N__45537),
            .I(n12976));
    Odrv4 I__9842 (
            .O(N__45532),
            .I(n12976));
    Odrv4 I__9841 (
            .O(N__45527),
            .I(n12976));
    CascadeMux I__9840 (
            .O(N__45520),
            .I(n12976_cascade_));
    CascadeMux I__9839 (
            .O(N__45517),
            .I(N__45514));
    InMux I__9838 (
            .O(N__45514),
            .I(N__45511));
    LocalMux I__9837 (
            .O(N__45511),
            .I(N__45507));
    InMux I__9836 (
            .O(N__45510),
            .I(N__45504));
    Span4Mux_v I__9835 (
            .O(N__45507),
            .I(N__45501));
    LocalMux I__9834 (
            .O(N__45504),
            .I(comm_buf_6_2));
    Odrv4 I__9833 (
            .O(N__45501),
            .I(comm_buf_6_2));
    CascadeMux I__9832 (
            .O(N__45496),
            .I(n12_adj_1760_cascade_));
    CascadeMux I__9831 (
            .O(N__45493),
            .I(n20834_cascade_));
    InMux I__9830 (
            .O(N__45490),
            .I(N__45487));
    LocalMux I__9829 (
            .O(N__45487),
            .I(n30_adj_1681));
    InMux I__9828 (
            .O(N__45484),
            .I(N__45481));
    LocalMux I__9827 (
            .O(N__45481),
            .I(n33));
    InMux I__9826 (
            .O(N__45478),
            .I(N__45475));
    LocalMux I__9825 (
            .O(N__45475),
            .I(n32));
    CascadeMux I__9824 (
            .O(N__45472),
            .I(n34_cascade_));
    InMux I__9823 (
            .O(N__45469),
            .I(N__45466));
    LocalMux I__9822 (
            .O(N__45466),
            .I(n31_adj_1680));
    CascadeMux I__9821 (
            .O(N__45463),
            .I(n49_cascade_));
    InMux I__9820 (
            .O(N__45460),
            .I(N__45455));
    InMux I__9819 (
            .O(N__45459),
            .I(N__45451));
    InMux I__9818 (
            .O(N__45458),
            .I(N__45448));
    LocalMux I__9817 (
            .O(N__45455),
            .I(N__45445));
    InMux I__9816 (
            .O(N__45454),
            .I(N__45442));
    LocalMux I__9815 (
            .O(N__45451),
            .I(N__45437));
    LocalMux I__9814 (
            .O(N__45448),
            .I(N__45437));
    Odrv12 I__9813 (
            .O(N__45445),
            .I(\comm_spi.n24022 ));
    LocalMux I__9812 (
            .O(N__45442),
            .I(\comm_spi.n24022 ));
    Odrv4 I__9811 (
            .O(N__45437),
            .I(\comm_spi.n24022 ));
    CascadeMux I__9810 (
            .O(N__45430),
            .I(n8856_cascade_));
    CascadeMux I__9809 (
            .O(N__45427),
            .I(N__45423));
    InMux I__9808 (
            .O(N__45426),
            .I(N__45418));
    InMux I__9807 (
            .O(N__45423),
            .I(N__45415));
    InMux I__9806 (
            .O(N__45422),
            .I(N__45411));
    InMux I__9805 (
            .O(N__45421),
            .I(N__45408));
    LocalMux I__9804 (
            .O(N__45418),
            .I(N__45405));
    LocalMux I__9803 (
            .O(N__45415),
            .I(N__45402));
    InMux I__9802 (
            .O(N__45414),
            .I(N__45397));
    LocalMux I__9801 (
            .O(N__45411),
            .I(N__45394));
    LocalMux I__9800 (
            .O(N__45408),
            .I(N__45391));
    Span4Mux_v I__9799 (
            .O(N__45405),
            .I(N__45388));
    Span4Mux_h I__9798 (
            .O(N__45402),
            .I(N__45385));
    InMux I__9797 (
            .O(N__45401),
            .I(N__45380));
    InMux I__9796 (
            .O(N__45400),
            .I(N__45380));
    LocalMux I__9795 (
            .O(N__45397),
            .I(N__45373));
    Span4Mux_h I__9794 (
            .O(N__45394),
            .I(N__45373));
    Span4Mux_v I__9793 (
            .O(N__45391),
            .I(N__45373));
    Span4Mux_v I__9792 (
            .O(N__45388),
            .I(N__45369));
    Span4Mux_v I__9791 (
            .O(N__45385),
            .I(N__45366));
    LocalMux I__9790 (
            .O(N__45380),
            .I(N__45361));
    Span4Mux_h I__9789 (
            .O(N__45373),
            .I(N__45361));
    InMux I__9788 (
            .O(N__45372),
            .I(N__45358));
    Span4Mux_h I__9787 (
            .O(N__45369),
            .I(N__45355));
    Span4Mux_v I__9786 (
            .O(N__45366),
            .I(N__45352));
    Span4Mux_v I__9785 (
            .O(N__45361),
            .I(N__45349));
    LocalMux I__9784 (
            .O(N__45358),
            .I(n13273));
    Odrv4 I__9783 (
            .O(N__45355),
            .I(n13273));
    Odrv4 I__9782 (
            .O(N__45352),
            .I(n13273));
    Odrv4 I__9781 (
            .O(N__45349),
            .I(n13273));
    CascadeMux I__9780 (
            .O(N__45340),
            .I(N__45336));
    CascadeMux I__9779 (
            .O(N__45339),
            .I(N__45332));
    InMux I__9778 (
            .O(N__45336),
            .I(N__45329));
    InMux I__9777 (
            .O(N__45335),
            .I(N__45322));
    InMux I__9776 (
            .O(N__45332),
            .I(N__45319));
    LocalMux I__9775 (
            .O(N__45329),
            .I(N__45316));
    CascadeMux I__9774 (
            .O(N__45328),
            .I(N__45313));
    InMux I__9773 (
            .O(N__45327),
            .I(N__45309));
    InMux I__9772 (
            .O(N__45326),
            .I(N__45304));
    InMux I__9771 (
            .O(N__45325),
            .I(N__45304));
    LocalMux I__9770 (
            .O(N__45322),
            .I(N__45301));
    LocalMux I__9769 (
            .O(N__45319),
            .I(N__45298));
    Span4Mux_v I__9768 (
            .O(N__45316),
            .I(N__45295));
    InMux I__9767 (
            .O(N__45313),
            .I(N__45292));
    InMux I__9766 (
            .O(N__45312),
            .I(N__45289));
    LocalMux I__9765 (
            .O(N__45309),
            .I(N__45284));
    LocalMux I__9764 (
            .O(N__45304),
            .I(N__45284));
    Span4Mux_v I__9763 (
            .O(N__45301),
            .I(N__45276));
    Span4Mux_v I__9762 (
            .O(N__45298),
            .I(N__45276));
    Span4Mux_h I__9761 (
            .O(N__45295),
            .I(N__45276));
    LocalMux I__9760 (
            .O(N__45292),
            .I(N__45273));
    LocalMux I__9759 (
            .O(N__45289),
            .I(N__45270));
    Span4Mux_v I__9758 (
            .O(N__45284),
            .I(N__45267));
    InMux I__9757 (
            .O(N__45283),
            .I(N__45264));
    Sp12to4 I__9756 (
            .O(N__45276),
            .I(N__45259));
    Span12Mux_v I__9755 (
            .O(N__45273),
            .I(N__45259));
    Span4Mux_v I__9754 (
            .O(N__45270),
            .I(N__45254));
    Span4Mux_v I__9753 (
            .O(N__45267),
            .I(N__45254));
    LocalMux I__9752 (
            .O(N__45264),
            .I(comm_buf_0_5));
    Odrv12 I__9751 (
            .O(N__45259),
            .I(comm_buf_0_5));
    Odrv4 I__9750 (
            .O(N__45254),
            .I(comm_buf_0_5));
    CascadeMux I__9749 (
            .O(N__45247),
            .I(\comm_spi.imosi_cascade_ ));
    InMux I__9748 (
            .O(N__45244),
            .I(N__45241));
    LocalMux I__9747 (
            .O(N__45241),
            .I(\comm_spi.n24019 ));
    InMux I__9746 (
            .O(N__45238),
            .I(N__45235));
    LocalMux I__9745 (
            .O(N__45235),
            .I(\comm_spi.n15344 ));
    InMux I__9744 (
            .O(N__45232),
            .I(N__45229));
    LocalMux I__9743 (
            .O(N__45229),
            .I(\comm_spi.n15345 ));
    CascadeMux I__9742 (
            .O(N__45226),
            .I(\comm_spi.n24019_cascade_ ));
    InMux I__9741 (
            .O(N__45223),
            .I(N__45219));
    InMux I__9740 (
            .O(N__45222),
            .I(N__45216));
    LocalMux I__9739 (
            .O(N__45219),
            .I(N__45211));
    LocalMux I__9738 (
            .O(N__45216),
            .I(N__45211));
    Odrv4 I__9737 (
            .O(N__45211),
            .I(secclk_cnt_0));
    InMux I__9736 (
            .O(N__45208),
            .I(N__45204));
    InMux I__9735 (
            .O(N__45207),
            .I(N__45201));
    LocalMux I__9734 (
            .O(N__45204),
            .I(N__45198));
    LocalMux I__9733 (
            .O(N__45201),
            .I(N__45193));
    Span4Mux_v I__9732 (
            .O(N__45198),
            .I(N__45193));
    Odrv4 I__9731 (
            .O(N__45193),
            .I(secclk_cnt_18));
    CascadeMux I__9730 (
            .O(N__45190),
            .I(N__45187));
    InMux I__9729 (
            .O(N__45187),
            .I(N__45184));
    LocalMux I__9728 (
            .O(N__45184),
            .I(N__45180));
    InMux I__9727 (
            .O(N__45183),
            .I(N__45177));
    Span4Mux_h I__9726 (
            .O(N__45180),
            .I(N__45174));
    LocalMux I__9725 (
            .O(N__45177),
            .I(secclk_cnt_11));
    Odrv4 I__9724 (
            .O(N__45174),
            .I(secclk_cnt_11));
    InMux I__9723 (
            .O(N__45169),
            .I(N__45165));
    InMux I__9722 (
            .O(N__45168),
            .I(N__45162));
    LocalMux I__9721 (
            .O(N__45165),
            .I(N__45159));
    LocalMux I__9720 (
            .O(N__45162),
            .I(secclk_cnt_4));
    Odrv4 I__9719 (
            .O(N__45159),
            .I(secclk_cnt_4));
    InMux I__9718 (
            .O(N__45154),
            .I(N__45151));
    LocalMux I__9717 (
            .O(N__45151),
            .I(n28));
    InMux I__9716 (
            .O(N__45148),
            .I(N__45144));
    InMux I__9715 (
            .O(N__45147),
            .I(N__45141));
    LocalMux I__9714 (
            .O(N__45144),
            .I(N__45136));
    LocalMux I__9713 (
            .O(N__45141),
            .I(N__45136));
    Span4Mux_h I__9712 (
            .O(N__45136),
            .I(N__45132));
    InMux I__9711 (
            .O(N__45135),
            .I(N__45129));
    Span4Mux_v I__9710 (
            .O(N__45132),
            .I(N__45126));
    LocalMux I__9709 (
            .O(N__45129),
            .I(data_index_6));
    Odrv4 I__9708 (
            .O(N__45126),
            .I(data_index_6));
    InMux I__9707 (
            .O(N__45121),
            .I(N__45118));
    LocalMux I__9706 (
            .O(N__45118),
            .I(n8_adj_1621));
    CascadeMux I__9705 (
            .O(N__45115),
            .I(n8_adj_1621_cascade_));
    InMux I__9704 (
            .O(N__45112),
            .I(N__45106));
    InMux I__9703 (
            .O(N__45111),
            .I(N__45106));
    LocalMux I__9702 (
            .O(N__45106),
            .I(N__45103));
    Span4Mux_v I__9701 (
            .O(N__45103),
            .I(N__45100));
    Odrv4 I__9700 (
            .O(N__45100),
            .I(n7_adj_1620));
    CascadeMux I__9699 (
            .O(N__45097),
            .I(N__45094));
    CascadeBuf I__9698 (
            .O(N__45094),
            .I(N__45091));
    CascadeMux I__9697 (
            .O(N__45091),
            .I(N__45088));
    CascadeBuf I__9696 (
            .O(N__45088),
            .I(N__45085));
    CascadeMux I__9695 (
            .O(N__45085),
            .I(N__45082));
    CascadeBuf I__9694 (
            .O(N__45082),
            .I(N__45079));
    CascadeMux I__9693 (
            .O(N__45079),
            .I(N__45076));
    CascadeBuf I__9692 (
            .O(N__45076),
            .I(N__45073));
    CascadeMux I__9691 (
            .O(N__45073),
            .I(N__45070));
    CascadeBuf I__9690 (
            .O(N__45070),
            .I(N__45067));
    CascadeMux I__9689 (
            .O(N__45067),
            .I(N__45064));
    CascadeBuf I__9688 (
            .O(N__45064),
            .I(N__45061));
    CascadeMux I__9687 (
            .O(N__45061),
            .I(N__45058));
    CascadeBuf I__9686 (
            .O(N__45058),
            .I(N__45054));
    CascadeMux I__9685 (
            .O(N__45057),
            .I(N__45051));
    CascadeMux I__9684 (
            .O(N__45054),
            .I(N__45048));
    CascadeBuf I__9683 (
            .O(N__45051),
            .I(N__45045));
    CascadeBuf I__9682 (
            .O(N__45048),
            .I(N__45042));
    CascadeMux I__9681 (
            .O(N__45045),
            .I(N__45039));
    CascadeMux I__9680 (
            .O(N__45042),
            .I(N__45036));
    InMux I__9679 (
            .O(N__45039),
            .I(N__45033));
    CascadeBuf I__9678 (
            .O(N__45036),
            .I(N__45030));
    LocalMux I__9677 (
            .O(N__45033),
            .I(N__45027));
    CascadeMux I__9676 (
            .O(N__45030),
            .I(N__45024));
    Span12Mux_s10_h I__9675 (
            .O(N__45027),
            .I(N__45021));
    InMux I__9674 (
            .O(N__45024),
            .I(N__45018));
    Span12Mux_v I__9673 (
            .O(N__45021),
            .I(N__45015));
    LocalMux I__9672 (
            .O(N__45018),
            .I(N__45012));
    Odrv12 I__9671 (
            .O(N__45015),
            .I(data_index_9_N_236_6));
    Odrv12 I__9670 (
            .O(N__45012),
            .I(data_index_9_N_236_6));
    InMux I__9669 (
            .O(N__45007),
            .I(N__45003));
    InMux I__9668 (
            .O(N__45006),
            .I(N__45000));
    LocalMux I__9667 (
            .O(N__45003),
            .I(N__44994));
    LocalMux I__9666 (
            .O(N__45000),
            .I(N__44994));
    InMux I__9665 (
            .O(N__44999),
            .I(N__44991));
    Span4Mux_h I__9664 (
            .O(N__44994),
            .I(N__44988));
    LocalMux I__9663 (
            .O(N__44991),
            .I(N__44983));
    Span4Mux_h I__9662 (
            .O(N__44988),
            .I(N__44983));
    Odrv4 I__9661 (
            .O(N__44983),
            .I(data_index_7));
    InMux I__9660 (
            .O(N__44980),
            .I(N__44977));
    LocalMux I__9659 (
            .O(N__44977),
            .I(N__44974));
    Odrv4 I__9658 (
            .O(N__44974),
            .I(n8_adj_1617));
    InMux I__9657 (
            .O(N__44971),
            .I(N__44967));
    InMux I__9656 (
            .O(N__44970),
            .I(N__44964));
    LocalMux I__9655 (
            .O(N__44967),
            .I(N__44959));
    LocalMux I__9654 (
            .O(N__44964),
            .I(N__44959));
    Span4Mux_v I__9653 (
            .O(N__44959),
            .I(N__44956));
    Odrv4 I__9652 (
            .O(N__44956),
            .I(n7_adj_1616));
    InMux I__9651 (
            .O(N__44953),
            .I(N__44949));
    InMux I__9650 (
            .O(N__44952),
            .I(N__44946));
    LocalMux I__9649 (
            .O(N__44949),
            .I(N__44941));
    LocalMux I__9648 (
            .O(N__44946),
            .I(N__44941));
    Span4Mux_v I__9647 (
            .O(N__44941),
            .I(N__44937));
    InMux I__9646 (
            .O(N__44940),
            .I(N__44934));
    Span4Mux_h I__9645 (
            .O(N__44937),
            .I(N__44931));
    LocalMux I__9644 (
            .O(N__44934),
            .I(data_index_8));
    Odrv4 I__9643 (
            .O(N__44931),
            .I(data_index_8));
    InMux I__9642 (
            .O(N__44926),
            .I(N__44920));
    InMux I__9641 (
            .O(N__44925),
            .I(N__44920));
    LocalMux I__9640 (
            .O(N__44920),
            .I(n8_adj_1619));
    InMux I__9639 (
            .O(N__44917),
            .I(N__44911));
    InMux I__9638 (
            .O(N__44916),
            .I(N__44911));
    LocalMux I__9637 (
            .O(N__44911),
            .I(N__44908));
    Span4Mux_v I__9636 (
            .O(N__44908),
            .I(N__44905));
    Odrv4 I__9635 (
            .O(N__44905),
            .I(n7_adj_1618));
    CascadeMux I__9634 (
            .O(N__44902),
            .I(N__44899));
    CascadeBuf I__9633 (
            .O(N__44899),
            .I(N__44896));
    CascadeMux I__9632 (
            .O(N__44896),
            .I(N__44893));
    CascadeBuf I__9631 (
            .O(N__44893),
            .I(N__44890));
    CascadeMux I__9630 (
            .O(N__44890),
            .I(N__44887));
    CascadeBuf I__9629 (
            .O(N__44887),
            .I(N__44884));
    CascadeMux I__9628 (
            .O(N__44884),
            .I(N__44881));
    CascadeBuf I__9627 (
            .O(N__44881),
            .I(N__44878));
    CascadeMux I__9626 (
            .O(N__44878),
            .I(N__44875));
    CascadeBuf I__9625 (
            .O(N__44875),
            .I(N__44872));
    CascadeMux I__9624 (
            .O(N__44872),
            .I(N__44869));
    CascadeBuf I__9623 (
            .O(N__44869),
            .I(N__44866));
    CascadeMux I__9622 (
            .O(N__44866),
            .I(N__44863));
    CascadeBuf I__9621 (
            .O(N__44863),
            .I(N__44859));
    CascadeMux I__9620 (
            .O(N__44862),
            .I(N__44856));
    CascadeMux I__9619 (
            .O(N__44859),
            .I(N__44853));
    CascadeBuf I__9618 (
            .O(N__44856),
            .I(N__44850));
    CascadeBuf I__9617 (
            .O(N__44853),
            .I(N__44847));
    CascadeMux I__9616 (
            .O(N__44850),
            .I(N__44844));
    CascadeMux I__9615 (
            .O(N__44847),
            .I(N__44841));
    InMux I__9614 (
            .O(N__44844),
            .I(N__44838));
    CascadeBuf I__9613 (
            .O(N__44841),
            .I(N__44835));
    LocalMux I__9612 (
            .O(N__44838),
            .I(N__44832));
    CascadeMux I__9611 (
            .O(N__44835),
            .I(N__44829));
    Span12Mux_h I__9610 (
            .O(N__44832),
            .I(N__44826));
    InMux I__9609 (
            .O(N__44829),
            .I(N__44823));
    Span12Mux_v I__9608 (
            .O(N__44826),
            .I(N__44820));
    LocalMux I__9607 (
            .O(N__44823),
            .I(N__44817));
    Odrv12 I__9606 (
            .O(N__44820),
            .I(data_index_9_N_236_7));
    Odrv12 I__9605 (
            .O(N__44817),
            .I(data_index_9_N_236_7));
    InMux I__9604 (
            .O(N__44812),
            .I(N__44809));
    LocalMux I__9603 (
            .O(N__44809),
            .I(\SIG_DDS.n22671 ));
    CascadeMux I__9602 (
            .O(N__44806),
            .I(N__44803));
    InMux I__9601 (
            .O(N__44803),
            .I(N__44800));
    LocalMux I__9600 (
            .O(N__44800),
            .I(N__44797));
    Odrv4 I__9599 (
            .O(N__44797),
            .I(\SIG_DDS.n10 ));
    SRMux I__9598 (
            .O(N__44794),
            .I(N__44791));
    LocalMux I__9597 (
            .O(N__44791),
            .I(N__44788));
    Odrv12 I__9596 (
            .O(N__44788),
            .I(\comm_spi.imosi_N_841 ));
    InMux I__9595 (
            .O(N__44785),
            .I(N__44780));
    InMux I__9594 (
            .O(N__44784),
            .I(N__44777));
    InMux I__9593 (
            .O(N__44783),
            .I(N__44774));
    LocalMux I__9592 (
            .O(N__44780),
            .I(N__44769));
    LocalMux I__9591 (
            .O(N__44777),
            .I(N__44769));
    LocalMux I__9590 (
            .O(N__44774),
            .I(\comm_spi.n15331 ));
    Odrv4 I__9589 (
            .O(N__44769),
            .I(\comm_spi.n15331 ));
    CascadeMux I__9588 (
            .O(N__44764),
            .I(N__44760));
    CascadeMux I__9587 (
            .O(N__44763),
            .I(N__44756));
    InMux I__9586 (
            .O(N__44760),
            .I(N__44751));
    InMux I__9585 (
            .O(N__44759),
            .I(N__44751));
    InMux I__9584 (
            .O(N__44756),
            .I(N__44748));
    LocalMux I__9583 (
            .O(N__44751),
            .I(\SIG_DDS.bit_cnt_2 ));
    LocalMux I__9582 (
            .O(N__44748),
            .I(\SIG_DDS.bit_cnt_2 ));
    CascadeMux I__9581 (
            .O(N__44743),
            .I(N__44739));
    InMux I__9580 (
            .O(N__44742),
            .I(N__44734));
    InMux I__9579 (
            .O(N__44739),
            .I(N__44729));
    InMux I__9578 (
            .O(N__44738),
            .I(N__44729));
    InMux I__9577 (
            .O(N__44737),
            .I(N__44726));
    LocalMux I__9576 (
            .O(N__44734),
            .I(\SIG_DDS.bit_cnt_1 ));
    LocalMux I__9575 (
            .O(N__44729),
            .I(\SIG_DDS.bit_cnt_1 ));
    LocalMux I__9574 (
            .O(N__44726),
            .I(\SIG_DDS.bit_cnt_1 ));
    CascadeMux I__9573 (
            .O(N__44719),
            .I(N__44716));
    InMux I__9572 (
            .O(N__44716),
            .I(N__44711));
    InMux I__9571 (
            .O(N__44715),
            .I(N__44708));
    InMux I__9570 (
            .O(N__44714),
            .I(N__44704));
    LocalMux I__9569 (
            .O(N__44711),
            .I(N__44700));
    LocalMux I__9568 (
            .O(N__44708),
            .I(N__44697));
    CascadeMux I__9567 (
            .O(N__44707),
            .I(N__44694));
    LocalMux I__9566 (
            .O(N__44704),
            .I(N__44690));
    InMux I__9565 (
            .O(N__44703),
            .I(N__44687));
    Span4Mux_h I__9564 (
            .O(N__44700),
            .I(N__44684));
    Span4Mux_v I__9563 (
            .O(N__44697),
            .I(N__44681));
    InMux I__9562 (
            .O(N__44694),
            .I(N__44678));
    CascadeMux I__9561 (
            .O(N__44693),
            .I(N__44674));
    Span4Mux_h I__9560 (
            .O(N__44690),
            .I(N__44665));
    LocalMux I__9559 (
            .O(N__44687),
            .I(N__44665));
    Span4Mux_h I__9558 (
            .O(N__44684),
            .I(N__44665));
    Span4Mux_h I__9557 (
            .O(N__44681),
            .I(N__44665));
    LocalMux I__9556 (
            .O(N__44678),
            .I(N__44662));
    InMux I__9555 (
            .O(N__44677),
            .I(N__44657));
    InMux I__9554 (
            .O(N__44674),
            .I(N__44657));
    Span4Mux_v I__9553 (
            .O(N__44665),
            .I(N__44654));
    Odrv12 I__9552 (
            .O(N__44662),
            .I(comm_buf_0_4));
    LocalMux I__9551 (
            .O(N__44657),
            .I(comm_buf_0_4));
    Odrv4 I__9550 (
            .O(N__44654),
            .I(comm_buf_0_4));
    CascadeMux I__9549 (
            .O(N__44647),
            .I(N__44643));
    CascadeMux I__9548 (
            .O(N__44646),
            .I(N__44639));
    InMux I__9547 (
            .O(N__44643),
            .I(N__44636));
    InMux I__9546 (
            .O(N__44642),
            .I(N__44633));
    InMux I__9545 (
            .O(N__44639),
            .I(N__44627));
    LocalMux I__9544 (
            .O(N__44636),
            .I(N__44624));
    LocalMux I__9543 (
            .O(N__44633),
            .I(N__44621));
    InMux I__9542 (
            .O(N__44632),
            .I(N__44618));
    CascadeMux I__9541 (
            .O(N__44631),
            .I(N__44614));
    CascadeMux I__9540 (
            .O(N__44630),
            .I(N__44610));
    LocalMux I__9539 (
            .O(N__44627),
            .I(N__44607));
    Span4Mux_v I__9538 (
            .O(N__44624),
            .I(N__44604));
    Span4Mux_v I__9537 (
            .O(N__44621),
            .I(N__44599));
    LocalMux I__9536 (
            .O(N__44618),
            .I(N__44599));
    CascadeMux I__9535 (
            .O(N__44617),
            .I(N__44596));
    InMux I__9534 (
            .O(N__44614),
            .I(N__44593));
    InMux I__9533 (
            .O(N__44613),
            .I(N__44589));
    InMux I__9532 (
            .O(N__44610),
            .I(N__44586));
    Span4Mux_v I__9531 (
            .O(N__44607),
            .I(N__44583));
    Span4Mux_v I__9530 (
            .O(N__44604),
            .I(N__44578));
    Span4Mux_h I__9529 (
            .O(N__44599),
            .I(N__44578));
    InMux I__9528 (
            .O(N__44596),
            .I(N__44575));
    LocalMux I__9527 (
            .O(N__44593),
            .I(N__44572));
    InMux I__9526 (
            .O(N__44592),
            .I(N__44569));
    LocalMux I__9525 (
            .O(N__44589),
            .I(N__44566));
    LocalMux I__9524 (
            .O(N__44586),
            .I(N__44558));
    Span4Mux_h I__9523 (
            .O(N__44583),
            .I(N__44558));
    Span4Mux_v I__9522 (
            .O(N__44578),
            .I(N__44558));
    LocalMux I__9521 (
            .O(N__44575),
            .I(N__44555));
    Span4Mux_h I__9520 (
            .O(N__44572),
            .I(N__44552));
    LocalMux I__9519 (
            .O(N__44569),
            .I(N__44549));
    Span4Mux_v I__9518 (
            .O(N__44566),
            .I(N__44546));
    InMux I__9517 (
            .O(N__44565),
            .I(N__44543));
    Span4Mux_v I__9516 (
            .O(N__44558),
            .I(N__44540));
    Odrv12 I__9515 (
            .O(N__44555),
            .I(comm_buf_0_1));
    Odrv4 I__9514 (
            .O(N__44552),
            .I(comm_buf_0_1));
    Odrv4 I__9513 (
            .O(N__44549),
            .I(comm_buf_0_1));
    Odrv4 I__9512 (
            .O(N__44546),
            .I(comm_buf_0_1));
    LocalMux I__9511 (
            .O(N__44543),
            .I(comm_buf_0_1));
    Odrv4 I__9510 (
            .O(N__44540),
            .I(comm_buf_0_1));
    InMux I__9509 (
            .O(N__44527),
            .I(N__44523));
    InMux I__9508 (
            .O(N__44526),
            .I(N__44520));
    LocalMux I__9507 (
            .O(N__44523),
            .I(\SIG_DDS.bit_cnt_3 ));
    LocalMux I__9506 (
            .O(N__44520),
            .I(\SIG_DDS.bit_cnt_3 ));
    InMux I__9505 (
            .O(N__44515),
            .I(N__44512));
    LocalMux I__9504 (
            .O(N__44512),
            .I(N__44509));
    Span4Mux_h I__9503 (
            .O(N__44509),
            .I(N__44505));
    InMux I__9502 (
            .O(N__44508),
            .I(N__44502));
    Odrv4 I__9501 (
            .O(N__44505),
            .I(n8_adj_1615));
    LocalMux I__9500 (
            .O(N__44502),
            .I(n8_adj_1615));
    InMux I__9499 (
            .O(N__44497),
            .I(N__44493));
    InMux I__9498 (
            .O(N__44496),
            .I(N__44490));
    LocalMux I__9497 (
            .O(N__44493),
            .I(N__44487));
    LocalMux I__9496 (
            .O(N__44490),
            .I(N__44484));
    Span4Mux_v I__9495 (
            .O(N__44487),
            .I(N__44479));
    Span4Mux_v I__9494 (
            .O(N__44484),
            .I(N__44479));
    Odrv4 I__9493 (
            .O(N__44479),
            .I(n7_adj_1614));
    CascadeMux I__9492 (
            .O(N__44476),
            .I(N__44473));
    CascadeBuf I__9491 (
            .O(N__44473),
            .I(N__44470));
    CascadeMux I__9490 (
            .O(N__44470),
            .I(N__44467));
    CascadeBuf I__9489 (
            .O(N__44467),
            .I(N__44464));
    CascadeMux I__9488 (
            .O(N__44464),
            .I(N__44461));
    CascadeBuf I__9487 (
            .O(N__44461),
            .I(N__44458));
    CascadeMux I__9486 (
            .O(N__44458),
            .I(N__44455));
    CascadeBuf I__9485 (
            .O(N__44455),
            .I(N__44452));
    CascadeMux I__9484 (
            .O(N__44452),
            .I(N__44449));
    CascadeBuf I__9483 (
            .O(N__44449),
            .I(N__44446));
    CascadeMux I__9482 (
            .O(N__44446),
            .I(N__44443));
    CascadeBuf I__9481 (
            .O(N__44443),
            .I(N__44440));
    CascadeMux I__9480 (
            .O(N__44440),
            .I(N__44437));
    CascadeBuf I__9479 (
            .O(N__44437),
            .I(N__44434));
    CascadeMux I__9478 (
            .O(N__44434),
            .I(N__44430));
    CascadeMux I__9477 (
            .O(N__44433),
            .I(N__44427));
    CascadeBuf I__9476 (
            .O(N__44430),
            .I(N__44424));
    CascadeBuf I__9475 (
            .O(N__44427),
            .I(N__44421));
    CascadeMux I__9474 (
            .O(N__44424),
            .I(N__44418));
    CascadeMux I__9473 (
            .O(N__44421),
            .I(N__44415));
    CascadeBuf I__9472 (
            .O(N__44418),
            .I(N__44412));
    InMux I__9471 (
            .O(N__44415),
            .I(N__44409));
    CascadeMux I__9470 (
            .O(N__44412),
            .I(N__44406));
    LocalMux I__9469 (
            .O(N__44409),
            .I(N__44403));
    InMux I__9468 (
            .O(N__44406),
            .I(N__44400));
    Span12Mux_h I__9467 (
            .O(N__44403),
            .I(N__44397));
    LocalMux I__9466 (
            .O(N__44400),
            .I(N__44394));
    Span12Mux_v I__9465 (
            .O(N__44397),
            .I(N__44391));
    Span4Mux_h I__9464 (
            .O(N__44394),
            .I(N__44388));
    Odrv12 I__9463 (
            .O(N__44391),
            .I(data_index_9_N_236_9));
    Odrv4 I__9462 (
            .O(N__44388),
            .I(data_index_9_N_236_9));
    InMux I__9461 (
            .O(N__44383),
            .I(N__44378));
    InMux I__9460 (
            .O(N__44382),
            .I(N__44375));
    InMux I__9459 (
            .O(N__44381),
            .I(N__44372));
    LocalMux I__9458 (
            .O(N__44378),
            .I(req_data_cnt_15));
    LocalMux I__9457 (
            .O(N__44375),
            .I(req_data_cnt_15));
    LocalMux I__9456 (
            .O(N__44372),
            .I(req_data_cnt_15));
    InMux I__9455 (
            .O(N__44365),
            .I(N__44362));
    LocalMux I__9454 (
            .O(N__44362),
            .I(N__44359));
    Span4Mux_h I__9453 (
            .O(N__44359),
            .I(N__44356));
    Span4Mux_h I__9452 (
            .O(N__44356),
            .I(N__44353));
    Odrv4 I__9451 (
            .O(N__44353),
            .I(n22314));
    InMux I__9450 (
            .O(N__44350),
            .I(N__44347));
    LocalMux I__9449 (
            .O(N__44347),
            .I(n22169));
    InMux I__9448 (
            .O(N__44344),
            .I(N__44341));
    LocalMux I__9447 (
            .O(N__44341),
            .I(N__44337));
    InMux I__9446 (
            .O(N__44340),
            .I(N__44333));
    Span12Mux_h I__9445 (
            .O(N__44337),
            .I(N__44330));
    InMux I__9444 (
            .O(N__44336),
            .I(N__44327));
    LocalMux I__9443 (
            .O(N__44333),
            .I(req_data_cnt_3));
    Odrv12 I__9442 (
            .O(N__44330),
            .I(req_data_cnt_3));
    LocalMux I__9441 (
            .O(N__44327),
            .I(req_data_cnt_3));
    CascadeMux I__9440 (
            .O(N__44320),
            .I(n23312_cascade_));
    CascadeMux I__9439 (
            .O(N__44317),
            .I(n23315_cascade_));
    InMux I__9438 (
            .O(N__44314),
            .I(N__44311));
    LocalMux I__9437 (
            .O(N__44311),
            .I(N__44308));
    Sp12to4 I__9436 (
            .O(N__44308),
            .I(N__44305));
    Span12Mux_v I__9435 (
            .O(N__44305),
            .I(N__44302));
    Odrv12 I__9434 (
            .O(N__44302),
            .I(n111_adj_1744));
    CascadeMux I__9433 (
            .O(N__44299),
            .I(n30_adj_1741_cascade_));
    CascadeMux I__9432 (
            .O(N__44296),
            .I(N__44292));
    CascadeMux I__9431 (
            .O(N__44295),
            .I(N__44289));
    InMux I__9430 (
            .O(N__44292),
            .I(N__44285));
    InMux I__9429 (
            .O(N__44289),
            .I(N__44280));
    InMux I__9428 (
            .O(N__44288),
            .I(N__44280));
    LocalMux I__9427 (
            .O(N__44285),
            .I(N__44277));
    LocalMux I__9426 (
            .O(N__44280),
            .I(acadc_skipCount_3));
    Odrv4 I__9425 (
            .O(N__44277),
            .I(acadc_skipCount_3));
    InMux I__9424 (
            .O(N__44272),
            .I(N__44269));
    LocalMux I__9423 (
            .O(N__44269),
            .I(N__44266));
    Span4Mux_v I__9422 (
            .O(N__44266),
            .I(N__44263));
    Odrv4 I__9421 (
            .O(N__44263),
            .I(n19_adj_1739));
    CascadeMux I__9420 (
            .O(N__44260),
            .I(N__44257));
    InMux I__9419 (
            .O(N__44257),
            .I(N__44254));
    LocalMux I__9418 (
            .O(N__44254),
            .I(N__44251));
    Span4Mux_h I__9417 (
            .O(N__44251),
            .I(N__44248));
    Sp12to4 I__9416 (
            .O(N__44248),
            .I(N__44244));
    CascadeMux I__9415 (
            .O(N__44247),
            .I(N__44241));
    Span12Mux_v I__9414 (
            .O(N__44244),
            .I(N__44238));
    InMux I__9413 (
            .O(N__44241),
            .I(N__44235));
    Odrv12 I__9412 (
            .O(N__44238),
            .I(buf_readRTD_3));
    LocalMux I__9411 (
            .O(N__44235),
            .I(buf_readRTD_3));
    InMux I__9410 (
            .O(N__44230),
            .I(N__44225));
    InMux I__9409 (
            .O(N__44229),
            .I(N__44222));
    CascadeMux I__9408 (
            .O(N__44228),
            .I(N__44219));
    LocalMux I__9407 (
            .O(N__44225),
            .I(N__44214));
    LocalMux I__9406 (
            .O(N__44222),
            .I(N__44214));
    InMux I__9405 (
            .O(N__44219),
            .I(N__44211));
    Span12Mux_h I__9404 (
            .O(N__44214),
            .I(N__44208));
    LocalMux I__9403 (
            .O(N__44211),
            .I(buf_adcdata_iac_11));
    Odrv12 I__9402 (
            .O(N__44208),
            .I(buf_adcdata_iac_11));
    InMux I__9401 (
            .O(N__44203),
            .I(N__44200));
    LocalMux I__9400 (
            .O(N__44200),
            .I(N__44197));
    Span4Mux_h I__9399 (
            .O(N__44197),
            .I(N__44194));
    Odrv4 I__9398 (
            .O(N__44194),
            .I(n16_adj_1738));
    CascadeMux I__9397 (
            .O(N__44191),
            .I(n23558_cascade_));
    InMux I__9396 (
            .O(N__44188),
            .I(N__44185));
    LocalMux I__9395 (
            .O(N__44185),
            .I(n23561));
    InMux I__9394 (
            .O(N__44182),
            .I(N__44176));
    InMux I__9393 (
            .O(N__44181),
            .I(N__44176));
    LocalMux I__9392 (
            .O(N__44176),
            .I(N__44173));
    Odrv4 I__9391 (
            .O(N__44173),
            .I(n7_adj_1624));
    InMux I__9390 (
            .O(N__44170),
            .I(N__44167));
    LocalMux I__9389 (
            .O(N__44167),
            .I(n8_adj_1625));
    InMux I__9388 (
            .O(N__44164),
            .I(N__44160));
    InMux I__9387 (
            .O(N__44163),
            .I(N__44157));
    LocalMux I__9386 (
            .O(N__44160),
            .I(N__44151));
    LocalMux I__9385 (
            .O(N__44157),
            .I(N__44151));
    InMux I__9384 (
            .O(N__44156),
            .I(N__44148));
    Span4Mux_h I__9383 (
            .O(N__44151),
            .I(N__44145));
    LocalMux I__9382 (
            .O(N__44148),
            .I(data_index_4));
    Odrv4 I__9381 (
            .O(N__44145),
            .I(data_index_4));
    InMux I__9380 (
            .O(N__44140),
            .I(N__44137));
    LocalMux I__9379 (
            .O(N__44137),
            .I(n23546));
    InMux I__9378 (
            .O(N__44134),
            .I(N__44131));
    LocalMux I__9377 (
            .O(N__44131),
            .I(n30));
    InMux I__9376 (
            .O(N__44128),
            .I(N__44125));
    LocalMux I__9375 (
            .O(N__44125),
            .I(N__44122));
    Span4Mux_h I__9374 (
            .O(N__44122),
            .I(N__44119));
    Odrv4 I__9373 (
            .O(N__44119),
            .I(n17_adj_1594));
    InMux I__9372 (
            .O(N__44116),
            .I(N__44112));
    InMux I__9371 (
            .O(N__44115),
            .I(N__44109));
    LocalMux I__9370 (
            .O(N__44112),
            .I(N__44106));
    LocalMux I__9369 (
            .O(N__44109),
            .I(N__44100));
    Span4Mux_h I__9368 (
            .O(N__44106),
            .I(N__44100));
    InMux I__9367 (
            .O(N__44105),
            .I(N__44097));
    Odrv4 I__9366 (
            .O(N__44100),
            .I(acadc_skipCount_8));
    LocalMux I__9365 (
            .O(N__44097),
            .I(acadc_skipCount_8));
    CascadeMux I__9364 (
            .O(N__44092),
            .I(N__44089));
    InMux I__9363 (
            .O(N__44089),
            .I(N__44086));
    LocalMux I__9362 (
            .O(N__44086),
            .I(N__44083));
    Odrv4 I__9361 (
            .O(N__44083),
            .I(n24_adj_1800));
    InMux I__9360 (
            .O(N__44080),
            .I(N__44075));
    CascadeMux I__9359 (
            .O(N__44079),
            .I(N__44072));
    InMux I__9358 (
            .O(N__44078),
            .I(N__44069));
    LocalMux I__9357 (
            .O(N__44075),
            .I(N__44066));
    InMux I__9356 (
            .O(N__44072),
            .I(N__44063));
    LocalMux I__9355 (
            .O(N__44069),
            .I(req_data_cnt_9));
    Odrv4 I__9354 (
            .O(N__44066),
            .I(req_data_cnt_9));
    LocalMux I__9353 (
            .O(N__44063),
            .I(req_data_cnt_9));
    InMux I__9352 (
            .O(N__44056),
            .I(N__44053));
    LocalMux I__9351 (
            .O(N__44053),
            .I(N__44050));
    Sp12to4 I__9350 (
            .O(N__44050),
            .I(N__44047));
    Odrv12 I__9349 (
            .O(N__44047),
            .I(n18_adj_1699));
    CEMux I__9348 (
            .O(N__44044),
            .I(N__44041));
    LocalMux I__9347 (
            .O(N__44041),
            .I(N__44037));
    CascadeMux I__9346 (
            .O(N__44040),
            .I(N__44034));
    Span4Mux_h I__9345 (
            .O(N__44037),
            .I(N__44031));
    InMux I__9344 (
            .O(N__44034),
            .I(N__44028));
    Span4Mux_h I__9343 (
            .O(N__44031),
            .I(N__44025));
    LocalMux I__9342 (
            .O(N__44028),
            .I(N__44022));
    Odrv4 I__9341 (
            .O(N__44025),
            .I(n13257));
    Odrv4 I__9340 (
            .O(N__44022),
            .I(n13257));
    InMux I__9339 (
            .O(N__44017),
            .I(N__44014));
    LocalMux I__9338 (
            .O(N__44014),
            .I(N__44011));
    Span4Mux_v I__9337 (
            .O(N__44011),
            .I(N__44007));
    InMux I__9336 (
            .O(N__44010),
            .I(N__44004));
    Span4Mux_h I__9335 (
            .O(N__44007),
            .I(N__44001));
    LocalMux I__9334 (
            .O(N__44004),
            .I(acadc_skipcnt_1));
    Odrv4 I__9333 (
            .O(N__44001),
            .I(acadc_skipcnt_1));
    CascadeMux I__9332 (
            .O(N__43996),
            .I(N__43993));
    InMux I__9331 (
            .O(N__43993),
            .I(N__43990));
    LocalMux I__9330 (
            .O(N__43990),
            .I(N__43987));
    Span4Mux_v I__9329 (
            .O(N__43987),
            .I(N__43983));
    InMux I__9328 (
            .O(N__43986),
            .I(N__43980));
    Span4Mux_v I__9327 (
            .O(N__43983),
            .I(N__43977));
    LocalMux I__9326 (
            .O(N__43980),
            .I(acadc_skipcnt_4));
    Odrv4 I__9325 (
            .O(N__43977),
            .I(acadc_skipcnt_4));
    InMux I__9324 (
            .O(N__43972),
            .I(N__43969));
    LocalMux I__9323 (
            .O(N__43969),
            .I(N__43966));
    Span4Mux_h I__9322 (
            .O(N__43966),
            .I(N__43963));
    Odrv4 I__9321 (
            .O(N__43963),
            .I(n18));
    InMux I__9320 (
            .O(N__43960),
            .I(N__43957));
    LocalMux I__9319 (
            .O(N__43957),
            .I(N__43952));
    CascadeMux I__9318 (
            .O(N__43956),
            .I(N__43949));
    InMux I__9317 (
            .O(N__43955),
            .I(N__43944));
    Span4Mux_h I__9316 (
            .O(N__43952),
            .I(N__43941));
    InMux I__9315 (
            .O(N__43949),
            .I(N__43934));
    InMux I__9314 (
            .O(N__43948),
            .I(N__43934));
    InMux I__9313 (
            .O(N__43947),
            .I(N__43930));
    LocalMux I__9312 (
            .O(N__43944),
            .I(N__43927));
    Span4Mux_h I__9311 (
            .O(N__43941),
            .I(N__43924));
    CascadeMux I__9310 (
            .O(N__43940),
            .I(N__43921));
    InMux I__9309 (
            .O(N__43939),
            .I(N__43918));
    LocalMux I__9308 (
            .O(N__43934),
            .I(N__43915));
    InMux I__9307 (
            .O(N__43933),
            .I(N__43911));
    LocalMux I__9306 (
            .O(N__43930),
            .I(N__43908));
    Span4Mux_h I__9305 (
            .O(N__43927),
            .I(N__43905));
    Span4Mux_v I__9304 (
            .O(N__43924),
            .I(N__43902));
    InMux I__9303 (
            .O(N__43921),
            .I(N__43899));
    LocalMux I__9302 (
            .O(N__43918),
            .I(N__43894));
    Span4Mux_h I__9301 (
            .O(N__43915),
            .I(N__43894));
    InMux I__9300 (
            .O(N__43914),
            .I(N__43891));
    LocalMux I__9299 (
            .O(N__43911),
            .I(N__43886));
    Span12Mux_h I__9298 (
            .O(N__43908),
            .I(N__43886));
    Odrv4 I__9297 (
            .O(N__43905),
            .I(comm_buf_0_0));
    Odrv4 I__9296 (
            .O(N__43902),
            .I(comm_buf_0_0));
    LocalMux I__9295 (
            .O(N__43899),
            .I(comm_buf_0_0));
    Odrv4 I__9294 (
            .O(N__43894),
            .I(comm_buf_0_0));
    LocalMux I__9293 (
            .O(N__43891),
            .I(comm_buf_0_0));
    Odrv12 I__9292 (
            .O(N__43886),
            .I(comm_buf_0_0));
    InMux I__9291 (
            .O(N__43873),
            .I(N__43869));
    InMux I__9290 (
            .O(N__43872),
            .I(N__43866));
    LocalMux I__9289 (
            .O(N__43869),
            .I(N__43862));
    LocalMux I__9288 (
            .O(N__43866),
            .I(N__43859));
    InMux I__9287 (
            .O(N__43865),
            .I(N__43856));
    Span4Mux_v I__9286 (
            .O(N__43862),
            .I(N__43853));
    Span4Mux_h I__9285 (
            .O(N__43859),
            .I(N__43848));
    LocalMux I__9284 (
            .O(N__43856),
            .I(N__43848));
    Odrv4 I__9283 (
            .O(N__43853),
            .I(n11172));
    Odrv4 I__9282 (
            .O(N__43848),
            .I(n11172));
    InMux I__9281 (
            .O(N__43843),
            .I(N__43839));
    CascadeMux I__9280 (
            .O(N__43842),
            .I(N__43836));
    LocalMux I__9279 (
            .O(N__43839),
            .I(N__43832));
    InMux I__9278 (
            .O(N__43836),
            .I(N__43829));
    InMux I__9277 (
            .O(N__43835),
            .I(N__43825));
    Span4Mux_v I__9276 (
            .O(N__43832),
            .I(N__43822));
    LocalMux I__9275 (
            .O(N__43829),
            .I(N__43819));
    InMux I__9274 (
            .O(N__43828),
            .I(N__43815));
    LocalMux I__9273 (
            .O(N__43825),
            .I(N__43808));
    Sp12to4 I__9272 (
            .O(N__43822),
            .I(N__43808));
    Span12Mux_v I__9271 (
            .O(N__43819),
            .I(N__43808));
    InMux I__9270 (
            .O(N__43818),
            .I(N__43805));
    LocalMux I__9269 (
            .O(N__43815),
            .I(eis_start));
    Odrv12 I__9268 (
            .O(N__43808),
            .I(eis_start));
    LocalMux I__9267 (
            .O(N__43805),
            .I(eis_start));
    CascadeMux I__9266 (
            .O(N__43798),
            .I(n8_adj_1625_cascade_));
    CascadeMux I__9265 (
            .O(N__43795),
            .I(N__43792));
    CascadeBuf I__9264 (
            .O(N__43792),
            .I(N__43789));
    CascadeMux I__9263 (
            .O(N__43789),
            .I(N__43786));
    CascadeBuf I__9262 (
            .O(N__43786),
            .I(N__43783));
    CascadeMux I__9261 (
            .O(N__43783),
            .I(N__43780));
    CascadeBuf I__9260 (
            .O(N__43780),
            .I(N__43777));
    CascadeMux I__9259 (
            .O(N__43777),
            .I(N__43774));
    CascadeBuf I__9258 (
            .O(N__43774),
            .I(N__43771));
    CascadeMux I__9257 (
            .O(N__43771),
            .I(N__43768));
    CascadeBuf I__9256 (
            .O(N__43768),
            .I(N__43765));
    CascadeMux I__9255 (
            .O(N__43765),
            .I(N__43762));
    CascadeBuf I__9254 (
            .O(N__43762),
            .I(N__43759));
    CascadeMux I__9253 (
            .O(N__43759),
            .I(N__43755));
    CascadeMux I__9252 (
            .O(N__43758),
            .I(N__43752));
    CascadeBuf I__9251 (
            .O(N__43755),
            .I(N__43749));
    CascadeBuf I__9250 (
            .O(N__43752),
            .I(N__43746));
    CascadeMux I__9249 (
            .O(N__43749),
            .I(N__43743));
    CascadeMux I__9248 (
            .O(N__43746),
            .I(N__43740));
    CascadeBuf I__9247 (
            .O(N__43743),
            .I(N__43737));
    InMux I__9246 (
            .O(N__43740),
            .I(N__43734));
    CascadeMux I__9245 (
            .O(N__43737),
            .I(N__43731));
    LocalMux I__9244 (
            .O(N__43734),
            .I(N__43728));
    CascadeBuf I__9243 (
            .O(N__43731),
            .I(N__43725));
    Span4Mux_h I__9242 (
            .O(N__43728),
            .I(N__43722));
    CascadeMux I__9241 (
            .O(N__43725),
            .I(N__43719));
    Span4Mux_v I__9240 (
            .O(N__43722),
            .I(N__43716));
    InMux I__9239 (
            .O(N__43719),
            .I(N__43713));
    Span4Mux_v I__9238 (
            .O(N__43716),
            .I(N__43710));
    LocalMux I__9237 (
            .O(N__43713),
            .I(N__43707));
    Sp12to4 I__9236 (
            .O(N__43710),
            .I(N__43702));
    Span12Mux_s11_v I__9235 (
            .O(N__43707),
            .I(N__43702));
    Odrv12 I__9234 (
            .O(N__43702),
            .I(data_index_9_N_236_4));
    InMux I__9233 (
            .O(N__43699),
            .I(N__43696));
    LocalMux I__9232 (
            .O(N__43696),
            .I(N__43693));
    Span12Mux_h I__9231 (
            .O(N__43693),
            .I(N__43690));
    Odrv12 I__9230 (
            .O(N__43690),
            .I(n19_adj_1722));
    CascadeMux I__9229 (
            .O(N__43687),
            .I(N__43684));
    InMux I__9228 (
            .O(N__43684),
            .I(N__43681));
    LocalMux I__9227 (
            .O(N__43681),
            .I(N__43678));
    Span4Mux_v I__9226 (
            .O(N__43678),
            .I(N__43675));
    Span4Mux_v I__9225 (
            .O(N__43675),
            .I(N__43672));
    Sp12to4 I__9224 (
            .O(N__43672),
            .I(N__43668));
    InMux I__9223 (
            .O(N__43671),
            .I(N__43665));
    Odrv12 I__9222 (
            .O(N__43668),
            .I(buf_readRTD_6));
    LocalMux I__9221 (
            .O(N__43665),
            .I(buf_readRTD_6));
    InMux I__9220 (
            .O(N__43660),
            .I(N__43657));
    LocalMux I__9219 (
            .O(N__43657),
            .I(n23288));
    CascadeMux I__9218 (
            .O(N__43654),
            .I(n22396_cascade_));
    CascadeMux I__9217 (
            .O(N__43651),
            .I(N__43647));
    CascadeMux I__9216 (
            .O(N__43650),
            .I(N__43644));
    InMux I__9215 (
            .O(N__43647),
            .I(N__43641));
    InMux I__9214 (
            .O(N__43644),
            .I(N__43638));
    LocalMux I__9213 (
            .O(N__43641),
            .I(n6));
    LocalMux I__9212 (
            .O(N__43638),
            .I(n6));
    InMux I__9211 (
            .O(N__43633),
            .I(N__43629));
    InMux I__9210 (
            .O(N__43632),
            .I(N__43626));
    LocalMux I__9209 (
            .O(N__43629),
            .I(N__43623));
    LocalMux I__9208 (
            .O(N__43626),
            .I(n22061));
    Odrv4 I__9207 (
            .O(N__43623),
            .I(n22061));
    InMux I__9206 (
            .O(N__43618),
            .I(N__43613));
    InMux I__9205 (
            .O(N__43617),
            .I(N__43606));
    InMux I__9204 (
            .O(N__43616),
            .I(N__43606));
    LocalMux I__9203 (
            .O(N__43613),
            .I(N__43603));
    InMux I__9202 (
            .O(N__43612),
            .I(N__43600));
    InMux I__9201 (
            .O(N__43611),
            .I(N__43597));
    LocalMux I__9200 (
            .O(N__43606),
            .I(N__43592));
    Span4Mux_h I__9199 (
            .O(N__43603),
            .I(N__43592));
    LocalMux I__9198 (
            .O(N__43600),
            .I(N__43589));
    LocalMux I__9197 (
            .O(N__43597),
            .I(N__43586));
    Span4Mux_h I__9196 (
            .O(N__43592),
            .I(N__43583));
    Span4Mux_v I__9195 (
            .O(N__43589),
            .I(N__43578));
    Span4Mux_h I__9194 (
            .O(N__43586),
            .I(N__43578));
    Odrv4 I__9193 (
            .O(N__43583),
            .I(n21929));
    Odrv4 I__9192 (
            .O(N__43578),
            .I(n21929));
    InMux I__9191 (
            .O(N__43573),
            .I(N__43570));
    LocalMux I__9190 (
            .O(N__43570),
            .I(n22_adj_1801));
    InMux I__9189 (
            .O(N__43567),
            .I(N__43564));
    LocalMux I__9188 (
            .O(N__43564),
            .I(N__43561));
    Span4Mux_h I__9187 (
            .O(N__43561),
            .I(N__43558));
    Odrv4 I__9186 (
            .O(N__43558),
            .I(n112_adj_1799));
    InMux I__9185 (
            .O(N__43555),
            .I(N__43552));
    LocalMux I__9184 (
            .O(N__43552),
            .I(N__43549));
    Span4Mux_h I__9183 (
            .O(N__43549),
            .I(N__43546));
    Odrv4 I__9182 (
            .O(N__43546),
            .I(comm_buf_0_7_N_543_1));
    InMux I__9181 (
            .O(N__43543),
            .I(N__43540));
    LocalMux I__9180 (
            .O(N__43540),
            .I(N__43537));
    Span4Mux_v I__9179 (
            .O(N__43537),
            .I(N__43533));
    CascadeMux I__9178 (
            .O(N__43536),
            .I(N__43530));
    Span4Mux_h I__9177 (
            .O(N__43533),
            .I(N__43527));
    InMux I__9176 (
            .O(N__43530),
            .I(N__43524));
    Odrv4 I__9175 (
            .O(N__43527),
            .I(buf_adcdata_vdc_16));
    LocalMux I__9174 (
            .O(N__43524),
            .I(buf_adcdata_vdc_16));
    CascadeMux I__9173 (
            .O(N__43519),
            .I(n23504_cascade_));
    InMux I__9172 (
            .O(N__43516),
            .I(N__43513));
    LocalMux I__9171 (
            .O(N__43513),
            .I(N__43510));
    Span4Mux_h I__9170 (
            .O(N__43510),
            .I(N__43506));
    InMux I__9169 (
            .O(N__43509),
            .I(N__43503));
    Span4Mux_h I__9168 (
            .O(N__43506),
            .I(N__43500));
    LocalMux I__9167 (
            .O(N__43503),
            .I(N__43497));
    Span4Mux_h I__9166 (
            .O(N__43500),
            .I(N__43493));
    Span4Mux_h I__9165 (
            .O(N__43497),
            .I(N__43490));
    InMux I__9164 (
            .O(N__43496),
            .I(N__43487));
    Span4Mux_h I__9163 (
            .O(N__43493),
            .I(N__43484));
    Span4Mux_h I__9162 (
            .O(N__43490),
            .I(N__43481));
    LocalMux I__9161 (
            .O(N__43487),
            .I(buf_adcdata_vac_16));
    Odrv4 I__9160 (
            .O(N__43484),
            .I(buf_adcdata_vac_16));
    Odrv4 I__9159 (
            .O(N__43481),
            .I(buf_adcdata_vac_16));
    InMux I__9158 (
            .O(N__43474),
            .I(N__43471));
    LocalMux I__9157 (
            .O(N__43471),
            .I(N__43468));
    Span4Mux_v I__9156 (
            .O(N__43468),
            .I(N__43465));
    Odrv4 I__9155 (
            .O(N__43465),
            .I(n22288));
    CEMux I__9154 (
            .O(N__43462),
            .I(N__43459));
    LocalMux I__9153 (
            .O(N__43459),
            .I(N__43455));
    InMux I__9152 (
            .O(N__43458),
            .I(N__43452));
    Span4Mux_v I__9151 (
            .O(N__43455),
            .I(N__43447));
    LocalMux I__9150 (
            .O(N__43452),
            .I(N__43447));
    Odrv4 I__9149 (
            .O(N__43447),
            .I(n12838));
    InMux I__9148 (
            .O(N__43444),
            .I(N__43441));
    LocalMux I__9147 (
            .O(N__43441),
            .I(N__43438));
    Odrv12 I__9146 (
            .O(N__43438),
            .I(n23306));
    InMux I__9145 (
            .O(N__43435),
            .I(N__43432));
    LocalMux I__9144 (
            .O(N__43432),
            .I(N__43429));
    Odrv4 I__9143 (
            .O(N__43429),
            .I(n8_adj_1504));
    CascadeMux I__9142 (
            .O(N__43426),
            .I(n6_cascade_));
    InMux I__9141 (
            .O(N__43423),
            .I(N__43419));
    InMux I__9140 (
            .O(N__43422),
            .I(N__43416));
    LocalMux I__9139 (
            .O(N__43419),
            .I(N__43412));
    LocalMux I__9138 (
            .O(N__43416),
            .I(N__43409));
    InMux I__9137 (
            .O(N__43415),
            .I(N__43406));
    Span4Mux_h I__9136 (
            .O(N__43412),
            .I(N__43403));
    Span4Mux_v I__9135 (
            .O(N__43409),
            .I(N__43398));
    LocalMux I__9134 (
            .O(N__43406),
            .I(N__43398));
    Span4Mux_v I__9133 (
            .O(N__43403),
            .I(N__43395));
    Span4Mux_h I__9132 (
            .O(N__43398),
            .I(N__43392));
    Odrv4 I__9131 (
            .O(N__43395),
            .I(n21938));
    Odrv4 I__9130 (
            .O(N__43392),
            .I(n21938));
    InMux I__9129 (
            .O(N__43387),
            .I(N__43384));
    LocalMux I__9128 (
            .O(N__43384),
            .I(N__43381));
    Span4Mux_h I__9127 (
            .O(N__43381),
            .I(N__43378));
    Span4Mux_h I__9126 (
            .O(N__43378),
            .I(N__43375));
    Span4Mux_v I__9125 (
            .O(N__43375),
            .I(N__43372));
    Odrv4 I__9124 (
            .O(N__43372),
            .I(buf_data_vac_3));
    InMux I__9123 (
            .O(N__43369),
            .I(N__43366));
    LocalMux I__9122 (
            .O(N__43366),
            .I(N__43363));
    Span4Mux_v I__9121 (
            .O(N__43363),
            .I(N__43360));
    Span4Mux_h I__9120 (
            .O(N__43360),
            .I(N__43357));
    Odrv4 I__9119 (
            .O(N__43357),
            .I(buf_data_vac_2));
    InMux I__9118 (
            .O(N__43354),
            .I(N__43351));
    LocalMux I__9117 (
            .O(N__43351),
            .I(comm_buf_5_2));
    InMux I__9116 (
            .O(N__43348),
            .I(N__43345));
    LocalMux I__9115 (
            .O(N__43345),
            .I(N__43342));
    Span4Mux_v I__9114 (
            .O(N__43342),
            .I(N__43339));
    Span4Mux_h I__9113 (
            .O(N__43339),
            .I(N__43336));
    Odrv4 I__9112 (
            .O(N__43336),
            .I(buf_data_vac_1));
    InMux I__9111 (
            .O(N__43333),
            .I(N__43330));
    LocalMux I__9110 (
            .O(N__43330),
            .I(N__43327));
    Span4Mux_v I__9109 (
            .O(N__43327),
            .I(N__43324));
    Odrv4 I__9108 (
            .O(N__43324),
            .I(comm_buf_5_1));
    CascadeMux I__9107 (
            .O(N__43321),
            .I(N__43318));
    InMux I__9106 (
            .O(N__43318),
            .I(N__43315));
    LocalMux I__9105 (
            .O(N__43315),
            .I(N__43312));
    Span4Mux_v I__9104 (
            .O(N__43312),
            .I(N__43309));
    Span4Mux_h I__9103 (
            .O(N__43309),
            .I(N__43306));
    Span4Mux_h I__9102 (
            .O(N__43306),
            .I(N__43302));
    InMux I__9101 (
            .O(N__43305),
            .I(N__43299));
    Odrv4 I__9100 (
            .O(N__43302),
            .I(buf_readRTD_8));
    LocalMux I__9099 (
            .O(N__43299),
            .I(buf_readRTD_8));
    InMux I__9098 (
            .O(N__43294),
            .I(N__43291));
    LocalMux I__9097 (
            .O(N__43291),
            .I(N__43288));
    Odrv4 I__9096 (
            .O(N__43288),
            .I(n18816));
    InMux I__9095 (
            .O(N__43285),
            .I(N__43281));
    InMux I__9094 (
            .O(N__43284),
            .I(N__43278));
    LocalMux I__9093 (
            .O(N__43281),
            .I(N__43274));
    LocalMux I__9092 (
            .O(N__43278),
            .I(N__43271));
    InMux I__9091 (
            .O(N__43277),
            .I(N__43268));
    Span4Mux_h I__9090 (
            .O(N__43274),
            .I(N__43265));
    Span4Mux_h I__9089 (
            .O(N__43271),
            .I(N__43260));
    LocalMux I__9088 (
            .O(N__43268),
            .I(N__43260));
    Span4Mux_v I__9087 (
            .O(N__43265),
            .I(N__43257));
    Span4Mux_v I__9086 (
            .O(N__43260),
            .I(N__43254));
    Odrv4 I__9085 (
            .O(N__43257),
            .I(comm_tx_buf_0));
    Odrv4 I__9084 (
            .O(N__43254),
            .I(comm_tx_buf_0));
    InMux I__9083 (
            .O(N__43249),
            .I(N__43246));
    LocalMux I__9082 (
            .O(N__43246),
            .I(N__43243));
    Odrv4 I__9081 (
            .O(N__43243),
            .I(comm_buf_3_0));
    InMux I__9080 (
            .O(N__43240),
            .I(N__43237));
    LocalMux I__9079 (
            .O(N__43237),
            .I(n22338));
    InMux I__9078 (
            .O(N__43234),
            .I(N__43231));
    LocalMux I__9077 (
            .O(N__43231),
            .I(n18815));
    CascadeMux I__9076 (
            .O(N__43228),
            .I(N__43223));
    InMux I__9075 (
            .O(N__43227),
            .I(N__43220));
    InMux I__9074 (
            .O(N__43226),
            .I(N__43217));
    InMux I__9073 (
            .O(N__43223),
            .I(N__43214));
    LocalMux I__9072 (
            .O(N__43220),
            .I(N__43209));
    LocalMux I__9071 (
            .O(N__43217),
            .I(N__43209));
    LocalMux I__9070 (
            .O(N__43214),
            .I(N__43206));
    Span4Mux_v I__9069 (
            .O(N__43209),
            .I(N__43203));
    Odrv12 I__9068 (
            .O(N__43206),
            .I(comm_buf_2_0));
    Odrv4 I__9067 (
            .O(N__43203),
            .I(comm_buf_2_0));
    InMux I__9066 (
            .O(N__43198),
            .I(N__43195));
    LocalMux I__9065 (
            .O(N__43195),
            .I(N__43192));
    Span4Mux_h I__9064 (
            .O(N__43192),
            .I(N__43189));
    Odrv4 I__9063 (
            .O(N__43189),
            .I(n18823));
    InMux I__9062 (
            .O(N__43186),
            .I(N__43183));
    LocalMux I__9061 (
            .O(N__43183),
            .I(N__43180));
    Span4Mux_h I__9060 (
            .O(N__43180),
            .I(N__43177));
    Span4Mux_h I__9059 (
            .O(N__43177),
            .I(N__43174));
    Odrv4 I__9058 (
            .O(N__43174),
            .I(buf_data_vac_0));
    InMux I__9057 (
            .O(N__43171),
            .I(N__43168));
    LocalMux I__9056 (
            .O(N__43168),
            .I(comm_buf_5_0));
    InMux I__9055 (
            .O(N__43165),
            .I(N__43162));
    LocalMux I__9054 (
            .O(N__43162),
            .I(N__43159));
    Span4Mux_v I__9053 (
            .O(N__43159),
            .I(N__43156));
    Span4Mux_v I__9052 (
            .O(N__43156),
            .I(N__43153));
    Sp12to4 I__9051 (
            .O(N__43153),
            .I(N__43150));
    Odrv12 I__9050 (
            .O(N__43150),
            .I(buf_data_vac_7));
    InMux I__9049 (
            .O(N__43147),
            .I(N__43144));
    LocalMux I__9048 (
            .O(N__43144),
            .I(comm_buf_5_7));
    InMux I__9047 (
            .O(N__43141),
            .I(N__43138));
    LocalMux I__9046 (
            .O(N__43138),
            .I(N__43135));
    Span4Mux_v I__9045 (
            .O(N__43135),
            .I(N__43132));
    Sp12to4 I__9044 (
            .O(N__43132),
            .I(N__43129));
    Odrv12 I__9043 (
            .O(N__43129),
            .I(buf_data_vac_6));
    InMux I__9042 (
            .O(N__43126),
            .I(N__43123));
    LocalMux I__9041 (
            .O(N__43123),
            .I(N__43120));
    Span4Mux_h I__9040 (
            .O(N__43120),
            .I(N__43117));
    Odrv4 I__9039 (
            .O(N__43117),
            .I(comm_buf_5_6));
    InMux I__9038 (
            .O(N__43114),
            .I(N__43111));
    LocalMux I__9037 (
            .O(N__43111),
            .I(N__43108));
    Span4Mux_v I__9036 (
            .O(N__43108),
            .I(N__43105));
    Sp12to4 I__9035 (
            .O(N__43105),
            .I(N__43102));
    Odrv12 I__9034 (
            .O(N__43102),
            .I(buf_data_vac_5));
    InMux I__9033 (
            .O(N__43099),
            .I(N__43096));
    LocalMux I__9032 (
            .O(N__43096),
            .I(N__43093));
    Span4Mux_v I__9031 (
            .O(N__43093),
            .I(N__43090));
    Sp12to4 I__9030 (
            .O(N__43090),
            .I(N__43087));
    Odrv12 I__9029 (
            .O(N__43087),
            .I(buf_data_vac_4));
    InMux I__9028 (
            .O(N__43084),
            .I(N__43081));
    LocalMux I__9027 (
            .O(N__43081),
            .I(N__43078));
    Span4Mux_h I__9026 (
            .O(N__43078),
            .I(N__43075));
    Odrv4 I__9025 (
            .O(N__43075),
            .I(comm_buf_5_4));
    InMux I__9024 (
            .O(N__43072),
            .I(N__43068));
    InMux I__9023 (
            .O(N__43071),
            .I(N__43065));
    LocalMux I__9022 (
            .O(N__43068),
            .I(comm_buf_6_7));
    LocalMux I__9021 (
            .O(N__43065),
            .I(comm_buf_6_7));
    InMux I__9020 (
            .O(N__43060),
            .I(N__43057));
    LocalMux I__9019 (
            .O(N__43057),
            .I(N__43053));
    InMux I__9018 (
            .O(N__43056),
            .I(N__43050));
    Span4Mux_h I__9017 (
            .O(N__43053),
            .I(N__43047));
    LocalMux I__9016 (
            .O(N__43050),
            .I(comm_test_buf_24_17));
    Odrv4 I__9015 (
            .O(N__43047),
            .I(comm_test_buf_24_17));
    CascadeMux I__9014 (
            .O(N__43042),
            .I(N__43038));
    InMux I__9013 (
            .O(N__43041),
            .I(N__43035));
    InMux I__9012 (
            .O(N__43038),
            .I(N__43032));
    LocalMux I__9011 (
            .O(N__43035),
            .I(N__43029));
    LocalMux I__9010 (
            .O(N__43032),
            .I(comm_buf_6_0));
    Odrv12 I__9009 (
            .O(N__43029),
            .I(comm_buf_6_0));
    CascadeMux I__9008 (
            .O(N__43024),
            .I(n18818_cascade_));
    CascadeMux I__9007 (
            .O(N__43021),
            .I(n23372_cascade_));
    InMux I__9006 (
            .O(N__43018),
            .I(N__43014));
    InMux I__9005 (
            .O(N__43017),
            .I(N__43011));
    LocalMux I__9004 (
            .O(N__43014),
            .I(secclk_cnt_20));
    LocalMux I__9003 (
            .O(N__43011),
            .I(secclk_cnt_20));
    CascadeMux I__9002 (
            .O(N__43006),
            .I(n20922_cascade_));
    InMux I__9001 (
            .O(N__43003),
            .I(N__43000));
    LocalMux I__9000 (
            .O(N__43000),
            .I(N__42997));
    Odrv4 I__8999 (
            .O(N__42997),
            .I(n14_adj_1678));
    InMux I__8998 (
            .O(N__42994),
            .I(N__42990));
    InMux I__8997 (
            .O(N__42993),
            .I(N__42987));
    LocalMux I__8996 (
            .O(N__42990),
            .I(secclk_cnt_9));
    LocalMux I__8995 (
            .O(N__42987),
            .I(secclk_cnt_9));
    InMux I__8994 (
            .O(N__42982),
            .I(N__42978));
    InMux I__8993 (
            .O(N__42981),
            .I(N__42975));
    LocalMux I__8992 (
            .O(N__42978),
            .I(N__42972));
    LocalMux I__8991 (
            .O(N__42975),
            .I(secclk_cnt_17));
    Odrv4 I__8990 (
            .O(N__42972),
            .I(secclk_cnt_17));
    InMux I__8989 (
            .O(N__42967),
            .I(N__42964));
    LocalMux I__8988 (
            .O(N__42964),
            .I(n10_adj_1679));
    InMux I__8987 (
            .O(N__42961),
            .I(N__42957));
    InMux I__8986 (
            .O(N__42960),
            .I(N__42954));
    LocalMux I__8985 (
            .O(N__42957),
            .I(secclk_cnt_6));
    LocalMux I__8984 (
            .O(N__42954),
            .I(secclk_cnt_6));
    InMux I__8983 (
            .O(N__42949),
            .I(N__42945));
    InMux I__8982 (
            .O(N__42948),
            .I(N__42942));
    LocalMux I__8981 (
            .O(N__42945),
            .I(secclk_cnt_14));
    LocalMux I__8980 (
            .O(N__42942),
            .I(secclk_cnt_14));
    CascadeMux I__8979 (
            .O(N__42937),
            .I(N__42933));
    InMux I__8978 (
            .O(N__42936),
            .I(N__42930));
    InMux I__8977 (
            .O(N__42933),
            .I(N__42927));
    LocalMux I__8976 (
            .O(N__42930),
            .I(secclk_cnt_10));
    LocalMux I__8975 (
            .O(N__42927),
            .I(secclk_cnt_10));
    InMux I__8974 (
            .O(N__42922),
            .I(N__42918));
    InMux I__8973 (
            .O(N__42921),
            .I(N__42915));
    LocalMux I__8972 (
            .O(N__42918),
            .I(secclk_cnt_3));
    LocalMux I__8971 (
            .O(N__42915),
            .I(secclk_cnt_3));
    InMux I__8970 (
            .O(N__42910),
            .I(N__42907));
    LocalMux I__8969 (
            .O(N__42907),
            .I(n27));
    InMux I__8968 (
            .O(N__42904),
            .I(N__42900));
    InMux I__8967 (
            .O(N__42903),
            .I(N__42897));
    LocalMux I__8966 (
            .O(N__42900),
            .I(secclk_cnt_16));
    LocalMux I__8965 (
            .O(N__42897),
            .I(secclk_cnt_16));
    InMux I__8964 (
            .O(N__42892),
            .I(N__42888));
    InMux I__8963 (
            .O(N__42891),
            .I(N__42885));
    LocalMux I__8962 (
            .O(N__42888),
            .I(secclk_cnt_7));
    LocalMux I__8961 (
            .O(N__42885),
            .I(secclk_cnt_7));
    CascadeMux I__8960 (
            .O(N__42880),
            .I(N__42876));
    InMux I__8959 (
            .O(N__42879),
            .I(N__42873));
    InMux I__8958 (
            .O(N__42876),
            .I(N__42870));
    LocalMux I__8957 (
            .O(N__42873),
            .I(secclk_cnt_13));
    LocalMux I__8956 (
            .O(N__42870),
            .I(secclk_cnt_13));
    InMux I__8955 (
            .O(N__42865),
            .I(N__42861));
    InMux I__8954 (
            .O(N__42864),
            .I(N__42858));
    LocalMux I__8953 (
            .O(N__42861),
            .I(secclk_cnt_2));
    LocalMux I__8952 (
            .O(N__42858),
            .I(secclk_cnt_2));
    InMux I__8951 (
            .O(N__42853),
            .I(N__42850));
    LocalMux I__8950 (
            .O(N__42850),
            .I(n26_adj_1715));
    SRMux I__8949 (
            .O(N__42847),
            .I(N__42842));
    SRMux I__8948 (
            .O(N__42846),
            .I(N__42839));
    SRMux I__8947 (
            .O(N__42845),
            .I(N__42836));
    LocalMux I__8946 (
            .O(N__42842),
            .I(N__42833));
    LocalMux I__8945 (
            .O(N__42839),
            .I(N__42830));
    LocalMux I__8944 (
            .O(N__42836),
            .I(N__42827));
    Span4Mux_v I__8943 (
            .O(N__42833),
            .I(N__42821));
    Span4Mux_v I__8942 (
            .O(N__42830),
            .I(N__42821));
    Span4Mux_h I__8941 (
            .O(N__42827),
            .I(N__42818));
    InMux I__8940 (
            .O(N__42826),
            .I(N__42815));
    Odrv4 I__8939 (
            .O(N__42821),
            .I(n15420));
    Odrv4 I__8938 (
            .O(N__42818),
            .I(n15420));
    LocalMux I__8937 (
            .O(N__42815),
            .I(n15420));
    IoInMux I__8936 (
            .O(N__42808),
            .I(N__42805));
    LocalMux I__8935 (
            .O(N__42805),
            .I(N__42802));
    Span4Mux_s2_v I__8934 (
            .O(N__42802),
            .I(N__42799));
    Span4Mux_h I__8933 (
            .O(N__42799),
            .I(N__42796));
    Sp12to4 I__8932 (
            .O(N__42796),
            .I(N__42793));
    Span12Mux_h I__8931 (
            .O(N__42793),
            .I(N__42789));
    InMux I__8930 (
            .O(N__42792),
            .I(N__42786));
    Odrv12 I__8929 (
            .O(N__42789),
            .I(TEST_LED));
    LocalMux I__8928 (
            .O(N__42786),
            .I(TEST_LED));
    CascadeMux I__8927 (
            .O(N__42781),
            .I(N__42778));
    InMux I__8926 (
            .O(N__42778),
            .I(N__42775));
    LocalMux I__8925 (
            .O(N__42775),
            .I(N__42772));
    Span4Mux_h I__8924 (
            .O(N__42772),
            .I(N__42769));
    Odrv4 I__8923 (
            .O(N__42769),
            .I(n9_adj_1596));
    InMux I__8922 (
            .O(N__42766),
            .I(N__42763));
    LocalMux I__8921 (
            .O(N__42763),
            .I(\comm_spi.n15327 ));
    IoInMux I__8920 (
            .O(N__42760),
            .I(N__42754));
    ClkMux I__8919 (
            .O(N__42759),
            .I(N__42750));
    ClkMux I__8918 (
            .O(N__42758),
            .I(N__42744));
    ClkMux I__8917 (
            .O(N__42757),
            .I(N__42741));
    LocalMux I__8916 (
            .O(N__42754),
            .I(N__42734));
    ClkMux I__8915 (
            .O(N__42753),
            .I(N__42731));
    LocalMux I__8914 (
            .O(N__42750),
            .I(N__42728));
    ClkMux I__8913 (
            .O(N__42749),
            .I(N__42725));
    ClkMux I__8912 (
            .O(N__42748),
            .I(N__42722));
    ClkMux I__8911 (
            .O(N__42747),
            .I(N__42714));
    LocalMux I__8910 (
            .O(N__42744),
            .I(N__42711));
    LocalMux I__8909 (
            .O(N__42741),
            .I(N__42708));
    ClkMux I__8908 (
            .O(N__42740),
            .I(N__42705));
    ClkMux I__8907 (
            .O(N__42739),
            .I(N__42702));
    ClkMux I__8906 (
            .O(N__42738),
            .I(N__42699));
    ClkMux I__8905 (
            .O(N__42737),
            .I(N__42691));
    IoSpan4Mux I__8904 (
            .O(N__42734),
            .I(N__42687));
    LocalMux I__8903 (
            .O(N__42731),
            .I(N__42684));
    Span4Mux_v I__8902 (
            .O(N__42728),
            .I(N__42679));
    LocalMux I__8901 (
            .O(N__42725),
            .I(N__42679));
    LocalMux I__8900 (
            .O(N__42722),
            .I(N__42676));
    ClkMux I__8899 (
            .O(N__42721),
            .I(N__42673));
    ClkMux I__8898 (
            .O(N__42720),
            .I(N__42670));
    ClkMux I__8897 (
            .O(N__42719),
            .I(N__42667));
    ClkMux I__8896 (
            .O(N__42718),
            .I(N__42664));
    ClkMux I__8895 (
            .O(N__42717),
            .I(N__42660));
    LocalMux I__8894 (
            .O(N__42714),
            .I(N__42657));
    Span4Mux_v I__8893 (
            .O(N__42711),
            .I(N__42646));
    Span4Mux_h I__8892 (
            .O(N__42708),
            .I(N__42646));
    LocalMux I__8891 (
            .O(N__42705),
            .I(N__42646));
    LocalMux I__8890 (
            .O(N__42702),
            .I(N__42646));
    LocalMux I__8889 (
            .O(N__42699),
            .I(N__42646));
    ClkMux I__8888 (
            .O(N__42698),
            .I(N__42643));
    ClkMux I__8887 (
            .O(N__42697),
            .I(N__42640));
    ClkMux I__8886 (
            .O(N__42696),
            .I(N__42637));
    ClkMux I__8885 (
            .O(N__42695),
            .I(N__42634));
    ClkMux I__8884 (
            .O(N__42694),
            .I(N__42631));
    LocalMux I__8883 (
            .O(N__42691),
            .I(N__42628));
    ClkMux I__8882 (
            .O(N__42690),
            .I(N__42625));
    Sp12to4 I__8881 (
            .O(N__42687),
            .I(N__42622));
    Span4Mux_v I__8880 (
            .O(N__42684),
            .I(N__42617));
    Span4Mux_v I__8879 (
            .O(N__42679),
            .I(N__42617));
    Span4Mux_v I__8878 (
            .O(N__42676),
            .I(N__42606));
    LocalMux I__8877 (
            .O(N__42673),
            .I(N__42606));
    LocalMux I__8876 (
            .O(N__42670),
            .I(N__42606));
    LocalMux I__8875 (
            .O(N__42667),
            .I(N__42606));
    LocalMux I__8874 (
            .O(N__42664),
            .I(N__42606));
    ClkMux I__8873 (
            .O(N__42663),
            .I(N__42603));
    LocalMux I__8872 (
            .O(N__42660),
            .I(N__42600));
    Span4Mux_v I__8871 (
            .O(N__42657),
            .I(N__42593));
    Span4Mux_v I__8870 (
            .O(N__42646),
            .I(N__42593));
    LocalMux I__8869 (
            .O(N__42643),
            .I(N__42593));
    LocalMux I__8868 (
            .O(N__42640),
            .I(N__42590));
    LocalMux I__8867 (
            .O(N__42637),
            .I(N__42587));
    LocalMux I__8866 (
            .O(N__42634),
            .I(N__42584));
    LocalMux I__8865 (
            .O(N__42631),
            .I(N__42581));
    Span4Mux_h I__8864 (
            .O(N__42628),
            .I(N__42576));
    LocalMux I__8863 (
            .O(N__42625),
            .I(N__42576));
    Span12Mux_s6_h I__8862 (
            .O(N__42622),
            .I(N__42573));
    Span4Mux_h I__8861 (
            .O(N__42617),
            .I(N__42570));
    Span4Mux_v I__8860 (
            .O(N__42606),
            .I(N__42565));
    LocalMux I__8859 (
            .O(N__42603),
            .I(N__42565));
    Span4Mux_h I__8858 (
            .O(N__42600),
            .I(N__42560));
    Span4Mux_h I__8857 (
            .O(N__42593),
            .I(N__42560));
    Span4Mux_v I__8856 (
            .O(N__42590),
            .I(N__42555));
    Span4Mux_h I__8855 (
            .O(N__42587),
            .I(N__42555));
    Span4Mux_v I__8854 (
            .O(N__42584),
            .I(N__42548));
    Span4Mux_h I__8853 (
            .O(N__42581),
            .I(N__42548));
    Span4Mux_v I__8852 (
            .O(N__42576),
            .I(N__42548));
    Span12Mux_h I__8851 (
            .O(N__42573),
            .I(N__42543));
    Sp12to4 I__8850 (
            .O(N__42570),
            .I(N__42543));
    Span4Mux_h I__8849 (
            .O(N__42565),
            .I(N__42540));
    Span4Mux_h I__8848 (
            .O(N__42560),
            .I(N__42537));
    Span4Mux_h I__8847 (
            .O(N__42555),
            .I(N__42534));
    Span4Mux_h I__8846 (
            .O(N__42548),
            .I(N__42531));
    Odrv12 I__8845 (
            .O(N__42543),
            .I(VDC_CLK));
    Odrv4 I__8844 (
            .O(N__42540),
            .I(VDC_CLK));
    Odrv4 I__8843 (
            .O(N__42537),
            .I(VDC_CLK));
    Odrv4 I__8842 (
            .O(N__42534),
            .I(VDC_CLK));
    Odrv4 I__8841 (
            .O(N__42531),
            .I(VDC_CLK));
    InMux I__8840 (
            .O(N__42520),
            .I(N__42517));
    LocalMux I__8839 (
            .O(N__42517),
            .I(N__42514));
    Odrv4 I__8838 (
            .O(N__42514),
            .I(n4_adj_1676));
    SRMux I__8837 (
            .O(N__42511),
            .I(N__42508));
    LocalMux I__8836 (
            .O(N__42508),
            .I(N__42505));
    Span4Mux_v I__8835 (
            .O(N__42505),
            .I(N__42502));
    Odrv4 I__8834 (
            .O(N__42502),
            .I(\comm_spi.DOUT_7__N_835 ));
    InMux I__8833 (
            .O(N__42499),
            .I(N__42495));
    InMux I__8832 (
            .O(N__42498),
            .I(N__42492));
    LocalMux I__8831 (
            .O(N__42495),
            .I(N__42484));
    LocalMux I__8830 (
            .O(N__42492),
            .I(N__42484));
    InMux I__8829 (
            .O(N__42491),
            .I(N__42481));
    InMux I__8828 (
            .O(N__42490),
            .I(N__42478));
    InMux I__8827 (
            .O(N__42489),
            .I(N__42475));
    Span4Mux_v I__8826 (
            .O(N__42484),
            .I(N__42472));
    LocalMux I__8825 (
            .O(N__42481),
            .I(N__42469));
    LocalMux I__8824 (
            .O(N__42478),
            .I(N__42466));
    LocalMux I__8823 (
            .O(N__42475),
            .I(N__42463));
    Span4Mux_v I__8822 (
            .O(N__42472),
            .I(N__42460));
    Sp12to4 I__8821 (
            .O(N__42469),
            .I(N__42453));
    Sp12to4 I__8820 (
            .O(N__42466),
            .I(N__42453));
    Sp12to4 I__8819 (
            .O(N__42463),
            .I(N__42453));
    Sp12to4 I__8818 (
            .O(N__42460),
            .I(N__42448));
    Span12Mux_v I__8817 (
            .O(N__42453),
            .I(N__42448));
    Span12Mux_h I__8816 (
            .O(N__42448),
            .I(N__42445));
    Odrv12 I__8815 (
            .O(N__42445),
            .I(ICE_SPI_SCLK));
    SRMux I__8814 (
            .O(N__42442),
            .I(N__42439));
    LocalMux I__8813 (
            .O(N__42439),
            .I(N__42436));
    Span4Mux_h I__8812 (
            .O(N__42436),
            .I(N__42433));
    Odrv4 I__8811 (
            .O(N__42433),
            .I(\comm_spi.iclk_N_851 ));
    InMux I__8810 (
            .O(N__42430),
            .I(N__42426));
    InMux I__8809 (
            .O(N__42429),
            .I(N__42423));
    LocalMux I__8808 (
            .O(N__42426),
            .I(secclk_cnt_15));
    LocalMux I__8807 (
            .O(N__42423),
            .I(secclk_cnt_15));
    InMux I__8806 (
            .O(N__42418),
            .I(N__42414));
    InMux I__8805 (
            .O(N__42417),
            .I(N__42411));
    LocalMux I__8804 (
            .O(N__42414),
            .I(secclk_cnt_8));
    LocalMux I__8803 (
            .O(N__42411),
            .I(secclk_cnt_8));
    CascadeMux I__8802 (
            .O(N__42406),
            .I(N__42402));
    InMux I__8801 (
            .O(N__42405),
            .I(N__42399));
    InMux I__8800 (
            .O(N__42402),
            .I(N__42396));
    LocalMux I__8799 (
            .O(N__42399),
            .I(secclk_cnt_1));
    LocalMux I__8798 (
            .O(N__42396),
            .I(secclk_cnt_1));
    InMux I__8797 (
            .O(N__42391),
            .I(N__42387));
    InMux I__8796 (
            .O(N__42390),
            .I(N__42384));
    LocalMux I__8795 (
            .O(N__42387),
            .I(secclk_cnt_5));
    LocalMux I__8794 (
            .O(N__42384),
            .I(secclk_cnt_5));
    CascadeMux I__8793 (
            .O(N__42379),
            .I(n25_adj_1717_cascade_));
    InMux I__8792 (
            .O(N__42376),
            .I(N__42373));
    LocalMux I__8791 (
            .O(N__42373),
            .I(N__42369));
    InMux I__8790 (
            .O(N__42372),
            .I(N__42366));
    Span4Mux_h I__8789 (
            .O(N__42369),
            .I(N__42363));
    LocalMux I__8788 (
            .O(N__42366),
            .I(comm_test_buf_24_23));
    Odrv4 I__8787 (
            .O(N__42363),
            .I(comm_test_buf_24_23));
    InMux I__8786 (
            .O(N__42358),
            .I(N__42355));
    LocalMux I__8785 (
            .O(N__42355),
            .I(N__42352));
    Span4Mux_v I__8784 (
            .O(N__42352),
            .I(N__42347));
    InMux I__8783 (
            .O(N__42351),
            .I(N__42344));
    InMux I__8782 (
            .O(N__42350),
            .I(N__42341));
    Odrv4 I__8781 (
            .O(N__42347),
            .I(buf_dds0_2));
    LocalMux I__8780 (
            .O(N__42344),
            .I(buf_dds0_2));
    LocalMux I__8779 (
            .O(N__42341),
            .I(buf_dds0_2));
    InMux I__8778 (
            .O(N__42334),
            .I(N__42329));
    InMux I__8777 (
            .O(N__42333),
            .I(N__42326));
    InMux I__8776 (
            .O(N__42332),
            .I(N__42323));
    LocalMux I__8775 (
            .O(N__42329),
            .I(N__42320));
    LocalMux I__8774 (
            .O(N__42326),
            .I(N__42317));
    LocalMux I__8773 (
            .O(N__42323),
            .I(N__42314));
    Span4Mux_h I__8772 (
            .O(N__42320),
            .I(N__42311));
    Span4Mux_v I__8771 (
            .O(N__42317),
            .I(N__42306));
    Span4Mux_v I__8770 (
            .O(N__42314),
            .I(N__42306));
    Odrv4 I__8769 (
            .O(N__42311),
            .I(data_index_9));
    Odrv4 I__8768 (
            .O(N__42306),
            .I(data_index_9));
    CascadeMux I__8767 (
            .O(N__42301),
            .I(n8_adj_1617_cascade_));
    CascadeMux I__8766 (
            .O(N__42298),
            .I(N__42295));
    CascadeBuf I__8765 (
            .O(N__42295),
            .I(N__42292));
    CascadeMux I__8764 (
            .O(N__42292),
            .I(N__42289));
    CascadeBuf I__8763 (
            .O(N__42289),
            .I(N__42286));
    CascadeMux I__8762 (
            .O(N__42286),
            .I(N__42283));
    CascadeBuf I__8761 (
            .O(N__42283),
            .I(N__42280));
    CascadeMux I__8760 (
            .O(N__42280),
            .I(N__42277));
    CascadeBuf I__8759 (
            .O(N__42277),
            .I(N__42274));
    CascadeMux I__8758 (
            .O(N__42274),
            .I(N__42271));
    CascadeBuf I__8757 (
            .O(N__42271),
            .I(N__42268));
    CascadeMux I__8756 (
            .O(N__42268),
            .I(N__42265));
    CascadeBuf I__8755 (
            .O(N__42265),
            .I(N__42262));
    CascadeMux I__8754 (
            .O(N__42262),
            .I(N__42259));
    CascadeBuf I__8753 (
            .O(N__42259),
            .I(N__42255));
    CascadeMux I__8752 (
            .O(N__42258),
            .I(N__42252));
    CascadeMux I__8751 (
            .O(N__42255),
            .I(N__42249));
    CascadeBuf I__8750 (
            .O(N__42252),
            .I(N__42246));
    CascadeBuf I__8749 (
            .O(N__42249),
            .I(N__42243));
    CascadeMux I__8748 (
            .O(N__42246),
            .I(N__42240));
    CascadeMux I__8747 (
            .O(N__42243),
            .I(N__42237));
    InMux I__8746 (
            .O(N__42240),
            .I(N__42234));
    CascadeBuf I__8745 (
            .O(N__42237),
            .I(N__42231));
    LocalMux I__8744 (
            .O(N__42234),
            .I(N__42228));
    CascadeMux I__8743 (
            .O(N__42231),
            .I(N__42225));
    Span12Mux_h I__8742 (
            .O(N__42228),
            .I(N__42222));
    InMux I__8741 (
            .O(N__42225),
            .I(N__42219));
    Span12Mux_v I__8740 (
            .O(N__42222),
            .I(N__42216));
    LocalMux I__8739 (
            .O(N__42219),
            .I(N__42213));
    Odrv12 I__8738 (
            .O(N__42216),
            .I(data_index_9_N_236_8));
    Odrv12 I__8737 (
            .O(N__42213),
            .I(data_index_9_N_236_8));
    CEMux I__8736 (
            .O(N__42208),
            .I(N__42202));
    CEMux I__8735 (
            .O(N__42207),
            .I(N__42199));
    CEMux I__8734 (
            .O(N__42206),
            .I(N__42196));
    CEMux I__8733 (
            .O(N__42205),
            .I(N__42193));
    LocalMux I__8732 (
            .O(N__42202),
            .I(N__42190));
    LocalMux I__8731 (
            .O(N__42199),
            .I(N__42187));
    LocalMux I__8730 (
            .O(N__42196),
            .I(N__42182));
    LocalMux I__8729 (
            .O(N__42193),
            .I(N__42182));
    Span4Mux_v I__8728 (
            .O(N__42190),
            .I(N__42179));
    Span4Mux_h I__8727 (
            .O(N__42187),
            .I(N__42176));
    Span4Mux_h I__8726 (
            .O(N__42182),
            .I(N__42173));
    Odrv4 I__8725 (
            .O(N__42179),
            .I(\SIG_DDS.n13338 ));
    Odrv4 I__8724 (
            .O(N__42176),
            .I(\SIG_DDS.n13338 ));
    Odrv4 I__8723 (
            .O(N__42173),
            .I(\SIG_DDS.n13338 ));
    SRMux I__8722 (
            .O(N__42166),
            .I(N__42163));
    LocalMux I__8721 (
            .O(N__42163),
            .I(N__42160));
    Span4Mux_h I__8720 (
            .O(N__42160),
            .I(N__42157));
    Odrv4 I__8719 (
            .O(N__42157),
            .I(\comm_spi.iclk_N_850 ));
    InMux I__8718 (
            .O(N__42154),
            .I(N__42149));
    InMux I__8717 (
            .O(N__42153),
            .I(N__42146));
    InMux I__8716 (
            .O(N__42152),
            .I(N__42143));
    LocalMux I__8715 (
            .O(N__42149),
            .I(N__42140));
    LocalMux I__8714 (
            .O(N__42146),
            .I(buf_dds0_1));
    LocalMux I__8713 (
            .O(N__42143),
            .I(buf_dds0_1));
    Odrv4 I__8712 (
            .O(N__42140),
            .I(buf_dds0_1));
    InMux I__8711 (
            .O(N__42133),
            .I(N__42129));
    InMux I__8710 (
            .O(N__42132),
            .I(N__42126));
    LocalMux I__8709 (
            .O(N__42129),
            .I(N__42122));
    LocalMux I__8708 (
            .O(N__42126),
            .I(N__42119));
    InMux I__8707 (
            .O(N__42125),
            .I(N__42116));
    Span4Mux_h I__8706 (
            .O(N__42122),
            .I(N__42113));
    Span12Mux_s11_v I__8705 (
            .O(N__42119),
            .I(N__42110));
    LocalMux I__8704 (
            .O(N__42116),
            .I(buf_dds1_1));
    Odrv4 I__8703 (
            .O(N__42113),
            .I(buf_dds1_1));
    Odrv12 I__8702 (
            .O(N__42110),
            .I(buf_dds1_1));
    InMux I__8701 (
            .O(N__42103),
            .I(N__42100));
    LocalMux I__8700 (
            .O(N__42100),
            .I(N__42097));
    Span4Mux_h I__8699 (
            .O(N__42097),
            .I(N__42092));
    InMux I__8698 (
            .O(N__42096),
            .I(N__42089));
    InMux I__8697 (
            .O(N__42095),
            .I(N__42086));
    Span4Mux_h I__8696 (
            .O(N__42092),
            .I(N__42083));
    LocalMux I__8695 (
            .O(N__42089),
            .I(buf_dds1_2));
    LocalMux I__8694 (
            .O(N__42086),
            .I(buf_dds1_2));
    Odrv4 I__8693 (
            .O(N__42083),
            .I(buf_dds1_2));
    InMux I__8692 (
            .O(N__42076),
            .I(N__42073));
    LocalMux I__8691 (
            .O(N__42073),
            .I(N__42070));
    Span4Mux_v I__8690 (
            .O(N__42070),
            .I(N__42066));
    InMux I__8689 (
            .O(N__42069),
            .I(N__42063));
    Span4Mux_h I__8688 (
            .O(N__42066),
            .I(N__42060));
    LocalMux I__8687 (
            .O(N__42063),
            .I(N__42057));
    Span4Mux_h I__8686 (
            .O(N__42060),
            .I(N__42053));
    Span4Mux_h I__8685 (
            .O(N__42057),
            .I(N__42050));
    InMux I__8684 (
            .O(N__42056),
            .I(N__42047));
    Span4Mux_h I__8683 (
            .O(N__42053),
            .I(N__42044));
    Span4Mux_v I__8682 (
            .O(N__42050),
            .I(N__42041));
    LocalMux I__8681 (
            .O(N__42047),
            .I(buf_adcdata_iac_10));
    Odrv4 I__8680 (
            .O(N__42044),
            .I(buf_adcdata_iac_10));
    Odrv4 I__8679 (
            .O(N__42041),
            .I(buf_adcdata_iac_10));
    CascadeMux I__8678 (
            .O(N__42034),
            .I(n16_adj_1746_cascade_));
    InMux I__8677 (
            .O(N__42031),
            .I(N__42028));
    LocalMux I__8676 (
            .O(N__42028),
            .I(N__42025));
    Span4Mux_h I__8675 (
            .O(N__42025),
            .I(N__42022));
    Sp12to4 I__8674 (
            .O(N__42022),
            .I(N__42018));
    InMux I__8673 (
            .O(N__42021),
            .I(N__42015));
    Span12Mux_v I__8672 (
            .O(N__42018),
            .I(N__42010));
    LocalMux I__8671 (
            .O(N__42015),
            .I(N__42010));
    Odrv12 I__8670 (
            .O(N__42010),
            .I(\comm_spi.n15341 ));
    InMux I__8669 (
            .O(N__42007),
            .I(N__42004));
    LocalMux I__8668 (
            .O(N__42004),
            .I(N__42000));
    InMux I__8667 (
            .O(N__42003),
            .I(N__41997));
    Span4Mux_v I__8666 (
            .O(N__42000),
            .I(N__41994));
    LocalMux I__8665 (
            .O(N__41997),
            .I(N__41991));
    Odrv4 I__8664 (
            .O(N__41994),
            .I(\comm_spi.n15340 ));
    Odrv12 I__8663 (
            .O(N__41991),
            .I(\comm_spi.n15340 ));
    InMux I__8662 (
            .O(N__41986),
            .I(N__41982));
    InMux I__8661 (
            .O(N__41985),
            .I(N__41977));
    LocalMux I__8660 (
            .O(N__41982),
            .I(N__41974));
    InMux I__8659 (
            .O(N__41981),
            .I(N__41971));
    InMux I__8658 (
            .O(N__41980),
            .I(N__41967));
    LocalMux I__8657 (
            .O(N__41977),
            .I(N__41964));
    Span4Mux_v I__8656 (
            .O(N__41974),
            .I(N__41958));
    LocalMux I__8655 (
            .O(N__41971),
            .I(N__41958));
    InMux I__8654 (
            .O(N__41970),
            .I(N__41955));
    LocalMux I__8653 (
            .O(N__41967),
            .I(N__41950));
    Span4Mux_v I__8652 (
            .O(N__41964),
            .I(N__41950));
    InMux I__8651 (
            .O(N__41963),
            .I(N__41947));
    Span4Mux_h I__8650 (
            .O(N__41958),
            .I(N__41940));
    LocalMux I__8649 (
            .O(N__41955),
            .I(N__41940));
    Span4Mux_v I__8648 (
            .O(N__41950),
            .I(N__41940));
    LocalMux I__8647 (
            .O(N__41947),
            .I(\comm_spi.n15333 ));
    Odrv4 I__8646 (
            .O(N__41940),
            .I(\comm_spi.n15333 ));
    InMux I__8645 (
            .O(N__41935),
            .I(N__41932));
    LocalMux I__8644 (
            .O(N__41932),
            .I(N__41929));
    Span4Mux_v I__8643 (
            .O(N__41929),
            .I(N__41926));
    Span4Mux_h I__8642 (
            .O(N__41926),
            .I(N__41923));
    Sp12to4 I__8641 (
            .O(N__41923),
            .I(N__41920));
    Span12Mux_h I__8640 (
            .O(N__41920),
            .I(N__41917));
    Odrv12 I__8639 (
            .O(N__41917),
            .I(\comm_spi.n15334 ));
    SRMux I__8638 (
            .O(N__41914),
            .I(N__41910));
    SRMux I__8637 (
            .O(N__41913),
            .I(N__41907));
    LocalMux I__8636 (
            .O(N__41910),
            .I(N__41904));
    LocalMux I__8635 (
            .O(N__41907),
            .I(N__41900));
    Span4Mux_v I__8634 (
            .O(N__41904),
            .I(N__41897));
    SRMux I__8633 (
            .O(N__41903),
            .I(N__41894));
    Span4Mux_h I__8632 (
            .O(N__41900),
            .I(N__41891));
    Span4Mux_h I__8631 (
            .O(N__41897),
            .I(N__41886));
    LocalMux I__8630 (
            .O(N__41894),
            .I(N__41886));
    Span4Mux_h I__8629 (
            .O(N__41891),
            .I(N__41883));
    Span4Mux_v I__8628 (
            .O(N__41886),
            .I(N__41880));
    Span4Mux_v I__8627 (
            .O(N__41883),
            .I(N__41877));
    Odrv4 I__8626 (
            .O(N__41880),
            .I(\comm_spi.data_tx_7__N_854 ));
    Odrv4 I__8625 (
            .O(N__41877),
            .I(\comm_spi.data_tx_7__N_854 ));
    InMux I__8624 (
            .O(N__41872),
            .I(N__41868));
    InMux I__8623 (
            .O(N__41871),
            .I(N__41864));
    LocalMux I__8622 (
            .O(N__41868),
            .I(N__41861));
    InMux I__8621 (
            .O(N__41867),
            .I(N__41858));
    LocalMux I__8620 (
            .O(N__41864),
            .I(N__41855));
    Span4Mux_h I__8619 (
            .O(N__41861),
            .I(N__41852));
    LocalMux I__8618 (
            .O(N__41858),
            .I(N__41849));
    Span4Mux_v I__8617 (
            .O(N__41855),
            .I(N__41846));
    Span4Mux_v I__8616 (
            .O(N__41852),
            .I(N__41843));
    Odrv4 I__8615 (
            .O(N__41849),
            .I(comm_test_buf_24_1));
    Odrv4 I__8614 (
            .O(N__41846),
            .I(comm_test_buf_24_1));
    Odrv4 I__8613 (
            .O(N__41843),
            .I(comm_test_buf_24_1));
    InMux I__8612 (
            .O(N__41836),
            .I(N__41833));
    LocalMux I__8611 (
            .O(N__41833),
            .I(N__41830));
    Span4Mux_v I__8610 (
            .O(N__41830),
            .I(N__41827));
    Odrv4 I__8609 (
            .O(N__41827),
            .I(n111_adj_1798));
    InMux I__8608 (
            .O(N__41824),
            .I(N__41821));
    LocalMux I__8607 (
            .O(N__41821),
            .I(N__41818));
    Span4Mux_v I__8606 (
            .O(N__41818),
            .I(N__41815));
    Span4Mux_v I__8605 (
            .O(N__41815),
            .I(N__41812));
    Odrv4 I__8604 (
            .O(N__41812),
            .I(n21965));
    CascadeMux I__8603 (
            .O(N__41809),
            .I(n12056_cascade_));
    InMux I__8602 (
            .O(N__41806),
            .I(N__41803));
    LocalMux I__8601 (
            .O(N__41803),
            .I(N__41800));
    Span4Mux_h I__8600 (
            .O(N__41800),
            .I(N__41797));
    Span4Mux_h I__8599 (
            .O(N__41797),
            .I(N__41794));
    Odrv4 I__8598 (
            .O(N__41794),
            .I(buf_data_iac_12));
    InMux I__8597 (
            .O(N__41791),
            .I(N__41786));
    InMux I__8596 (
            .O(N__41790),
            .I(N__41783));
    InMux I__8595 (
            .O(N__41789),
            .I(N__41780));
    LocalMux I__8594 (
            .O(N__41786),
            .I(data_index_2));
    LocalMux I__8593 (
            .O(N__41783),
            .I(data_index_2));
    LocalMux I__8592 (
            .O(N__41780),
            .I(data_index_2));
    InMux I__8591 (
            .O(N__41773),
            .I(N__41770));
    LocalMux I__8590 (
            .O(N__41770),
            .I(n8_adj_1628));
    CascadeMux I__8589 (
            .O(N__41767),
            .I(n8_adj_1628_cascade_));
    InMux I__8588 (
            .O(N__41764),
            .I(N__41758));
    InMux I__8587 (
            .O(N__41763),
            .I(N__41758));
    LocalMux I__8586 (
            .O(N__41758),
            .I(n7_adj_1627));
    CascadeMux I__8585 (
            .O(N__41755),
            .I(N__41752));
    CascadeBuf I__8584 (
            .O(N__41752),
            .I(N__41749));
    CascadeMux I__8583 (
            .O(N__41749),
            .I(N__41746));
    CascadeBuf I__8582 (
            .O(N__41746),
            .I(N__41743));
    CascadeMux I__8581 (
            .O(N__41743),
            .I(N__41740));
    CascadeBuf I__8580 (
            .O(N__41740),
            .I(N__41737));
    CascadeMux I__8579 (
            .O(N__41737),
            .I(N__41734));
    CascadeBuf I__8578 (
            .O(N__41734),
            .I(N__41731));
    CascadeMux I__8577 (
            .O(N__41731),
            .I(N__41728));
    CascadeBuf I__8576 (
            .O(N__41728),
            .I(N__41725));
    CascadeMux I__8575 (
            .O(N__41725),
            .I(N__41722));
    CascadeBuf I__8574 (
            .O(N__41722),
            .I(N__41719));
    CascadeMux I__8573 (
            .O(N__41719),
            .I(N__41715));
    CascadeMux I__8572 (
            .O(N__41718),
            .I(N__41712));
    CascadeBuf I__8571 (
            .O(N__41715),
            .I(N__41709));
    CascadeBuf I__8570 (
            .O(N__41712),
            .I(N__41706));
    CascadeMux I__8569 (
            .O(N__41709),
            .I(N__41703));
    CascadeMux I__8568 (
            .O(N__41706),
            .I(N__41700));
    CascadeBuf I__8567 (
            .O(N__41703),
            .I(N__41697));
    InMux I__8566 (
            .O(N__41700),
            .I(N__41694));
    CascadeMux I__8565 (
            .O(N__41697),
            .I(N__41691));
    LocalMux I__8564 (
            .O(N__41694),
            .I(N__41688));
    CascadeBuf I__8563 (
            .O(N__41691),
            .I(N__41685));
    Span4Mux_h I__8562 (
            .O(N__41688),
            .I(N__41682));
    CascadeMux I__8561 (
            .O(N__41685),
            .I(N__41679));
    Span4Mux_v I__8560 (
            .O(N__41682),
            .I(N__41676));
    InMux I__8559 (
            .O(N__41679),
            .I(N__41673));
    Span4Mux_v I__8558 (
            .O(N__41676),
            .I(N__41670));
    LocalMux I__8557 (
            .O(N__41673),
            .I(N__41667));
    Span4Mux_h I__8556 (
            .O(N__41670),
            .I(N__41664));
    Span4Mux_h I__8555 (
            .O(N__41667),
            .I(N__41661));
    Span4Mux_h I__8554 (
            .O(N__41664),
            .I(N__41656));
    Span4Mux_h I__8553 (
            .O(N__41661),
            .I(N__41656));
    Odrv4 I__8552 (
            .O(N__41656),
            .I(data_index_9_N_236_2));
    InMux I__8551 (
            .O(N__41653),
            .I(N__41649));
    InMux I__8550 (
            .O(N__41652),
            .I(N__41646));
    LocalMux I__8549 (
            .O(N__41649),
            .I(n18865));
    LocalMux I__8548 (
            .O(N__41646),
            .I(n18865));
    InMux I__8547 (
            .O(N__41641),
            .I(N__41637));
    InMux I__8546 (
            .O(N__41640),
            .I(N__41634));
    LocalMux I__8545 (
            .O(N__41637),
            .I(N__41631));
    LocalMux I__8544 (
            .O(N__41634),
            .I(n7_adj_1626));
    Odrv4 I__8543 (
            .O(N__41631),
            .I(n7_adj_1626));
    InMux I__8542 (
            .O(N__41626),
            .I(N__41621));
    InMux I__8541 (
            .O(N__41625),
            .I(N__41618));
    InMux I__8540 (
            .O(N__41624),
            .I(N__41615));
    LocalMux I__8539 (
            .O(N__41621),
            .I(data_index_3));
    LocalMux I__8538 (
            .O(N__41618),
            .I(data_index_3));
    LocalMux I__8537 (
            .O(N__41615),
            .I(data_index_3));
    InMux I__8536 (
            .O(N__41608),
            .I(N__41605));
    LocalMux I__8535 (
            .O(N__41605),
            .I(N__41602));
    Span4Mux_h I__8534 (
            .O(N__41602),
            .I(N__41598));
    InMux I__8533 (
            .O(N__41601),
            .I(N__41595));
    Span4Mux_h I__8532 (
            .O(N__41598),
            .I(N__41592));
    LocalMux I__8531 (
            .O(N__41595),
            .I(acadc_skipcnt_8));
    Odrv4 I__8530 (
            .O(N__41592),
            .I(acadc_skipcnt_8));
    CascadeMux I__8529 (
            .O(N__41587),
            .I(N__41584));
    InMux I__8528 (
            .O(N__41584),
            .I(N__41581));
    LocalMux I__8527 (
            .O(N__41581),
            .I(N__41578));
    Odrv4 I__8526 (
            .O(N__41578),
            .I(n20));
    InMux I__8525 (
            .O(N__41575),
            .I(N__41572));
    LocalMux I__8524 (
            .O(N__41572),
            .I(n14_adj_1599));
    InMux I__8523 (
            .O(N__41569),
            .I(N__41566));
    LocalMux I__8522 (
            .O(N__41566),
            .I(N__41563));
    Odrv4 I__8521 (
            .O(N__41563),
            .I(n17));
    CascadeMux I__8520 (
            .O(N__41560),
            .I(n26_cascade_));
    InMux I__8519 (
            .O(N__41557),
            .I(N__41554));
    LocalMux I__8518 (
            .O(N__41554),
            .I(n30_adj_1743));
    InMux I__8517 (
            .O(N__41551),
            .I(N__41548));
    LocalMux I__8516 (
            .O(N__41548),
            .I(N__41545));
    Span4Mux_h I__8515 (
            .O(N__41545),
            .I(N__41541));
    InMux I__8514 (
            .O(N__41544),
            .I(N__41538));
    Odrv4 I__8513 (
            .O(N__41541),
            .I(n31));
    LocalMux I__8512 (
            .O(N__41538),
            .I(n31));
    InMux I__8511 (
            .O(N__41533),
            .I(N__41530));
    LocalMux I__8510 (
            .O(N__41530),
            .I(N__41527));
    Span4Mux_h I__8509 (
            .O(N__41527),
            .I(N__41523));
    InMux I__8508 (
            .O(N__41526),
            .I(N__41520));
    Span4Mux_v I__8507 (
            .O(N__41523),
            .I(N__41517));
    LocalMux I__8506 (
            .O(N__41520),
            .I(acadc_skipcnt_3));
    Odrv4 I__8505 (
            .O(N__41517),
            .I(acadc_skipcnt_3));
    InMux I__8504 (
            .O(N__41512),
            .I(N__41507));
    CascadeMux I__8503 (
            .O(N__41511),
            .I(N__41504));
    CascadeMux I__8502 (
            .O(N__41510),
            .I(N__41501));
    LocalMux I__8501 (
            .O(N__41507),
            .I(N__41498));
    InMux I__8500 (
            .O(N__41504),
            .I(N__41495));
    InMux I__8499 (
            .O(N__41501),
            .I(N__41492));
    Span4Mux_h I__8498 (
            .O(N__41498),
            .I(N__41487));
    LocalMux I__8497 (
            .O(N__41495),
            .I(N__41487));
    LocalMux I__8496 (
            .O(N__41492),
            .I(acadc_skipCount_15));
    Odrv4 I__8495 (
            .O(N__41487),
            .I(acadc_skipCount_15));
    InMux I__8494 (
            .O(N__41482),
            .I(N__41479));
    LocalMux I__8493 (
            .O(N__41479),
            .I(N__41476));
    Span4Mux_h I__8492 (
            .O(N__41476),
            .I(N__41473));
    Odrv4 I__8491 (
            .O(N__41473),
            .I(n23_adj_1756));
    InMux I__8490 (
            .O(N__41470),
            .I(N__41467));
    LocalMux I__8489 (
            .O(N__41467),
            .I(n21_adj_1803));
    InMux I__8488 (
            .O(N__41464),
            .I(N__41461));
    LocalMux I__8487 (
            .O(N__41461),
            .I(N__41458));
    Odrv4 I__8486 (
            .O(N__41458),
            .I(n30_adj_1769));
    InMux I__8485 (
            .O(N__41455),
            .I(N__41452));
    LocalMux I__8484 (
            .O(N__41452),
            .I(N__41449));
    Odrv4 I__8483 (
            .O(N__41449),
            .I(n22167));
    CascadeMux I__8482 (
            .O(N__41446),
            .I(N__41443));
    InMux I__8481 (
            .O(N__41443),
            .I(N__41440));
    LocalMux I__8480 (
            .O(N__41440),
            .I(N__41437));
    Span4Mux_h I__8479 (
            .O(N__41437),
            .I(N__41434));
    Odrv4 I__8478 (
            .O(N__41434),
            .I(n22166));
    InMux I__8477 (
            .O(N__41431),
            .I(N__41428));
    LocalMux I__8476 (
            .O(N__41428),
            .I(N__41425));
    Span4Mux_h I__8475 (
            .O(N__41425),
            .I(N__41422));
    Span4Mux_h I__8474 (
            .O(N__41422),
            .I(N__41419));
    Odrv4 I__8473 (
            .O(N__41419),
            .I(n23471));
    CascadeMux I__8472 (
            .O(N__41416),
            .I(n23549_cascade_));
    InMux I__8471 (
            .O(N__41413),
            .I(N__41410));
    LocalMux I__8470 (
            .O(N__41410),
            .I(n22174));
    InMux I__8469 (
            .O(N__41407),
            .I(N__41404));
    LocalMux I__8468 (
            .O(N__41404),
            .I(N__41401));
    Span4Mux_v I__8467 (
            .O(N__41401),
            .I(N__41397));
    InMux I__8466 (
            .O(N__41400),
            .I(N__41394));
    Odrv4 I__8465 (
            .O(N__41397),
            .I(n112));
    LocalMux I__8464 (
            .O(N__41394),
            .I(n112));
    InMux I__8463 (
            .O(N__41389),
            .I(N__41386));
    LocalMux I__8462 (
            .O(N__41386),
            .I(N__41383));
    Span4Mux_v I__8461 (
            .O(N__41383),
            .I(N__41380));
    Span4Mux_h I__8460 (
            .O(N__41380),
            .I(N__41377));
    Span4Mux_h I__8459 (
            .O(N__41377),
            .I(N__41374));
    Odrv4 I__8458 (
            .O(N__41374),
            .I(n30_adj_1805));
    InMux I__8457 (
            .O(N__41371),
            .I(N__41367));
    InMux I__8456 (
            .O(N__41370),
            .I(N__41364));
    LocalMux I__8455 (
            .O(N__41367),
            .I(N__41361));
    LocalMux I__8454 (
            .O(N__41364),
            .I(N__41358));
    Odrv4 I__8453 (
            .O(N__41361),
            .I(n17650));
    Odrv12 I__8452 (
            .O(N__41358),
            .I(n17650));
    InMux I__8451 (
            .O(N__41353),
            .I(N__41350));
    LocalMux I__8450 (
            .O(N__41350),
            .I(N__41346));
    InMux I__8449 (
            .O(N__41349),
            .I(N__41343));
    Odrv4 I__8448 (
            .O(N__41346),
            .I(n12));
    LocalMux I__8447 (
            .O(N__41343),
            .I(n12));
    SRMux I__8446 (
            .O(N__41338),
            .I(N__41335));
    LocalMux I__8445 (
            .O(N__41335),
            .I(N__41332));
    Span4Mux_h I__8444 (
            .O(N__41332),
            .I(N__41329));
    Odrv4 I__8443 (
            .O(N__41329),
            .I(n15553));
    InMux I__8442 (
            .O(N__41326),
            .I(N__41323));
    LocalMux I__8441 (
            .O(N__41323),
            .I(N__41320));
    Span4Mux_v I__8440 (
            .O(N__41320),
            .I(N__41317));
    Span4Mux_h I__8439 (
            .O(N__41317),
            .I(N__41314));
    Odrv4 I__8438 (
            .O(N__41314),
            .I(n16_adj_1721));
    CascadeMux I__8437 (
            .O(N__41311),
            .I(N__41307));
    InMux I__8436 (
            .O(N__41310),
            .I(N__41304));
    InMux I__8435 (
            .O(N__41307),
            .I(N__41301));
    LocalMux I__8434 (
            .O(N__41304),
            .I(N__41298));
    LocalMux I__8433 (
            .O(N__41301),
            .I(N__41294));
    Span4Mux_v I__8432 (
            .O(N__41298),
            .I(N__41291));
    CascadeMux I__8431 (
            .O(N__41297),
            .I(N__41288));
    Span4Mux_h I__8430 (
            .O(N__41294),
            .I(N__41285));
    Sp12to4 I__8429 (
            .O(N__41291),
            .I(N__41282));
    InMux I__8428 (
            .O(N__41288),
            .I(N__41279));
    Span4Mux_h I__8427 (
            .O(N__41285),
            .I(N__41276));
    Span12Mux_h I__8426 (
            .O(N__41282),
            .I(N__41273));
    LocalMux I__8425 (
            .O(N__41279),
            .I(buf_adcdata_iac_14));
    Odrv4 I__8424 (
            .O(N__41276),
            .I(buf_adcdata_iac_14));
    Odrv12 I__8423 (
            .O(N__41273),
            .I(buf_adcdata_iac_14));
    CascadeMux I__8422 (
            .O(N__41266),
            .I(N__41262));
    InMux I__8421 (
            .O(N__41265),
            .I(N__41257));
    InMux I__8420 (
            .O(N__41262),
            .I(N__41257));
    LocalMux I__8419 (
            .O(N__41257),
            .I(n12015));
    CascadeMux I__8418 (
            .O(N__41254),
            .I(n8_cascade_));
    InMux I__8417 (
            .O(N__41251),
            .I(N__41248));
    LocalMux I__8416 (
            .O(N__41248),
            .I(N__41245));
    Span4Mux_v I__8415 (
            .O(N__41245),
            .I(N__41242));
    Span4Mux_h I__8414 (
            .O(N__41242),
            .I(N__41238));
    InMux I__8413 (
            .O(N__41241),
            .I(N__41235));
    Odrv4 I__8412 (
            .O(N__41238),
            .I(buf_adcdata_vdc_11));
    LocalMux I__8411 (
            .O(N__41235),
            .I(buf_adcdata_vdc_11));
    InMux I__8410 (
            .O(N__41230),
            .I(N__41227));
    LocalMux I__8409 (
            .O(N__41227),
            .I(N__41224));
    Span4Mux_v I__8408 (
            .O(N__41224),
            .I(N__41221));
    Span4Mux_h I__8407 (
            .O(N__41221),
            .I(N__41217));
    InMux I__8406 (
            .O(N__41220),
            .I(N__41214));
    Span4Mux_h I__8405 (
            .O(N__41217),
            .I(N__41209));
    LocalMux I__8404 (
            .O(N__41214),
            .I(N__41209));
    Span4Mux_v I__8403 (
            .O(N__41209),
            .I(N__41205));
    InMux I__8402 (
            .O(N__41208),
            .I(N__41202));
    Span4Mux_h I__8401 (
            .O(N__41205),
            .I(N__41199));
    LocalMux I__8400 (
            .O(N__41202),
            .I(buf_adcdata_vac_11));
    Odrv4 I__8399 (
            .O(N__41199),
            .I(buf_adcdata_vac_11));
    InMux I__8398 (
            .O(N__41194),
            .I(N__41191));
    LocalMux I__8397 (
            .O(N__41191),
            .I(n22092));
    CEMux I__8396 (
            .O(N__41188),
            .I(N__41184));
    InMux I__8395 (
            .O(N__41187),
            .I(N__41181));
    LocalMux I__8394 (
            .O(N__41184),
            .I(N__41178));
    LocalMux I__8393 (
            .O(N__41181),
            .I(N__41175));
    Span12Mux_h I__8392 (
            .O(N__41178),
            .I(N__41172));
    Span4Mux_h I__8391 (
            .O(N__41175),
            .I(N__41169));
    Odrv12 I__8390 (
            .O(N__41172),
            .I(n13211));
    Odrv4 I__8389 (
            .O(N__41169),
            .I(n13211));
    InMux I__8388 (
            .O(N__41164),
            .I(N__41161));
    LocalMux I__8387 (
            .O(N__41161),
            .I(N__41158));
    Span4Mux_h I__8386 (
            .O(N__41158),
            .I(N__41154));
    InMux I__8385 (
            .O(N__41157),
            .I(N__41151));
    Span4Mux_v I__8384 (
            .O(N__41154),
            .I(N__41148));
    LocalMux I__8383 (
            .O(N__41151),
            .I(acadc_skipcnt_5));
    Odrv4 I__8382 (
            .O(N__41148),
            .I(acadc_skipcnt_5));
    InMux I__8381 (
            .O(N__41143),
            .I(N__41140));
    LocalMux I__8380 (
            .O(N__41140),
            .I(N__41137));
    Span4Mux_v I__8379 (
            .O(N__41137),
            .I(N__41134));
    Span4Mux_h I__8378 (
            .O(N__41134),
            .I(N__41131));
    Odrv4 I__8377 (
            .O(N__41131),
            .I(buf_data_vac_18));
    InMux I__8376 (
            .O(N__41128),
            .I(N__41125));
    LocalMux I__8375 (
            .O(N__41125),
            .I(comm_buf_3_2));
    InMux I__8374 (
            .O(N__41122),
            .I(N__41119));
    LocalMux I__8373 (
            .O(N__41119),
            .I(N__41116));
    Span4Mux_h I__8372 (
            .O(N__41116),
            .I(N__41113));
    Span4Mux_h I__8371 (
            .O(N__41113),
            .I(N__41110));
    Odrv4 I__8370 (
            .O(N__41110),
            .I(buf_data_vac_17));
    InMux I__8369 (
            .O(N__41107),
            .I(N__41104));
    LocalMux I__8368 (
            .O(N__41104),
            .I(N__41101));
    Span4Mux_v I__8367 (
            .O(N__41101),
            .I(N__41098));
    Odrv4 I__8366 (
            .O(N__41098),
            .I(comm_buf_3_1));
    SRMux I__8365 (
            .O(N__41095),
            .I(N__41092));
    LocalMux I__8364 (
            .O(N__41092),
            .I(N__41089));
    Span4Mux_h I__8363 (
            .O(N__41089),
            .I(N__41086));
    Span4Mux_h I__8362 (
            .O(N__41086),
            .I(N__41083));
    Odrv4 I__8361 (
            .O(N__41083),
            .I(n15503));
    InMux I__8360 (
            .O(N__41080),
            .I(N__41077));
    LocalMux I__8359 (
            .O(N__41077),
            .I(N__41074));
    Odrv12 I__8358 (
            .O(N__41074),
            .I(n30_adj_1708));
    InMux I__8357 (
            .O(N__41071),
            .I(N__41068));
    LocalMux I__8356 (
            .O(N__41068),
            .I(N__41063));
    InMux I__8355 (
            .O(N__41067),
            .I(N__41058));
    InMux I__8354 (
            .O(N__41066),
            .I(N__41058));
    Span12Mux_h I__8353 (
            .O(N__41063),
            .I(N__41055));
    LocalMux I__8352 (
            .O(N__41058),
            .I(N__41052));
    Odrv12 I__8351 (
            .O(N__41055),
            .I(comm_test_buf_24_2));
    Odrv4 I__8350 (
            .O(N__41052),
            .I(comm_test_buf_24_2));
    InMux I__8349 (
            .O(N__41047),
            .I(N__41044));
    LocalMux I__8348 (
            .O(N__41044),
            .I(N__41041));
    Odrv4 I__8347 (
            .O(N__41041),
            .I(comm_buf_2_7_N_575_2));
    CEMux I__8346 (
            .O(N__41038),
            .I(N__41035));
    LocalMux I__8345 (
            .O(N__41035),
            .I(N__41032));
    Span4Mux_v I__8344 (
            .O(N__41032),
            .I(N__41028));
    InMux I__8343 (
            .O(N__41031),
            .I(N__41025));
    Odrv4 I__8342 (
            .O(N__41028),
            .I(n12880));
    LocalMux I__8341 (
            .O(N__41025),
            .I(n12880));
    InMux I__8340 (
            .O(N__41020),
            .I(N__41016));
    InMux I__8339 (
            .O(N__41019),
            .I(N__41012));
    LocalMux I__8338 (
            .O(N__41016),
            .I(N__41009));
    InMux I__8337 (
            .O(N__41015),
            .I(N__41006));
    LocalMux I__8336 (
            .O(N__41012),
            .I(N__41002));
    Span4Mux_h I__8335 (
            .O(N__41009),
            .I(N__40997));
    LocalMux I__8334 (
            .O(N__41006),
            .I(N__40997));
    InMux I__8333 (
            .O(N__41005),
            .I(N__40994));
    Span4Mux_h I__8332 (
            .O(N__41002),
            .I(N__40991));
    Span4Mux_v I__8331 (
            .O(N__40997),
            .I(N__40986));
    LocalMux I__8330 (
            .O(N__40994),
            .I(N__40986));
    Odrv4 I__8329 (
            .O(N__40991),
            .I(n21886));
    Odrv4 I__8328 (
            .O(N__40986),
            .I(n21886));
    CascadeMux I__8327 (
            .O(N__40981),
            .I(n12_cascade_));
    CascadeMux I__8326 (
            .O(N__40978),
            .I(N__40975));
    InMux I__8325 (
            .O(N__40975),
            .I(N__40970));
    InMux I__8324 (
            .O(N__40974),
            .I(N__40965));
    InMux I__8323 (
            .O(N__40973),
            .I(N__40965));
    LocalMux I__8322 (
            .O(N__40970),
            .I(N__40962));
    LocalMux I__8321 (
            .O(N__40965),
            .I(N__40959));
    Span4Mux_v I__8320 (
            .O(N__40962),
            .I(N__40956));
    Span4Mux_v I__8319 (
            .O(N__40959),
            .I(N__40953));
    Odrv4 I__8318 (
            .O(N__40956),
            .I(comm_buf_2_2));
    Odrv4 I__8317 (
            .O(N__40953),
            .I(comm_buf_2_2));
    InMux I__8316 (
            .O(N__40948),
            .I(N__40944));
    CascadeMux I__8315 (
            .O(N__40947),
            .I(N__40941));
    LocalMux I__8314 (
            .O(N__40944),
            .I(N__40936));
    InMux I__8313 (
            .O(N__40941),
            .I(N__40932));
    InMux I__8312 (
            .O(N__40940),
            .I(N__40929));
    CascadeMux I__8311 (
            .O(N__40939),
            .I(N__40926));
    Span4Mux_v I__8310 (
            .O(N__40936),
            .I(N__40921));
    InMux I__8309 (
            .O(N__40935),
            .I(N__40918));
    LocalMux I__8308 (
            .O(N__40932),
            .I(N__40915));
    LocalMux I__8307 (
            .O(N__40929),
            .I(N__40912));
    InMux I__8306 (
            .O(N__40926),
            .I(N__40907));
    InMux I__8305 (
            .O(N__40925),
            .I(N__40907));
    CascadeMux I__8304 (
            .O(N__40924),
            .I(N__40904));
    Span4Mux_h I__8303 (
            .O(N__40921),
            .I(N__40899));
    LocalMux I__8302 (
            .O(N__40918),
            .I(N__40899));
    Span4Mux_h I__8301 (
            .O(N__40915),
            .I(N__40894));
    Span4Mux_v I__8300 (
            .O(N__40912),
            .I(N__40894));
    LocalMux I__8299 (
            .O(N__40907),
            .I(N__40891));
    InMux I__8298 (
            .O(N__40904),
            .I(N__40887));
    Span4Mux_v I__8297 (
            .O(N__40899),
            .I(N__40884));
    Span4Mux_h I__8296 (
            .O(N__40894),
            .I(N__40879));
    Span4Mux_h I__8295 (
            .O(N__40891),
            .I(N__40879));
    InMux I__8294 (
            .O(N__40890),
            .I(N__40876));
    LocalMux I__8293 (
            .O(N__40887),
            .I(comm_buf_0_2));
    Odrv4 I__8292 (
            .O(N__40884),
            .I(comm_buf_0_2));
    Odrv4 I__8291 (
            .O(N__40879),
            .I(comm_buf_0_2));
    LocalMux I__8290 (
            .O(N__40876),
            .I(comm_buf_0_2));
    InMux I__8289 (
            .O(N__40867),
            .I(N__40864));
    LocalMux I__8288 (
            .O(N__40864),
            .I(N__40861));
    Span4Mux_h I__8287 (
            .O(N__40861),
            .I(N__40858));
    Odrv4 I__8286 (
            .O(N__40858),
            .I(n13207));
    InMux I__8285 (
            .O(N__40855),
            .I(N__40849));
    InMux I__8284 (
            .O(N__40854),
            .I(N__40849));
    LocalMux I__8283 (
            .O(N__40849),
            .I(N__40846));
    Span4Mux_v I__8282 (
            .O(N__40846),
            .I(N__40842));
    InMux I__8281 (
            .O(N__40845),
            .I(N__40839));
    Odrv4 I__8280 (
            .O(N__40842),
            .I(comm_tx_buf_2));
    LocalMux I__8279 (
            .O(N__40839),
            .I(comm_tx_buf_2));
    SRMux I__8278 (
            .O(N__40834),
            .I(N__40831));
    LocalMux I__8277 (
            .O(N__40831),
            .I(N__40828));
    Span4Mux_v I__8276 (
            .O(N__40828),
            .I(N__40825));
    Span4Mux_v I__8275 (
            .O(N__40825),
            .I(N__40822));
    Sp12to4 I__8274 (
            .O(N__40822),
            .I(N__40819));
    Odrv12 I__8273 (
            .O(N__40819),
            .I(\comm_spi.data_tx_7__N_877 ));
    InMux I__8272 (
            .O(N__40816),
            .I(N__40813));
    LocalMux I__8271 (
            .O(N__40813),
            .I(N__40810));
    Span4Mux_h I__8270 (
            .O(N__40810),
            .I(N__40807));
    Span4Mux_h I__8269 (
            .O(N__40807),
            .I(N__40804));
    Odrv4 I__8268 (
            .O(N__40804),
            .I(buf_data_vac_16));
    InMux I__8267 (
            .O(N__40801),
            .I(N__40798));
    LocalMux I__8266 (
            .O(N__40798),
            .I(N__40795));
    Span4Mux_v I__8265 (
            .O(N__40795),
            .I(N__40792));
    Sp12to4 I__8264 (
            .O(N__40792),
            .I(N__40789));
    Span12Mux_h I__8263 (
            .O(N__40789),
            .I(N__40786));
    Odrv12 I__8262 (
            .O(N__40786),
            .I(buf_data_vac_23));
    InMux I__8261 (
            .O(N__40783),
            .I(N__40780));
    LocalMux I__8260 (
            .O(N__40780),
            .I(N__40777));
    Odrv4 I__8259 (
            .O(N__40777),
            .I(comm_buf_3_7));
    InMux I__8258 (
            .O(N__40774),
            .I(N__40771));
    LocalMux I__8257 (
            .O(N__40771),
            .I(N__40768));
    Span4Mux_v I__8256 (
            .O(N__40768),
            .I(N__40765));
    Span4Mux_h I__8255 (
            .O(N__40765),
            .I(N__40762));
    Span4Mux_h I__8254 (
            .O(N__40762),
            .I(N__40759));
    Span4Mux_v I__8253 (
            .O(N__40759),
            .I(N__40756));
    Odrv4 I__8252 (
            .O(N__40756),
            .I(buf_data_vac_22));
    InMux I__8251 (
            .O(N__40753),
            .I(N__40750));
    LocalMux I__8250 (
            .O(N__40750),
            .I(N__40747));
    Span4Mux_v I__8249 (
            .O(N__40747),
            .I(N__40744));
    Span4Mux_h I__8248 (
            .O(N__40744),
            .I(N__40741));
    Odrv4 I__8247 (
            .O(N__40741),
            .I(comm_buf_3_6));
    InMux I__8246 (
            .O(N__40738),
            .I(N__40735));
    LocalMux I__8245 (
            .O(N__40735),
            .I(N__40732));
    Span4Mux_h I__8244 (
            .O(N__40732),
            .I(N__40729));
    Span4Mux_h I__8243 (
            .O(N__40729),
            .I(N__40726));
    Span4Mux_v I__8242 (
            .O(N__40726),
            .I(N__40723));
    Span4Mux_v I__8241 (
            .O(N__40723),
            .I(N__40720));
    Odrv4 I__8240 (
            .O(N__40720),
            .I(buf_data_vac_21));
    InMux I__8239 (
            .O(N__40717),
            .I(N__40714));
    LocalMux I__8238 (
            .O(N__40714),
            .I(N__40711));
    Span4Mux_h I__8237 (
            .O(N__40711),
            .I(N__40708));
    Span4Mux_v I__8236 (
            .O(N__40708),
            .I(N__40705));
    Span4Mux_h I__8235 (
            .O(N__40705),
            .I(N__40702));
    Odrv4 I__8234 (
            .O(N__40702),
            .I(buf_data_vac_20));
    InMux I__8233 (
            .O(N__40699),
            .I(N__40696));
    LocalMux I__8232 (
            .O(N__40696),
            .I(N__40693));
    Span4Mux_v I__8231 (
            .O(N__40693),
            .I(N__40690));
    Odrv4 I__8230 (
            .O(N__40690),
            .I(comm_buf_3_4));
    InMux I__8229 (
            .O(N__40687),
            .I(N__40684));
    LocalMux I__8228 (
            .O(N__40684),
            .I(N__40681));
    Span4Mux_h I__8227 (
            .O(N__40681),
            .I(N__40678));
    Span4Mux_h I__8226 (
            .O(N__40678),
            .I(N__40675));
    Span4Mux_h I__8225 (
            .O(N__40675),
            .I(N__40672));
    Odrv4 I__8224 (
            .O(N__40672),
            .I(buf_data_vac_19));
    InMux I__8223 (
            .O(N__40669),
            .I(N__40666));
    LocalMux I__8222 (
            .O(N__40666),
            .I(n4_adj_1664));
    InMux I__8221 (
            .O(N__40663),
            .I(N__40660));
    LocalMux I__8220 (
            .O(N__40660),
            .I(n1));
    InMux I__8219 (
            .O(N__40657),
            .I(N__40654));
    LocalMux I__8218 (
            .O(N__40654),
            .I(N__40651));
    Span4Mux_v I__8217 (
            .O(N__40651),
            .I(N__40647));
    CascadeMux I__8216 (
            .O(N__40650),
            .I(N__40644));
    Span4Mux_h I__8215 (
            .O(N__40647),
            .I(N__40640));
    InMux I__8214 (
            .O(N__40644),
            .I(N__40635));
    InMux I__8213 (
            .O(N__40643),
            .I(N__40635));
    Odrv4 I__8212 (
            .O(N__40640),
            .I(comm_tx_buf_7));
    LocalMux I__8211 (
            .O(N__40635),
            .I(comm_tx_buf_7));
    SRMux I__8210 (
            .O(N__40630),
            .I(N__40626));
    SRMux I__8209 (
            .O(N__40629),
            .I(N__40623));
    LocalMux I__8208 (
            .O(N__40626),
            .I(N__40620));
    LocalMux I__8207 (
            .O(N__40623),
            .I(N__40616));
    Span4Mux_v I__8206 (
            .O(N__40620),
            .I(N__40613));
    SRMux I__8205 (
            .O(N__40619),
            .I(N__40610));
    Span4Mux_v I__8204 (
            .O(N__40616),
            .I(N__40603));
    Span4Mux_h I__8203 (
            .O(N__40613),
            .I(N__40603));
    LocalMux I__8202 (
            .O(N__40610),
            .I(N__40603));
    Span4Mux_h I__8201 (
            .O(N__40603),
            .I(N__40600));
    Odrv4 I__8200 (
            .O(N__40600),
            .I(\comm_spi.data_tx_7__N_862 ));
    InMux I__8199 (
            .O(N__40597),
            .I(N__40594));
    LocalMux I__8198 (
            .O(N__40594),
            .I(n4_adj_1673));
    CascadeMux I__8197 (
            .O(N__40591),
            .I(n22342_cascade_));
    InMux I__8196 (
            .O(N__40588),
            .I(N__40585));
    LocalMux I__8195 (
            .O(N__40585),
            .I(n23396));
    CascadeMux I__8194 (
            .O(N__40582),
            .I(n1_adj_1671_cascade_));
    InMux I__8193 (
            .O(N__40579),
            .I(N__40576));
    LocalMux I__8192 (
            .O(N__40576),
            .I(N__40573));
    Odrv12 I__8191 (
            .O(N__40573),
            .I(n2_adj_1672));
    CascadeMux I__8190 (
            .O(N__40570),
            .I(N__40565));
    CascadeMux I__8189 (
            .O(N__40569),
            .I(N__40558));
    CascadeMux I__8188 (
            .O(N__40568),
            .I(N__40555));
    InMux I__8187 (
            .O(N__40565),
            .I(N__40552));
    CascadeMux I__8186 (
            .O(N__40564),
            .I(N__40549));
    InMux I__8185 (
            .O(N__40563),
            .I(N__40546));
    InMux I__8184 (
            .O(N__40562),
            .I(N__40543));
    InMux I__8183 (
            .O(N__40561),
            .I(N__40540));
    InMux I__8182 (
            .O(N__40558),
            .I(N__40536));
    InMux I__8181 (
            .O(N__40555),
            .I(N__40533));
    LocalMux I__8180 (
            .O(N__40552),
            .I(N__40530));
    InMux I__8179 (
            .O(N__40549),
            .I(N__40527));
    LocalMux I__8178 (
            .O(N__40546),
            .I(N__40523));
    LocalMux I__8177 (
            .O(N__40543),
            .I(N__40518));
    LocalMux I__8176 (
            .O(N__40540),
            .I(N__40518));
    InMux I__8175 (
            .O(N__40539),
            .I(N__40514));
    LocalMux I__8174 (
            .O(N__40536),
            .I(N__40509));
    LocalMux I__8173 (
            .O(N__40533),
            .I(N__40509));
    Span4Mux_v I__8172 (
            .O(N__40530),
            .I(N__40504));
    LocalMux I__8171 (
            .O(N__40527),
            .I(N__40504));
    InMux I__8170 (
            .O(N__40526),
            .I(N__40500));
    Sp12to4 I__8169 (
            .O(N__40523),
            .I(N__40497));
    Span4Mux_h I__8168 (
            .O(N__40518),
            .I(N__40494));
    InMux I__8167 (
            .O(N__40517),
            .I(N__40491));
    LocalMux I__8166 (
            .O(N__40514),
            .I(N__40484));
    Span4Mux_v I__8165 (
            .O(N__40509),
            .I(N__40484));
    Span4Mux_h I__8164 (
            .O(N__40504),
            .I(N__40484));
    InMux I__8163 (
            .O(N__40503),
            .I(N__40481));
    LocalMux I__8162 (
            .O(N__40500),
            .I(N__40476));
    Span12Mux_v I__8161 (
            .O(N__40497),
            .I(N__40476));
    Odrv4 I__8160 (
            .O(N__40494),
            .I(comm_buf_0_6));
    LocalMux I__8159 (
            .O(N__40491),
            .I(comm_buf_0_6));
    Odrv4 I__8158 (
            .O(N__40484),
            .I(comm_buf_0_6));
    LocalMux I__8157 (
            .O(N__40481),
            .I(comm_buf_0_6));
    Odrv12 I__8156 (
            .O(N__40476),
            .I(comm_buf_0_6));
    InMux I__8155 (
            .O(N__40465),
            .I(N__40462));
    LocalMux I__8154 (
            .O(N__40462),
            .I(N__40458));
    InMux I__8153 (
            .O(N__40461),
            .I(N__40455));
    Odrv4 I__8152 (
            .O(N__40458),
            .I(comm_buf_6_1));
    LocalMux I__8151 (
            .O(N__40455),
            .I(comm_buf_6_1));
    InMux I__8150 (
            .O(N__40450),
            .I(N__40447));
    LocalMux I__8149 (
            .O(N__40447),
            .I(N__40444));
    Span12Mux_h I__8148 (
            .O(N__40444),
            .I(N__40441));
    Odrv12 I__8147 (
            .O(N__40441),
            .I(buf_data_iac_2));
    InMux I__8146 (
            .O(N__40438),
            .I(N__40435));
    LocalMux I__8145 (
            .O(N__40435),
            .I(N__40432));
    Odrv4 I__8144 (
            .O(N__40432),
            .I(n22_adj_1707));
    CascadeMux I__8143 (
            .O(N__40429),
            .I(N__40426));
    InMux I__8142 (
            .O(N__40426),
            .I(N__40419));
    InMux I__8141 (
            .O(N__40425),
            .I(N__40419));
    InMux I__8140 (
            .O(N__40424),
            .I(N__40416));
    LocalMux I__8139 (
            .O(N__40419),
            .I(N__40413));
    LocalMux I__8138 (
            .O(N__40416),
            .I(N__40410));
    Span4Mux_v I__8137 (
            .O(N__40413),
            .I(N__40407));
    Span4Mux_h I__8136 (
            .O(N__40410),
            .I(N__40404));
    Odrv4 I__8135 (
            .O(N__40407),
            .I(comm_buf_2_7));
    Odrv4 I__8134 (
            .O(N__40404),
            .I(comm_buf_2_7));
    CascadeMux I__8133 (
            .O(N__40399),
            .I(n22331_cascade_));
    CascadeMux I__8132 (
            .O(N__40396),
            .I(n23360_cascade_));
    InMux I__8131 (
            .O(N__40393),
            .I(N__40390));
    LocalMux I__8130 (
            .O(N__40390),
            .I(n2_adj_1663));
    InMux I__8129 (
            .O(N__40387),
            .I(n20806));
    InMux I__8128 (
            .O(N__40384),
            .I(n20807));
    InMux I__8127 (
            .O(N__40381),
            .I(n20808));
    InMux I__8126 (
            .O(N__40378),
            .I(n20809));
    InMux I__8125 (
            .O(N__40375),
            .I(n20810));
    InMux I__8124 (
            .O(N__40372),
            .I(n20811));
    InMux I__8123 (
            .O(N__40369),
            .I(N__40365));
    InMux I__8122 (
            .O(N__40368),
            .I(N__40362));
    LocalMux I__8121 (
            .O(N__40365),
            .I(secclk_cnt_19));
    LocalMux I__8120 (
            .O(N__40362),
            .I(secclk_cnt_19));
    InMux I__8119 (
            .O(N__40357),
            .I(N__40353));
    InMux I__8118 (
            .O(N__40356),
            .I(N__40350));
    LocalMux I__8117 (
            .O(N__40353),
            .I(secclk_cnt_21));
    LocalMux I__8116 (
            .O(N__40350),
            .I(secclk_cnt_21));
    CascadeMux I__8115 (
            .O(N__40345),
            .I(N__40342));
    InMux I__8114 (
            .O(N__40342),
            .I(N__40338));
    InMux I__8113 (
            .O(N__40341),
            .I(N__40335));
    LocalMux I__8112 (
            .O(N__40338),
            .I(N__40332));
    LocalMux I__8111 (
            .O(N__40335),
            .I(secclk_cnt_12));
    Odrv4 I__8110 (
            .O(N__40332),
            .I(secclk_cnt_12));
    InMux I__8109 (
            .O(N__40327),
            .I(N__40323));
    InMux I__8108 (
            .O(N__40326),
            .I(N__40320));
    LocalMux I__8107 (
            .O(N__40323),
            .I(secclk_cnt_22));
    LocalMux I__8106 (
            .O(N__40320),
            .I(secclk_cnt_22));
    InMux I__8105 (
            .O(N__40315),
            .I(bfn_14_6_0_));
    InMux I__8104 (
            .O(N__40312),
            .I(n20798));
    InMux I__8103 (
            .O(N__40309),
            .I(n20799));
    InMux I__8102 (
            .O(N__40306),
            .I(n20800));
    InMux I__8101 (
            .O(N__40303),
            .I(n20801));
    InMux I__8100 (
            .O(N__40300),
            .I(n20802));
    InMux I__8099 (
            .O(N__40297),
            .I(n20803));
    InMux I__8098 (
            .O(N__40294),
            .I(n20804));
    InMux I__8097 (
            .O(N__40291),
            .I(bfn_14_7_0_));
    InMux I__8096 (
            .O(N__40288),
            .I(N__40284));
    InMux I__8095 (
            .O(N__40287),
            .I(N__40281));
    LocalMux I__8094 (
            .O(N__40284),
            .I(\comm_spi.n15322 ));
    LocalMux I__8093 (
            .O(N__40281),
            .I(\comm_spi.n15322 ));
    SRMux I__8092 (
            .O(N__40276),
            .I(N__40273));
    LocalMux I__8091 (
            .O(N__40273),
            .I(N__40270));
    Span4Mux_h I__8090 (
            .O(N__40270),
            .I(N__40267));
    Odrv4 I__8089 (
            .O(N__40267),
            .I(\comm_spi.data_tx_7__N_861 ));
    InMux I__8088 (
            .O(N__40264),
            .I(bfn_14_5_0_));
    InMux I__8087 (
            .O(N__40261),
            .I(n20790));
    InMux I__8086 (
            .O(N__40258),
            .I(n20791));
    InMux I__8085 (
            .O(N__40255),
            .I(n20792));
    InMux I__8084 (
            .O(N__40252),
            .I(n20793));
    InMux I__8083 (
            .O(N__40249),
            .I(n20794));
    InMux I__8082 (
            .O(N__40246),
            .I(n20795));
    InMux I__8081 (
            .O(N__40243),
            .I(n20796));
    CascadeMux I__8080 (
            .O(N__40240),
            .I(N__40237));
    InMux I__8079 (
            .O(N__40237),
            .I(N__40233));
    CascadeMux I__8078 (
            .O(N__40236),
            .I(N__40230));
    LocalMux I__8077 (
            .O(N__40233),
            .I(N__40227));
    InMux I__8076 (
            .O(N__40230),
            .I(N__40223));
    Span4Mux_h I__8075 (
            .O(N__40227),
            .I(N__40220));
    InMux I__8074 (
            .O(N__40226),
            .I(N__40217));
    LocalMux I__8073 (
            .O(N__40223),
            .I(N__40214));
    Span4Mux_v I__8072 (
            .O(N__40220),
            .I(N__40211));
    LocalMux I__8071 (
            .O(N__40217),
            .I(buf_dds0_8));
    Odrv4 I__8070 (
            .O(N__40214),
            .I(buf_dds0_8));
    Odrv4 I__8069 (
            .O(N__40211),
            .I(buf_dds0_8));
    InMux I__8068 (
            .O(N__40204),
            .I(N__40200));
    InMux I__8067 (
            .O(N__40203),
            .I(N__40197));
    LocalMux I__8066 (
            .O(N__40200),
            .I(N__40191));
    LocalMux I__8065 (
            .O(N__40197),
            .I(N__40191));
    InMux I__8064 (
            .O(N__40196),
            .I(N__40188));
    Span4Mux_h I__8063 (
            .O(N__40191),
            .I(N__40185));
    LocalMux I__8062 (
            .O(N__40188),
            .I(data_index_1));
    Odrv4 I__8061 (
            .O(N__40185),
            .I(data_index_1));
    InMux I__8060 (
            .O(N__40180),
            .I(N__40177));
    LocalMux I__8059 (
            .O(N__40177),
            .I(n8_adj_1630));
    CascadeMux I__8058 (
            .O(N__40174),
            .I(n8_adj_1630_cascade_));
    InMux I__8057 (
            .O(N__40171),
            .I(N__40165));
    InMux I__8056 (
            .O(N__40170),
            .I(N__40165));
    LocalMux I__8055 (
            .O(N__40165),
            .I(N__40162));
    Odrv12 I__8054 (
            .O(N__40162),
            .I(n7_adj_1629));
    CascadeMux I__8053 (
            .O(N__40159),
            .I(N__40156));
    CascadeBuf I__8052 (
            .O(N__40156),
            .I(N__40153));
    CascadeMux I__8051 (
            .O(N__40153),
            .I(N__40150));
    CascadeBuf I__8050 (
            .O(N__40150),
            .I(N__40147));
    CascadeMux I__8049 (
            .O(N__40147),
            .I(N__40144));
    CascadeBuf I__8048 (
            .O(N__40144),
            .I(N__40141));
    CascadeMux I__8047 (
            .O(N__40141),
            .I(N__40138));
    CascadeBuf I__8046 (
            .O(N__40138),
            .I(N__40135));
    CascadeMux I__8045 (
            .O(N__40135),
            .I(N__40132));
    CascadeBuf I__8044 (
            .O(N__40132),
            .I(N__40129));
    CascadeMux I__8043 (
            .O(N__40129),
            .I(N__40126));
    CascadeBuf I__8042 (
            .O(N__40126),
            .I(N__40123));
    CascadeMux I__8041 (
            .O(N__40123),
            .I(N__40120));
    CascadeBuf I__8040 (
            .O(N__40120),
            .I(N__40116));
    CascadeMux I__8039 (
            .O(N__40119),
            .I(N__40113));
    CascadeMux I__8038 (
            .O(N__40116),
            .I(N__40110));
    CascadeBuf I__8037 (
            .O(N__40113),
            .I(N__40107));
    CascadeBuf I__8036 (
            .O(N__40110),
            .I(N__40104));
    CascadeMux I__8035 (
            .O(N__40107),
            .I(N__40101));
    CascadeMux I__8034 (
            .O(N__40104),
            .I(N__40098));
    InMux I__8033 (
            .O(N__40101),
            .I(N__40095));
    CascadeBuf I__8032 (
            .O(N__40098),
            .I(N__40092));
    LocalMux I__8031 (
            .O(N__40095),
            .I(N__40089));
    CascadeMux I__8030 (
            .O(N__40092),
            .I(N__40086));
    Sp12to4 I__8029 (
            .O(N__40089),
            .I(N__40083));
    InMux I__8028 (
            .O(N__40086),
            .I(N__40080));
    Span12Mux_v I__8027 (
            .O(N__40083),
            .I(N__40077));
    LocalMux I__8026 (
            .O(N__40080),
            .I(N__40074));
    Odrv12 I__8025 (
            .O(N__40077),
            .I(data_index_9_N_236_1));
    Odrv12 I__8024 (
            .O(N__40074),
            .I(data_index_9_N_236_1));
    InMux I__8023 (
            .O(N__40069),
            .I(N__40066));
    LocalMux I__8022 (
            .O(N__40066),
            .I(N__40061));
    InMux I__8021 (
            .O(N__40065),
            .I(N__40058));
    InMux I__8020 (
            .O(N__40064),
            .I(N__40055));
    Span4Mux_v I__8019 (
            .O(N__40061),
            .I(N__40052));
    LocalMux I__8018 (
            .O(N__40058),
            .I(buf_dds0_3));
    LocalMux I__8017 (
            .O(N__40055),
            .I(buf_dds0_3));
    Odrv4 I__8016 (
            .O(N__40052),
            .I(buf_dds0_3));
    InMux I__8015 (
            .O(N__40045),
            .I(N__40041));
    CascadeMux I__8014 (
            .O(N__40044),
            .I(N__40038));
    LocalMux I__8013 (
            .O(N__40041),
            .I(N__40035));
    InMux I__8012 (
            .O(N__40038),
            .I(N__40032));
    Span4Mux_v I__8011 (
            .O(N__40035),
            .I(N__40027));
    LocalMux I__8010 (
            .O(N__40032),
            .I(N__40027));
    Odrv4 I__8009 (
            .O(N__40027),
            .I(tmp_buf_15));
    IoInMux I__8008 (
            .O(N__40024),
            .I(N__40021));
    LocalMux I__8007 (
            .O(N__40021),
            .I(N__40018));
    Span4Mux_s2_v I__8006 (
            .O(N__40018),
            .I(N__40015));
    Span4Mux_v I__8005 (
            .O(N__40015),
            .I(N__40012));
    Sp12to4 I__8004 (
            .O(N__40012),
            .I(N__40008));
    InMux I__8003 (
            .O(N__40011),
            .I(N__40005));
    Odrv12 I__8002 (
            .O(N__40008),
            .I(DDS_MOSI));
    LocalMux I__8001 (
            .O(N__40005),
            .I(DDS_MOSI));
    InMux I__8000 (
            .O(N__40000),
            .I(N__39997));
    LocalMux I__7999 (
            .O(N__39997),
            .I(\comm_spi.n24016 ));
    InMux I__7998 (
            .O(N__39994),
            .I(N__39991));
    LocalMux I__7997 (
            .O(N__39991),
            .I(\comm_spi.n15326 ));
    CascadeMux I__7996 (
            .O(N__39988),
            .I(\comm_spi.n24016_cascade_ ));
    CascadeMux I__7995 (
            .O(N__39985),
            .I(n14_adj_1610_cascade_));
    CascadeMux I__7994 (
            .O(N__39982),
            .I(N__39978));
    InMux I__7993 (
            .O(N__39981),
            .I(N__39975));
    InMux I__7992 (
            .O(N__39978),
            .I(N__39972));
    LocalMux I__7991 (
            .O(N__39975),
            .I(N__39969));
    LocalMux I__7990 (
            .O(N__39972),
            .I(acadc_skipcnt_0));
    Odrv4 I__7989 (
            .O(N__39969),
            .I(acadc_skipcnt_0));
    CascadeMux I__7988 (
            .O(N__39964),
            .I(N__39961));
    InMux I__7987 (
            .O(N__39961),
            .I(N__39958));
    LocalMux I__7986 (
            .O(N__39958),
            .I(N__39954));
    InMux I__7985 (
            .O(N__39957),
            .I(N__39951));
    Span4Mux_h I__7984 (
            .O(N__39954),
            .I(N__39948));
    LocalMux I__7983 (
            .O(N__39951),
            .I(acadc_skipcnt_6));
    Odrv4 I__7982 (
            .O(N__39948),
            .I(acadc_skipcnt_6));
    IoInMux I__7981 (
            .O(N__39943),
            .I(N__39940));
    LocalMux I__7980 (
            .O(N__39940),
            .I(N__39937));
    Span4Mux_s0_v I__7979 (
            .O(N__39937),
            .I(N__39934));
    Span4Mux_v I__7978 (
            .O(N__39934),
            .I(N__39931));
    Span4Mux_v I__7977 (
            .O(N__39931),
            .I(N__39928));
    Sp12to4 I__7976 (
            .O(N__39928),
            .I(N__39923));
    InMux I__7975 (
            .O(N__39927),
            .I(N__39920));
    InMux I__7974 (
            .O(N__39926),
            .I(N__39917));
    Odrv12 I__7973 (
            .O(N__39923),
            .I(SELIRNG0));
    LocalMux I__7972 (
            .O(N__39920),
            .I(SELIRNG0));
    LocalMux I__7971 (
            .O(N__39917),
            .I(SELIRNG0));
    InMux I__7970 (
            .O(N__39910),
            .I(N__39905));
    InMux I__7969 (
            .O(N__39909),
            .I(N__39902));
    InMux I__7968 (
            .O(N__39908),
            .I(N__39899));
    LocalMux I__7967 (
            .O(N__39905),
            .I(acadc_skipCount_10));
    LocalMux I__7966 (
            .O(N__39902),
            .I(acadc_skipCount_10));
    LocalMux I__7965 (
            .O(N__39899),
            .I(acadc_skipCount_10));
    IoInMux I__7964 (
            .O(N__39892),
            .I(N__39889));
    LocalMux I__7963 (
            .O(N__39889),
            .I(N__39886));
    Span4Mux_s0_h I__7962 (
            .O(N__39886),
            .I(N__39883));
    Sp12to4 I__7961 (
            .O(N__39883),
            .I(N__39880));
    Span12Mux_v I__7960 (
            .O(N__39880),
            .I(N__39876));
    CascadeMux I__7959 (
            .O(N__39879),
            .I(N__39872));
    Span12Mux_h I__7958 (
            .O(N__39876),
            .I(N__39869));
    InMux I__7957 (
            .O(N__39875),
            .I(N__39866));
    InMux I__7956 (
            .O(N__39872),
            .I(N__39863));
    Odrv12 I__7955 (
            .O(N__39869),
            .I(VDC_RNG0));
    LocalMux I__7954 (
            .O(N__39866),
            .I(VDC_RNG0));
    LocalMux I__7953 (
            .O(N__39863),
            .I(VDC_RNG0));
    CascadeMux I__7952 (
            .O(N__39856),
            .I(N__39851));
    CascadeMux I__7951 (
            .O(N__39855),
            .I(N__39848));
    InMux I__7950 (
            .O(N__39854),
            .I(N__39845));
    InMux I__7949 (
            .O(N__39851),
            .I(N__39840));
    InMux I__7948 (
            .O(N__39848),
            .I(N__39840));
    LocalMux I__7947 (
            .O(N__39845),
            .I(acadc_skipCount_12));
    LocalMux I__7946 (
            .O(N__39840),
            .I(acadc_skipCount_12));
    InMux I__7945 (
            .O(N__39835),
            .I(N__39832));
    LocalMux I__7944 (
            .O(N__39832),
            .I(N__39829));
    Span4Mux_v I__7943 (
            .O(N__39829),
            .I(N__39826));
    Span4Mux_h I__7942 (
            .O(N__39826),
            .I(N__39823));
    Odrv4 I__7941 (
            .O(N__39823),
            .I(n23_adj_1783));
    CascadeMux I__7940 (
            .O(N__39820),
            .I(N__39813));
    InMux I__7939 (
            .O(N__39819),
            .I(N__39801));
    InMux I__7938 (
            .O(N__39818),
            .I(N__39801));
    InMux I__7937 (
            .O(N__39817),
            .I(N__39794));
    InMux I__7936 (
            .O(N__39816),
            .I(N__39785));
    InMux I__7935 (
            .O(N__39813),
            .I(N__39785));
    InMux I__7934 (
            .O(N__39812),
            .I(N__39785));
    InMux I__7933 (
            .O(N__39811),
            .I(N__39785));
    InMux I__7932 (
            .O(N__39810),
            .I(N__39782));
    CascadeMux I__7931 (
            .O(N__39809),
            .I(N__39777));
    CascadeMux I__7930 (
            .O(N__39808),
            .I(N__39769));
    CascadeMux I__7929 (
            .O(N__39807),
            .I(N__39759));
    InMux I__7928 (
            .O(N__39806),
            .I(N__39755));
    LocalMux I__7927 (
            .O(N__39801),
            .I(N__39750));
    InMux I__7926 (
            .O(N__39800),
            .I(N__39747));
    InMux I__7925 (
            .O(N__39799),
            .I(N__39738));
    InMux I__7924 (
            .O(N__39798),
            .I(N__39738));
    InMux I__7923 (
            .O(N__39797),
            .I(N__39738));
    LocalMux I__7922 (
            .O(N__39794),
            .I(N__39733));
    LocalMux I__7921 (
            .O(N__39785),
            .I(N__39733));
    LocalMux I__7920 (
            .O(N__39782),
            .I(N__39729));
    InMux I__7919 (
            .O(N__39781),
            .I(N__39725));
    InMux I__7918 (
            .O(N__39780),
            .I(N__39716));
    InMux I__7917 (
            .O(N__39777),
            .I(N__39716));
    InMux I__7916 (
            .O(N__39776),
            .I(N__39716));
    InMux I__7915 (
            .O(N__39775),
            .I(N__39716));
    InMux I__7914 (
            .O(N__39774),
            .I(N__39704));
    InMux I__7913 (
            .O(N__39773),
            .I(N__39704));
    InMux I__7912 (
            .O(N__39772),
            .I(N__39704));
    InMux I__7911 (
            .O(N__39769),
            .I(N__39701));
    InMux I__7910 (
            .O(N__39768),
            .I(N__39690));
    InMux I__7909 (
            .O(N__39767),
            .I(N__39690));
    InMux I__7908 (
            .O(N__39766),
            .I(N__39690));
    InMux I__7907 (
            .O(N__39765),
            .I(N__39690));
    InMux I__7906 (
            .O(N__39764),
            .I(N__39690));
    InMux I__7905 (
            .O(N__39763),
            .I(N__39685));
    InMux I__7904 (
            .O(N__39762),
            .I(N__39685));
    InMux I__7903 (
            .O(N__39759),
            .I(N__39682));
    InMux I__7902 (
            .O(N__39758),
            .I(N__39679));
    LocalMux I__7901 (
            .O(N__39755),
            .I(N__39676));
    InMux I__7900 (
            .O(N__39754),
            .I(N__39672));
    InMux I__7899 (
            .O(N__39753),
            .I(N__39669));
    Span4Mux_v I__7898 (
            .O(N__39750),
            .I(N__39664));
    LocalMux I__7897 (
            .O(N__39747),
            .I(N__39664));
    InMux I__7896 (
            .O(N__39746),
            .I(N__39659));
    InMux I__7895 (
            .O(N__39745),
            .I(N__39659));
    LocalMux I__7894 (
            .O(N__39738),
            .I(N__39656));
    Span4Mux_v I__7893 (
            .O(N__39733),
            .I(N__39653));
    InMux I__7892 (
            .O(N__39732),
            .I(N__39648));
    Span4Mux_h I__7891 (
            .O(N__39729),
            .I(N__39645));
    InMux I__7890 (
            .O(N__39728),
            .I(N__39642));
    LocalMux I__7889 (
            .O(N__39725),
            .I(N__39637));
    LocalMux I__7888 (
            .O(N__39716),
            .I(N__39637));
    CascadeMux I__7887 (
            .O(N__39715),
            .I(N__39633));
    CascadeMux I__7886 (
            .O(N__39714),
            .I(N__39627));
    CascadeMux I__7885 (
            .O(N__39713),
            .I(N__39624));
    CascadeMux I__7884 (
            .O(N__39712),
            .I(N__39614));
    CascadeMux I__7883 (
            .O(N__39711),
            .I(N__39611));
    LocalMux I__7882 (
            .O(N__39704),
            .I(N__39605));
    LocalMux I__7881 (
            .O(N__39701),
            .I(N__39598));
    LocalMux I__7880 (
            .O(N__39690),
            .I(N__39598));
    LocalMux I__7879 (
            .O(N__39685),
            .I(N__39598));
    LocalMux I__7878 (
            .O(N__39682),
            .I(N__39593));
    LocalMux I__7877 (
            .O(N__39679),
            .I(N__39593));
    Span4Mux_v I__7876 (
            .O(N__39676),
            .I(N__39590));
    InMux I__7875 (
            .O(N__39675),
            .I(N__39587));
    LocalMux I__7874 (
            .O(N__39672),
            .I(N__39580));
    LocalMux I__7873 (
            .O(N__39669),
            .I(N__39580));
    Span4Mux_h I__7872 (
            .O(N__39664),
            .I(N__39580));
    LocalMux I__7871 (
            .O(N__39659),
            .I(N__39573));
    Span4Mux_v I__7870 (
            .O(N__39656),
            .I(N__39573));
    Span4Mux_v I__7869 (
            .O(N__39653),
            .I(N__39573));
    InMux I__7868 (
            .O(N__39652),
            .I(N__39568));
    InMux I__7867 (
            .O(N__39651),
            .I(N__39568));
    LocalMux I__7866 (
            .O(N__39648),
            .I(N__39565));
    Span4Mux_h I__7865 (
            .O(N__39645),
            .I(N__39562));
    LocalMux I__7864 (
            .O(N__39642),
            .I(N__39557));
    Span4Mux_v I__7863 (
            .O(N__39637),
            .I(N__39557));
    InMux I__7862 (
            .O(N__39636),
            .I(N__39545));
    InMux I__7861 (
            .O(N__39633),
            .I(N__39542));
    InMux I__7860 (
            .O(N__39632),
            .I(N__39537));
    InMux I__7859 (
            .O(N__39631),
            .I(N__39537));
    InMux I__7858 (
            .O(N__39630),
            .I(N__39534));
    InMux I__7857 (
            .O(N__39627),
            .I(N__39523));
    InMux I__7856 (
            .O(N__39624),
            .I(N__39523));
    InMux I__7855 (
            .O(N__39623),
            .I(N__39523));
    InMux I__7854 (
            .O(N__39622),
            .I(N__39523));
    InMux I__7853 (
            .O(N__39621),
            .I(N__39523));
    InMux I__7852 (
            .O(N__39620),
            .I(N__39520));
    InMux I__7851 (
            .O(N__39619),
            .I(N__39513));
    InMux I__7850 (
            .O(N__39618),
            .I(N__39513));
    InMux I__7849 (
            .O(N__39617),
            .I(N__39513));
    InMux I__7848 (
            .O(N__39614),
            .I(N__39502));
    InMux I__7847 (
            .O(N__39611),
            .I(N__39502));
    InMux I__7846 (
            .O(N__39610),
            .I(N__39502));
    InMux I__7845 (
            .O(N__39609),
            .I(N__39502));
    InMux I__7844 (
            .O(N__39608),
            .I(N__39502));
    Span4Mux_h I__7843 (
            .O(N__39605),
            .I(N__39499));
    Span4Mux_h I__7842 (
            .O(N__39598),
            .I(N__39496));
    Span12Mux_h I__7841 (
            .O(N__39593),
            .I(N__39493));
    Span4Mux_h I__7840 (
            .O(N__39590),
            .I(N__39490));
    LocalMux I__7839 (
            .O(N__39587),
            .I(N__39483));
    Span4Mux_v I__7838 (
            .O(N__39580),
            .I(N__39483));
    Span4Mux_h I__7837 (
            .O(N__39573),
            .I(N__39483));
    LocalMux I__7836 (
            .O(N__39568),
            .I(N__39474));
    Span4Mux_h I__7835 (
            .O(N__39565),
            .I(N__39474));
    Span4Mux_v I__7834 (
            .O(N__39562),
            .I(N__39474));
    Span4Mux_h I__7833 (
            .O(N__39557),
            .I(N__39474));
    InMux I__7832 (
            .O(N__39556),
            .I(N__39465));
    InMux I__7831 (
            .O(N__39555),
            .I(N__39465));
    InMux I__7830 (
            .O(N__39554),
            .I(N__39465));
    InMux I__7829 (
            .O(N__39553),
            .I(N__39465));
    InMux I__7828 (
            .O(N__39552),
            .I(N__39454));
    InMux I__7827 (
            .O(N__39551),
            .I(N__39454));
    InMux I__7826 (
            .O(N__39550),
            .I(N__39454));
    InMux I__7825 (
            .O(N__39549),
            .I(N__39454));
    InMux I__7824 (
            .O(N__39548),
            .I(N__39454));
    LocalMux I__7823 (
            .O(N__39545),
            .I(adc_state_0));
    LocalMux I__7822 (
            .O(N__39542),
            .I(adc_state_0));
    LocalMux I__7821 (
            .O(N__39537),
            .I(adc_state_0));
    LocalMux I__7820 (
            .O(N__39534),
            .I(adc_state_0));
    LocalMux I__7819 (
            .O(N__39523),
            .I(adc_state_0));
    LocalMux I__7818 (
            .O(N__39520),
            .I(adc_state_0));
    LocalMux I__7817 (
            .O(N__39513),
            .I(adc_state_0));
    LocalMux I__7816 (
            .O(N__39502),
            .I(adc_state_0));
    Odrv4 I__7815 (
            .O(N__39499),
            .I(adc_state_0));
    Odrv4 I__7814 (
            .O(N__39496),
            .I(adc_state_0));
    Odrv12 I__7813 (
            .O(N__39493),
            .I(adc_state_0));
    Odrv4 I__7812 (
            .O(N__39490),
            .I(adc_state_0));
    Odrv4 I__7811 (
            .O(N__39483),
            .I(adc_state_0));
    Odrv4 I__7810 (
            .O(N__39474),
            .I(adc_state_0));
    LocalMux I__7809 (
            .O(N__39465),
            .I(adc_state_0));
    LocalMux I__7808 (
            .O(N__39454),
            .I(adc_state_0));
    InMux I__7807 (
            .O(N__39421),
            .I(N__39415));
    InMux I__7806 (
            .O(N__39420),
            .I(N__39410));
    InMux I__7805 (
            .O(N__39419),
            .I(N__39410));
    CascadeMux I__7804 (
            .O(N__39418),
            .I(N__39407));
    LocalMux I__7803 (
            .O(N__39415),
            .I(N__39395));
    LocalMux I__7802 (
            .O(N__39410),
            .I(N__39392));
    InMux I__7801 (
            .O(N__39407),
            .I(N__39387));
    InMux I__7800 (
            .O(N__39406),
            .I(N__39387));
    InMux I__7799 (
            .O(N__39405),
            .I(N__39382));
    InMux I__7798 (
            .O(N__39404),
            .I(N__39379));
    InMux I__7797 (
            .O(N__39403),
            .I(N__39372));
    InMux I__7796 (
            .O(N__39402),
            .I(N__39372));
    InMux I__7795 (
            .O(N__39401),
            .I(N__39365));
    InMux I__7794 (
            .O(N__39400),
            .I(N__39365));
    InMux I__7793 (
            .O(N__39399),
            .I(N__39362));
    InMux I__7792 (
            .O(N__39398),
            .I(N__39357));
    Span4Mux_v I__7791 (
            .O(N__39395),
            .I(N__39352));
    Span4Mux_h I__7790 (
            .O(N__39392),
            .I(N__39352));
    LocalMux I__7789 (
            .O(N__39387),
            .I(N__39348));
    InMux I__7788 (
            .O(N__39386),
            .I(N__39345));
    InMux I__7787 (
            .O(N__39385),
            .I(N__39342));
    LocalMux I__7786 (
            .O(N__39382),
            .I(N__39338));
    LocalMux I__7785 (
            .O(N__39379),
            .I(N__39335));
    InMux I__7784 (
            .O(N__39378),
            .I(N__39329));
    InMux I__7783 (
            .O(N__39377),
            .I(N__39329));
    LocalMux I__7782 (
            .O(N__39372),
            .I(N__39326));
    InMux I__7781 (
            .O(N__39371),
            .I(N__39321));
    InMux I__7780 (
            .O(N__39370),
            .I(N__39321));
    LocalMux I__7779 (
            .O(N__39365),
            .I(N__39318));
    LocalMux I__7778 (
            .O(N__39362),
            .I(N__39315));
    InMux I__7777 (
            .O(N__39361),
            .I(N__39310));
    InMux I__7776 (
            .O(N__39360),
            .I(N__39310));
    LocalMux I__7775 (
            .O(N__39357),
            .I(N__39305));
    Span4Mux_v I__7774 (
            .O(N__39352),
            .I(N__39305));
    InMux I__7773 (
            .O(N__39351),
            .I(N__39302));
    Span4Mux_h I__7772 (
            .O(N__39348),
            .I(N__39297));
    LocalMux I__7771 (
            .O(N__39345),
            .I(N__39297));
    LocalMux I__7770 (
            .O(N__39342),
            .I(N__39294));
    InMux I__7769 (
            .O(N__39341),
            .I(N__39291));
    Span4Mux_h I__7768 (
            .O(N__39338),
            .I(N__39286));
    Span4Mux_v I__7767 (
            .O(N__39335),
            .I(N__39286));
    InMux I__7766 (
            .O(N__39334),
            .I(N__39283));
    LocalMux I__7765 (
            .O(N__39329),
            .I(N__39274));
    Span4Mux_v I__7764 (
            .O(N__39326),
            .I(N__39274));
    LocalMux I__7763 (
            .O(N__39321),
            .I(N__39274));
    Span4Mux_v I__7762 (
            .O(N__39318),
            .I(N__39274));
    Span4Mux_h I__7761 (
            .O(N__39315),
            .I(N__39271));
    LocalMux I__7760 (
            .O(N__39310),
            .I(N__39266));
    Span4Mux_v I__7759 (
            .O(N__39305),
            .I(N__39266));
    LocalMux I__7758 (
            .O(N__39302),
            .I(N__39263));
    Span4Mux_v I__7757 (
            .O(N__39297),
            .I(N__39260));
    Span4Mux_h I__7756 (
            .O(N__39294),
            .I(N__39257));
    LocalMux I__7755 (
            .O(N__39291),
            .I(N__39252));
    Span4Mux_v I__7754 (
            .O(N__39286),
            .I(N__39252));
    LocalMux I__7753 (
            .O(N__39283),
            .I(N__39249));
    Span4Mux_h I__7752 (
            .O(N__39274),
            .I(N__39246));
    Span4Mux_v I__7751 (
            .O(N__39271),
            .I(N__39241));
    Span4Mux_h I__7750 (
            .O(N__39266),
            .I(N__39241));
    Span4Mux_h I__7749 (
            .O(N__39263),
            .I(N__39232));
    Span4Mux_h I__7748 (
            .O(N__39260),
            .I(N__39232));
    Span4Mux_h I__7747 (
            .O(N__39257),
            .I(N__39232));
    Span4Mux_h I__7746 (
            .O(N__39252),
            .I(N__39232));
    Odrv4 I__7745 (
            .O(N__39249),
            .I(n21951));
    Odrv4 I__7744 (
            .O(N__39246),
            .I(n21951));
    Odrv4 I__7743 (
            .O(N__39241),
            .I(n21951));
    Odrv4 I__7742 (
            .O(N__39232),
            .I(n21951));
    CascadeMux I__7741 (
            .O(N__39223),
            .I(N__39220));
    InMux I__7740 (
            .O(N__39220),
            .I(N__39217));
    LocalMux I__7739 (
            .O(N__39217),
            .I(N__39213));
    CascadeMux I__7738 (
            .O(N__39216),
            .I(N__39210));
    Span12Mux_h I__7737 (
            .O(N__39213),
            .I(N__39206));
    InMux I__7736 (
            .O(N__39210),
            .I(N__39201));
    InMux I__7735 (
            .O(N__39209),
            .I(N__39201));
    Odrv12 I__7734 (
            .O(N__39206),
            .I(cmd_rdadctmp_17));
    LocalMux I__7733 (
            .O(N__39201),
            .I(cmd_rdadctmp_17));
    InMux I__7732 (
            .O(N__39196),
            .I(N__39193));
    LocalMux I__7731 (
            .O(N__39193),
            .I(N__39188));
    InMux I__7730 (
            .O(N__39192),
            .I(N__39183));
    InMux I__7729 (
            .O(N__39191),
            .I(N__39183));
    Odrv4 I__7728 (
            .O(N__39188),
            .I(req_data_cnt_10));
    LocalMux I__7727 (
            .O(N__39183),
            .I(req_data_cnt_10));
    SRMux I__7726 (
            .O(N__39178),
            .I(N__39174));
    InMux I__7725 (
            .O(N__39177),
            .I(N__39167));
    LocalMux I__7724 (
            .O(N__39174),
            .I(N__39164));
    InMux I__7723 (
            .O(N__39173),
            .I(N__39161));
    SRMux I__7722 (
            .O(N__39172),
            .I(N__39158));
    InMux I__7721 (
            .O(N__39171),
            .I(N__39155));
    InMux I__7720 (
            .O(N__39170),
            .I(N__39152));
    LocalMux I__7719 (
            .O(N__39167),
            .I(N__39149));
    Span4Mux_v I__7718 (
            .O(N__39164),
            .I(N__39145));
    LocalMux I__7717 (
            .O(N__39161),
            .I(N__39142));
    LocalMux I__7716 (
            .O(N__39158),
            .I(N__39137));
    LocalMux I__7715 (
            .O(N__39155),
            .I(N__39137));
    LocalMux I__7714 (
            .O(N__39152),
            .I(N__39134));
    Span12Mux_s10_v I__7713 (
            .O(N__39149),
            .I(N__39127));
    InMux I__7712 (
            .O(N__39148),
            .I(N__39124));
    Span4Mux_h I__7711 (
            .O(N__39145),
            .I(N__39119));
    Span4Mux_v I__7710 (
            .O(N__39142),
            .I(N__39119));
    Span4Mux_h I__7709 (
            .O(N__39137),
            .I(N__39116));
    Span12Mux_h I__7708 (
            .O(N__39134),
            .I(N__39113));
    InMux I__7707 (
            .O(N__39133),
            .I(N__39110));
    InMux I__7706 (
            .O(N__39132),
            .I(N__39105));
    InMux I__7705 (
            .O(N__39131),
            .I(N__39105));
    InMux I__7704 (
            .O(N__39130),
            .I(N__39102));
    Odrv12 I__7703 (
            .O(N__39127),
            .I(acadc_rst));
    LocalMux I__7702 (
            .O(N__39124),
            .I(acadc_rst));
    Odrv4 I__7701 (
            .O(N__39119),
            .I(acadc_rst));
    Odrv4 I__7700 (
            .O(N__39116),
            .I(acadc_rst));
    Odrv12 I__7699 (
            .O(N__39113),
            .I(acadc_rst));
    LocalMux I__7698 (
            .O(N__39110),
            .I(acadc_rst));
    LocalMux I__7697 (
            .O(N__39105),
            .I(acadc_rst));
    LocalMux I__7696 (
            .O(N__39102),
            .I(acadc_rst));
    CascadeMux I__7695 (
            .O(N__39085),
            .I(N__39082));
    CascadeBuf I__7694 (
            .O(N__39082),
            .I(N__39079));
    CascadeMux I__7693 (
            .O(N__39079),
            .I(N__39076));
    CascadeBuf I__7692 (
            .O(N__39076),
            .I(N__39073));
    CascadeMux I__7691 (
            .O(N__39073),
            .I(N__39070));
    CascadeBuf I__7690 (
            .O(N__39070),
            .I(N__39067));
    CascadeMux I__7689 (
            .O(N__39067),
            .I(N__39064));
    CascadeBuf I__7688 (
            .O(N__39064),
            .I(N__39061));
    CascadeMux I__7687 (
            .O(N__39061),
            .I(N__39058));
    CascadeBuf I__7686 (
            .O(N__39058),
            .I(N__39055));
    CascadeMux I__7685 (
            .O(N__39055),
            .I(N__39052));
    CascadeBuf I__7684 (
            .O(N__39052),
            .I(N__39049));
    CascadeMux I__7683 (
            .O(N__39049),
            .I(N__39046));
    CascadeBuf I__7682 (
            .O(N__39046),
            .I(N__39042));
    CascadeMux I__7681 (
            .O(N__39045),
            .I(N__39039));
    CascadeMux I__7680 (
            .O(N__39042),
            .I(N__39036));
    CascadeBuf I__7679 (
            .O(N__39039),
            .I(N__39033));
    CascadeBuf I__7678 (
            .O(N__39036),
            .I(N__39030));
    CascadeMux I__7677 (
            .O(N__39033),
            .I(N__39027));
    CascadeMux I__7676 (
            .O(N__39030),
            .I(N__39024));
    InMux I__7675 (
            .O(N__39027),
            .I(N__39021));
    CascadeBuf I__7674 (
            .O(N__39024),
            .I(N__39018));
    LocalMux I__7673 (
            .O(N__39021),
            .I(N__39015));
    CascadeMux I__7672 (
            .O(N__39018),
            .I(N__39012));
    Span4Mux_v I__7671 (
            .O(N__39015),
            .I(N__39009));
    InMux I__7670 (
            .O(N__39012),
            .I(N__39006));
    Span4Mux_v I__7669 (
            .O(N__39009),
            .I(N__39003));
    LocalMux I__7668 (
            .O(N__39006),
            .I(N__39000));
    Span4Mux_h I__7667 (
            .O(N__39003),
            .I(N__38997));
    Span4Mux_v I__7666 (
            .O(N__39000),
            .I(N__38994));
    Span4Mux_h I__7665 (
            .O(N__38997),
            .I(N__38991));
    Span4Mux_h I__7664 (
            .O(N__38994),
            .I(N__38988));
    Odrv4 I__7663 (
            .O(N__38991),
            .I(data_index_9_N_236_3));
    Odrv4 I__7662 (
            .O(N__38988),
            .I(data_index_9_N_236_3));
    InMux I__7661 (
            .O(N__38983),
            .I(N__38980));
    LocalMux I__7660 (
            .O(N__38980),
            .I(N__38976));
    InMux I__7659 (
            .O(N__38979),
            .I(N__38973));
    Span4Mux_h I__7658 (
            .O(N__38976),
            .I(N__38970));
    LocalMux I__7657 (
            .O(N__38973),
            .I(acadc_skipcnt_7));
    Odrv4 I__7656 (
            .O(N__38970),
            .I(acadc_skipcnt_7));
    InMux I__7655 (
            .O(N__38965),
            .I(N__38962));
    LocalMux I__7654 (
            .O(N__38962),
            .I(N__38958));
    InMux I__7653 (
            .O(N__38961),
            .I(N__38955));
    Span4Mux_h I__7652 (
            .O(N__38958),
            .I(N__38952));
    LocalMux I__7651 (
            .O(N__38955),
            .I(acadc_skipcnt_2));
    Odrv4 I__7650 (
            .O(N__38952),
            .I(acadc_skipcnt_2));
    InMux I__7649 (
            .O(N__38947),
            .I(N__38944));
    LocalMux I__7648 (
            .O(N__38944),
            .I(N__38940));
    InMux I__7647 (
            .O(N__38943),
            .I(N__38937));
    Span4Mux_h I__7646 (
            .O(N__38940),
            .I(N__38934));
    LocalMux I__7645 (
            .O(N__38937),
            .I(acadc_skipcnt_12));
    Odrv4 I__7644 (
            .O(N__38934),
            .I(acadc_skipcnt_12));
    InMux I__7643 (
            .O(N__38929),
            .I(N__38926));
    LocalMux I__7642 (
            .O(N__38926),
            .I(N__38922));
    InMux I__7641 (
            .O(N__38925),
            .I(N__38919));
    Span4Mux_h I__7640 (
            .O(N__38922),
            .I(N__38916));
    LocalMux I__7639 (
            .O(N__38919),
            .I(acadc_skipcnt_10));
    Odrv4 I__7638 (
            .O(N__38916),
            .I(acadc_skipcnt_10));
    InMux I__7637 (
            .O(N__38911),
            .I(N__38908));
    LocalMux I__7636 (
            .O(N__38908),
            .I(N__38905));
    Odrv4 I__7635 (
            .O(N__38905),
            .I(n23_adj_1514));
    InMux I__7634 (
            .O(N__38902),
            .I(N__38899));
    LocalMux I__7633 (
            .O(N__38899),
            .I(n24_adj_1513));
    CascadeMux I__7632 (
            .O(N__38896),
            .I(n21_cascade_));
    InMux I__7631 (
            .O(N__38893),
            .I(N__38890));
    LocalMux I__7630 (
            .O(N__38890),
            .I(n22));
    InMux I__7629 (
            .O(N__38887),
            .I(n20656));
    InMux I__7628 (
            .O(N__38884),
            .I(n20657));
    InMux I__7627 (
            .O(N__38881),
            .I(n20658));
    InMux I__7626 (
            .O(N__38878),
            .I(bfn_13_16_0_));
    InMux I__7625 (
            .O(N__38875),
            .I(n20660));
    InMux I__7624 (
            .O(N__38872),
            .I(N__38868));
    InMux I__7623 (
            .O(N__38871),
            .I(N__38863));
    LocalMux I__7622 (
            .O(N__38868),
            .I(N__38860));
    InMux I__7621 (
            .O(N__38867),
            .I(N__38857));
    InMux I__7620 (
            .O(N__38866),
            .I(N__38854));
    LocalMux I__7619 (
            .O(N__38863),
            .I(N__38851));
    Span4Mux_v I__7618 (
            .O(N__38860),
            .I(N__38846));
    LocalMux I__7617 (
            .O(N__38857),
            .I(N__38846));
    LocalMux I__7616 (
            .O(N__38854),
            .I(eis_stop));
    Odrv4 I__7615 (
            .O(N__38851),
            .I(eis_stop));
    Odrv4 I__7614 (
            .O(N__38846),
            .I(eis_stop));
    InMux I__7613 (
            .O(N__38839),
            .I(N__38836));
    LocalMux I__7612 (
            .O(N__38836),
            .I(N__38832));
    InMux I__7611 (
            .O(N__38835),
            .I(N__38829));
    Span4Mux_h I__7610 (
            .O(N__38832),
            .I(N__38826));
    LocalMux I__7609 (
            .O(N__38829),
            .I(acadc_skipcnt_13));
    Odrv4 I__7608 (
            .O(N__38826),
            .I(acadc_skipcnt_13));
    InMux I__7607 (
            .O(N__38821),
            .I(N__38818));
    LocalMux I__7606 (
            .O(N__38818),
            .I(N__38813));
    InMux I__7605 (
            .O(N__38817),
            .I(N__38808));
    InMux I__7604 (
            .O(N__38816),
            .I(N__38808));
    Odrv4 I__7603 (
            .O(N__38813),
            .I(acadc_skipCount_13));
    LocalMux I__7602 (
            .O(N__38808),
            .I(acadc_skipCount_13));
    IoInMux I__7601 (
            .O(N__38803),
            .I(N__38800));
    LocalMux I__7600 (
            .O(N__38800),
            .I(N__38797));
    Span12Mux_s3_h I__7599 (
            .O(N__38797),
            .I(N__38794));
    Span12Mux_h I__7598 (
            .O(N__38794),
            .I(N__38789));
    InMux I__7597 (
            .O(N__38793),
            .I(N__38786));
    InMux I__7596 (
            .O(N__38792),
            .I(N__38783));
    Odrv12 I__7595 (
            .O(N__38789),
            .I(VAC_OSR0));
    LocalMux I__7594 (
            .O(N__38786),
            .I(VAC_OSR0));
    LocalMux I__7593 (
            .O(N__38783),
            .I(VAC_OSR0));
    CascadeMux I__7592 (
            .O(N__38776),
            .I(N__38769));
    CascadeMux I__7591 (
            .O(N__38775),
            .I(N__38766));
    CascadeMux I__7590 (
            .O(N__38774),
            .I(N__38763));
    CascadeMux I__7589 (
            .O(N__38773),
            .I(N__38760));
    CascadeMux I__7588 (
            .O(N__38772),
            .I(N__38754));
    InMux I__7587 (
            .O(N__38769),
            .I(N__38747));
    InMux I__7586 (
            .O(N__38766),
            .I(N__38747));
    InMux I__7585 (
            .O(N__38763),
            .I(N__38747));
    InMux I__7584 (
            .O(N__38760),
            .I(N__38744));
    CascadeMux I__7583 (
            .O(N__38759),
            .I(N__38741));
    CascadeMux I__7582 (
            .O(N__38758),
            .I(N__38738));
    InMux I__7581 (
            .O(N__38757),
            .I(N__38733));
    InMux I__7580 (
            .O(N__38754),
            .I(N__38733));
    LocalMux I__7579 (
            .O(N__38747),
            .I(N__38730));
    LocalMux I__7578 (
            .O(N__38744),
            .I(N__38727));
    InMux I__7577 (
            .O(N__38741),
            .I(N__38722));
    InMux I__7576 (
            .O(N__38738),
            .I(N__38722));
    LocalMux I__7575 (
            .O(N__38733),
            .I(N__38719));
    Span4Mux_h I__7574 (
            .O(N__38730),
            .I(N__38712));
    Span4Mux_h I__7573 (
            .O(N__38727),
            .I(N__38712));
    LocalMux I__7572 (
            .O(N__38722),
            .I(N__38712));
    Odrv4 I__7571 (
            .O(N__38719),
            .I(n40));
    Odrv4 I__7570 (
            .O(N__38712),
            .I(n40));
    InMux I__7569 (
            .O(N__38707),
            .I(N__38704));
    LocalMux I__7568 (
            .O(N__38704),
            .I(N__38701));
    Odrv4 I__7567 (
            .O(N__38701),
            .I(n24_adj_1505));
    InMux I__7566 (
            .O(N__38698),
            .I(N__38695));
    LocalMux I__7565 (
            .O(N__38695),
            .I(N__38691));
    InMux I__7564 (
            .O(N__38694),
            .I(N__38687));
    Span4Mux_h I__7563 (
            .O(N__38691),
            .I(N__38684));
    CascadeMux I__7562 (
            .O(N__38690),
            .I(N__38681));
    LocalMux I__7561 (
            .O(N__38687),
            .I(N__38676));
    Span4Mux_h I__7560 (
            .O(N__38684),
            .I(N__38676));
    InMux I__7559 (
            .O(N__38681),
            .I(N__38673));
    Odrv4 I__7558 (
            .O(N__38676),
            .I(req_data_cnt_12));
    LocalMux I__7557 (
            .O(N__38673),
            .I(req_data_cnt_12));
    IoInMux I__7556 (
            .O(N__38668),
            .I(N__38665));
    LocalMux I__7555 (
            .O(N__38665),
            .I(N__38662));
    Span4Mux_s2_h I__7554 (
            .O(N__38662),
            .I(N__38658));
    InMux I__7553 (
            .O(N__38661),
            .I(N__38654));
    Sp12to4 I__7552 (
            .O(N__38658),
            .I(N__38651));
    InMux I__7551 (
            .O(N__38657),
            .I(N__38648));
    LocalMux I__7550 (
            .O(N__38654),
            .I(N__38645));
    Span12Mux_v I__7549 (
            .O(N__38651),
            .I(N__38642));
    LocalMux I__7548 (
            .O(N__38648),
            .I(N__38639));
    Span4Mux_v I__7547 (
            .O(N__38645),
            .I(N__38636));
    Span12Mux_h I__7546 (
            .O(N__38642),
            .I(N__38633));
    Span4Mux_h I__7545 (
            .O(N__38639),
            .I(N__38628));
    Span4Mux_h I__7544 (
            .O(N__38636),
            .I(N__38628));
    Odrv12 I__7543 (
            .O(N__38633),
            .I(VAC_OSR1));
    Odrv4 I__7542 (
            .O(N__38628),
            .I(VAC_OSR1));
    InMux I__7541 (
            .O(N__38623),
            .I(N__38620));
    LocalMux I__7540 (
            .O(N__38620),
            .I(N__38616));
    CascadeMux I__7539 (
            .O(N__38619),
            .I(N__38613));
    Span4Mux_v I__7538 (
            .O(N__38616),
            .I(N__38610));
    InMux I__7537 (
            .O(N__38613),
            .I(N__38607));
    Sp12to4 I__7536 (
            .O(N__38610),
            .I(N__38603));
    LocalMux I__7535 (
            .O(N__38607),
            .I(N__38600));
    InMux I__7534 (
            .O(N__38606),
            .I(N__38597));
    Span12Mux_h I__7533 (
            .O(N__38603),
            .I(N__38594));
    Span4Mux_h I__7532 (
            .O(N__38600),
            .I(N__38591));
    LocalMux I__7531 (
            .O(N__38597),
            .I(buf_adcdata_iac_21));
    Odrv12 I__7530 (
            .O(N__38594),
            .I(buf_adcdata_iac_21));
    Odrv4 I__7529 (
            .O(N__38591),
            .I(buf_adcdata_iac_21));
    InMux I__7528 (
            .O(N__38584),
            .I(N__38579));
    InMux I__7527 (
            .O(N__38583),
            .I(N__38576));
    InMux I__7526 (
            .O(N__38582),
            .I(N__38573));
    LocalMux I__7525 (
            .O(N__38579),
            .I(N__38570));
    LocalMux I__7524 (
            .O(N__38576),
            .I(N__38565));
    LocalMux I__7523 (
            .O(N__38573),
            .I(N__38565));
    Odrv12 I__7522 (
            .O(N__38570),
            .I(n9_adj_1600));
    Odrv4 I__7521 (
            .O(N__38565),
            .I(n9_adj_1600));
    InMux I__7520 (
            .O(N__38560),
            .I(bfn_13_15_0_));
    InMux I__7519 (
            .O(N__38557),
            .I(n20652));
    InMux I__7518 (
            .O(N__38554),
            .I(n20653));
    InMux I__7517 (
            .O(N__38551),
            .I(n20654));
    InMux I__7516 (
            .O(N__38548),
            .I(n20655));
    CascadeMux I__7515 (
            .O(N__38545),
            .I(n23450_cascade_));
    InMux I__7514 (
            .O(N__38542),
            .I(N__38539));
    LocalMux I__7513 (
            .O(N__38539),
            .I(N__38536));
    Span4Mux_h I__7512 (
            .O(N__38536),
            .I(N__38533));
    Odrv4 I__7511 (
            .O(N__38533),
            .I(n23327));
    InMux I__7510 (
            .O(N__38530),
            .I(N__38527));
    LocalMux I__7509 (
            .O(N__38527),
            .I(N__38524));
    Odrv4 I__7508 (
            .O(N__38524),
            .I(n23453));
    InMux I__7507 (
            .O(N__38521),
            .I(N__38518));
    LocalMux I__7506 (
            .O(N__38518),
            .I(N__38515));
    Odrv4 I__7505 (
            .O(N__38515),
            .I(n112_adj_1583));
    InMux I__7504 (
            .O(N__38512),
            .I(N__38509));
    LocalMux I__7503 (
            .O(N__38509),
            .I(N__38506));
    Span4Mux_v I__7502 (
            .O(N__38506),
            .I(N__38503));
    Odrv4 I__7501 (
            .O(N__38503),
            .I(n23522));
    InMux I__7500 (
            .O(N__38500),
            .I(N__38497));
    LocalMux I__7499 (
            .O(N__38497),
            .I(n22267));
    InMux I__7498 (
            .O(N__38494),
            .I(N__38491));
    LocalMux I__7497 (
            .O(N__38491),
            .I(n112_adj_1797));
    CascadeMux I__7496 (
            .O(N__38488),
            .I(N__38485));
    InMux I__7495 (
            .O(N__38485),
            .I(N__38482));
    LocalMux I__7494 (
            .O(N__38482),
            .I(N__38479));
    Odrv4 I__7493 (
            .O(N__38479),
            .I(comm_buf_0_7_N_543_2));
    InMux I__7492 (
            .O(N__38476),
            .I(N__38473));
    LocalMux I__7491 (
            .O(N__38473),
            .I(N__38469));
    InMux I__7490 (
            .O(N__38472),
            .I(N__38466));
    Span4Mux_h I__7489 (
            .O(N__38469),
            .I(N__38463));
    LocalMux I__7488 (
            .O(N__38466),
            .I(comm_test_buf_24_16));
    Odrv4 I__7487 (
            .O(N__38463),
            .I(comm_test_buf_24_16));
    InMux I__7486 (
            .O(N__38458),
            .I(N__38455));
    LocalMux I__7485 (
            .O(N__38455),
            .I(n111_adj_1584));
    InMux I__7484 (
            .O(N__38452),
            .I(N__38449));
    LocalMux I__7483 (
            .O(N__38449),
            .I(N__38446));
    Odrv4 I__7482 (
            .O(N__38446),
            .I(n20_adj_1804));
    InMux I__7481 (
            .O(N__38443),
            .I(N__38440));
    LocalMux I__7480 (
            .O(N__38440),
            .I(N__38437));
    Span4Mux_v I__7479 (
            .O(N__38437),
            .I(N__38433));
    InMux I__7478 (
            .O(N__38436),
            .I(N__38430));
    Odrv4 I__7477 (
            .O(N__38433),
            .I(\comm_spi.n15338 ));
    LocalMux I__7476 (
            .O(N__38430),
            .I(\comm_spi.n15338 ));
    SRMux I__7475 (
            .O(N__38425),
            .I(N__38422));
    LocalMux I__7474 (
            .O(N__38422),
            .I(N__38419));
    Odrv4 I__7473 (
            .O(N__38419),
            .I(n15496));
    CascadeMux I__7472 (
            .O(N__38416),
            .I(N__38413));
    InMux I__7471 (
            .O(N__38413),
            .I(N__38410));
    LocalMux I__7470 (
            .O(N__38410),
            .I(N__38407));
    Span4Mux_h I__7469 (
            .O(N__38407),
            .I(N__38404));
    Span4Mux_h I__7468 (
            .O(N__38404),
            .I(N__38401));
    Odrv4 I__7467 (
            .O(N__38401),
            .I(buf_data_iac_16));
    CascadeMux I__7466 (
            .O(N__38398),
            .I(n22270_cascade_));
    InMux I__7465 (
            .O(N__38395),
            .I(N__38392));
    LocalMux I__7464 (
            .O(N__38392),
            .I(N__38388));
    InMux I__7463 (
            .O(N__38391),
            .I(N__38385));
    Span4Mux_h I__7462 (
            .O(N__38388),
            .I(N__38382));
    LocalMux I__7461 (
            .O(N__38385),
            .I(comm_test_buf_24_9));
    Odrv4 I__7460 (
            .O(N__38382),
            .I(comm_test_buf_24_9));
    InMux I__7459 (
            .O(N__38377),
            .I(N__38374));
    LocalMux I__7458 (
            .O(N__38374),
            .I(comm_buf_0_7_N_543_0));
    InMux I__7457 (
            .O(N__38371),
            .I(N__38368));
    LocalMux I__7456 (
            .O(N__38368),
            .I(N__38364));
    InMux I__7455 (
            .O(N__38367),
            .I(N__38361));
    Span4Mux_v I__7454 (
            .O(N__38364),
            .I(N__38358));
    LocalMux I__7453 (
            .O(N__38361),
            .I(comm_test_buf_24_18));
    Odrv4 I__7452 (
            .O(N__38358),
            .I(comm_test_buf_24_18));
    InMux I__7451 (
            .O(N__38353),
            .I(N__38348));
    InMux I__7450 (
            .O(N__38352),
            .I(N__38345));
    InMux I__7449 (
            .O(N__38351),
            .I(N__38342));
    LocalMux I__7448 (
            .O(N__38348),
            .I(N__38339));
    LocalMux I__7447 (
            .O(N__38345),
            .I(N__38334));
    LocalMux I__7446 (
            .O(N__38342),
            .I(N__38334));
    Odrv4 I__7445 (
            .O(N__38339),
            .I(comm_test_buf_24_7));
    Odrv4 I__7444 (
            .O(N__38334),
            .I(comm_test_buf_24_7));
    InMux I__7443 (
            .O(N__38329),
            .I(N__38326));
    LocalMux I__7442 (
            .O(N__38326),
            .I(N__38323));
    Span4Mux_h I__7441 (
            .O(N__38323),
            .I(N__38319));
    InMux I__7440 (
            .O(N__38322),
            .I(N__38316));
    Odrv4 I__7439 (
            .O(N__38319),
            .I(comm_test_buf_24_15));
    LocalMux I__7438 (
            .O(N__38316),
            .I(comm_test_buf_24_15));
    InMux I__7437 (
            .O(N__38311),
            .I(N__38308));
    LocalMux I__7436 (
            .O(N__38308),
            .I(N__38304));
    InMux I__7435 (
            .O(N__38307),
            .I(N__38301));
    Span4Mux_h I__7434 (
            .O(N__38304),
            .I(N__38298));
    LocalMux I__7433 (
            .O(N__38301),
            .I(N__38294));
    Span4Mux_v I__7432 (
            .O(N__38298),
            .I(N__38291));
    InMux I__7431 (
            .O(N__38297),
            .I(N__38288));
    Span4Mux_h I__7430 (
            .O(N__38294),
            .I(N__38285));
    Odrv4 I__7429 (
            .O(N__38291),
            .I(comm_buf_2_1));
    LocalMux I__7428 (
            .O(N__38288),
            .I(comm_buf_2_1));
    Odrv4 I__7427 (
            .O(N__38285),
            .I(comm_buf_2_1));
    InMux I__7426 (
            .O(N__38278),
            .I(N__38275));
    LocalMux I__7425 (
            .O(N__38275),
            .I(N__38272));
    Span4Mux_h I__7424 (
            .O(N__38272),
            .I(N__38269));
    Odrv4 I__7423 (
            .O(N__38269),
            .I(n13201));
    InMux I__7422 (
            .O(N__38266),
            .I(N__38263));
    LocalMux I__7421 (
            .O(N__38263),
            .I(N__38260));
    Span4Mux_v I__7420 (
            .O(N__38260),
            .I(N__38257));
    Sp12to4 I__7419 (
            .O(N__38257),
            .I(N__38253));
    InMux I__7418 (
            .O(N__38256),
            .I(N__38250));
    Odrv12 I__7417 (
            .O(N__38253),
            .I(buf_readRTD_9));
    LocalMux I__7416 (
            .O(N__38250),
            .I(buf_readRTD_9));
    CascadeMux I__7415 (
            .O(N__38245),
            .I(N__38242));
    InMux I__7414 (
            .O(N__38242),
            .I(N__38239));
    LocalMux I__7413 (
            .O(N__38239),
            .I(N__38234));
    InMux I__7412 (
            .O(N__38238),
            .I(N__38230));
    InMux I__7411 (
            .O(N__38237),
            .I(N__38227));
    Span4Mux_v I__7410 (
            .O(N__38234),
            .I(N__38224));
    InMux I__7409 (
            .O(N__38233),
            .I(N__38221));
    LocalMux I__7408 (
            .O(N__38230),
            .I(N__38216));
    LocalMux I__7407 (
            .O(N__38227),
            .I(N__38216));
    Span4Mux_h I__7406 (
            .O(N__38224),
            .I(N__38212));
    LocalMux I__7405 (
            .O(N__38221),
            .I(N__38209));
    Span12Mux_v I__7404 (
            .O(N__38216),
            .I(N__38206));
    InMux I__7403 (
            .O(N__38215),
            .I(N__38203));
    Span4Mux_h I__7402 (
            .O(N__38212),
            .I(N__38198));
    Span4Mux_v I__7401 (
            .O(N__38209),
            .I(N__38198));
    Odrv12 I__7400 (
            .O(N__38206),
            .I(buf_cfgRTD_1));
    LocalMux I__7399 (
            .O(N__38203),
            .I(buf_cfgRTD_1));
    Odrv4 I__7398 (
            .O(N__38198),
            .I(buf_cfgRTD_1));
    InMux I__7397 (
            .O(N__38191),
            .I(N__38188));
    LocalMux I__7396 (
            .O(N__38188),
            .I(N__38185));
    Span4Mux_v I__7395 (
            .O(N__38185),
            .I(N__38182));
    Span4Mux_h I__7394 (
            .O(N__38182),
            .I(N__38178));
    InMux I__7393 (
            .O(N__38181),
            .I(N__38175));
    Odrv4 I__7392 (
            .O(N__38178),
            .I(\comm_spi.n15337 ));
    LocalMux I__7391 (
            .O(N__38175),
            .I(\comm_spi.n15337 ));
    CascadeMux I__7390 (
            .O(N__38170),
            .I(N__38167));
    InMux I__7389 (
            .O(N__38167),
            .I(N__38164));
    LocalMux I__7388 (
            .O(N__38164),
            .I(N__38161));
    Span4Mux_v I__7387 (
            .O(N__38161),
            .I(N__38157));
    CascadeMux I__7386 (
            .O(N__38160),
            .I(N__38154));
    Span4Mux_h I__7385 (
            .O(N__38157),
            .I(N__38151));
    InMux I__7384 (
            .O(N__38154),
            .I(N__38148));
    Sp12to4 I__7383 (
            .O(N__38151),
            .I(N__38145));
    LocalMux I__7382 (
            .O(N__38148),
            .I(cmd_rdadctmp_7));
    Odrv12 I__7381 (
            .O(N__38145),
            .I(cmd_rdadctmp_7));
    InMux I__7380 (
            .O(N__38140),
            .I(N__38136));
    InMux I__7379 (
            .O(N__38139),
            .I(N__38133));
    LocalMux I__7378 (
            .O(N__38136),
            .I(comm_buf_6_4));
    LocalMux I__7377 (
            .O(N__38133),
            .I(comm_buf_6_4));
    InMux I__7376 (
            .O(N__38128),
            .I(N__38125));
    LocalMux I__7375 (
            .O(N__38125),
            .I(N__38122));
    Span4Mux_v I__7374 (
            .O(N__38122),
            .I(N__38119));
    Span4Mux_h I__7373 (
            .O(N__38119),
            .I(N__38114));
    InMux I__7372 (
            .O(N__38118),
            .I(N__38111));
    InMux I__7371 (
            .O(N__38117),
            .I(N__38108));
    Span4Mux_v I__7370 (
            .O(N__38114),
            .I(N__38105));
    LocalMux I__7369 (
            .O(N__38111),
            .I(cmd_rdadctmp_8));
    LocalMux I__7368 (
            .O(N__38108),
            .I(cmd_rdadctmp_8));
    Odrv4 I__7367 (
            .O(N__38105),
            .I(cmd_rdadctmp_8));
    InMux I__7366 (
            .O(N__38098),
            .I(N__38094));
    CascadeMux I__7365 (
            .O(N__38097),
            .I(N__38091));
    LocalMux I__7364 (
            .O(N__38094),
            .I(N__38088));
    InMux I__7363 (
            .O(N__38091),
            .I(N__38084));
    Span12Mux_v I__7362 (
            .O(N__38088),
            .I(N__38081));
    InMux I__7361 (
            .O(N__38087),
            .I(N__38078));
    LocalMux I__7360 (
            .O(N__38084),
            .I(buf_adcdata_iac_0));
    Odrv12 I__7359 (
            .O(N__38081),
            .I(buf_adcdata_iac_0));
    LocalMux I__7358 (
            .O(N__38078),
            .I(buf_adcdata_iac_0));
    InMux I__7357 (
            .O(N__38071),
            .I(N__38068));
    LocalMux I__7356 (
            .O(N__38068),
            .I(N__38065));
    Span4Mux_h I__7355 (
            .O(N__38065),
            .I(N__38062));
    Span4Mux_v I__7354 (
            .O(N__38062),
            .I(N__38058));
    InMux I__7353 (
            .O(N__38061),
            .I(N__38055));
    Odrv4 I__7352 (
            .O(N__38058),
            .I(buf_adcdata_vdc_13));
    LocalMux I__7351 (
            .O(N__38055),
            .I(buf_adcdata_vdc_13));
    InMux I__7350 (
            .O(N__38050),
            .I(N__38047));
    LocalMux I__7349 (
            .O(N__38047),
            .I(N__38044));
    Span4Mux_v I__7348 (
            .O(N__38044),
            .I(N__38040));
    InMux I__7347 (
            .O(N__38043),
            .I(N__38037));
    Span4Mux_h I__7346 (
            .O(N__38040),
            .I(N__38033));
    LocalMux I__7345 (
            .O(N__38037),
            .I(N__38030));
    InMux I__7344 (
            .O(N__38036),
            .I(N__38027));
    Span4Mux_h I__7343 (
            .O(N__38033),
            .I(N__38022));
    Span4Mux_v I__7342 (
            .O(N__38030),
            .I(N__38022));
    LocalMux I__7341 (
            .O(N__38027),
            .I(buf_adcdata_vac_13));
    Odrv4 I__7340 (
            .O(N__38022),
            .I(buf_adcdata_vac_13));
    InMux I__7339 (
            .O(N__38017),
            .I(N__38014));
    LocalMux I__7338 (
            .O(N__38014),
            .I(N__38011));
    Span4Mux_v I__7337 (
            .O(N__38011),
            .I(N__38008));
    Span4Mux_h I__7336 (
            .O(N__38008),
            .I(N__38005));
    Span4Mux_h I__7335 (
            .O(N__38005),
            .I(N__38001));
    InMux I__7334 (
            .O(N__38004),
            .I(N__37998));
    Odrv4 I__7333 (
            .O(N__38001),
            .I(buf_readRTD_5));
    LocalMux I__7332 (
            .O(N__37998),
            .I(buf_readRTD_5));
    CascadeMux I__7331 (
            .O(N__37993),
            .I(n19_adj_1729_cascade_));
    InMux I__7330 (
            .O(N__37990),
            .I(N__37986));
    InMux I__7329 (
            .O(N__37989),
            .I(N__37983));
    LocalMux I__7328 (
            .O(N__37986),
            .I(N__37980));
    LocalMux I__7327 (
            .O(N__37983),
            .I(comm_buf_6_6));
    Odrv4 I__7326 (
            .O(N__37980),
            .I(comm_buf_6_6));
    CascadeMux I__7325 (
            .O(N__37975),
            .I(n9_adj_1600_cascade_));
    CascadeMux I__7324 (
            .O(N__37972),
            .I(n6776_cascade_));
    InMux I__7323 (
            .O(N__37969),
            .I(N__37966));
    LocalMux I__7322 (
            .O(N__37966),
            .I(N__37963));
    Span4Mux_v I__7321 (
            .O(N__37963),
            .I(N__37960));
    Odrv4 I__7320 (
            .O(N__37960),
            .I(n18890));
    InMux I__7319 (
            .O(N__37957),
            .I(N__37954));
    LocalMux I__7318 (
            .O(N__37954),
            .I(N__37951));
    Span4Mux_v I__7317 (
            .O(N__37951),
            .I(N__37948));
    Odrv4 I__7316 (
            .O(N__37948),
            .I(n23390));
    CascadeMux I__7315 (
            .O(N__37945),
            .I(n1_adj_1674_cascade_));
    InMux I__7314 (
            .O(N__37942),
            .I(N__37935));
    InMux I__7313 (
            .O(N__37941),
            .I(N__37935));
    InMux I__7312 (
            .O(N__37940),
            .I(N__37932));
    LocalMux I__7311 (
            .O(N__37935),
            .I(N__37929));
    LocalMux I__7310 (
            .O(N__37932),
            .I(N__37926));
    Odrv12 I__7309 (
            .O(N__37929),
            .I(comm_tx_buf_1));
    Odrv4 I__7308 (
            .O(N__37926),
            .I(comm_tx_buf_1));
    CascadeMux I__7307 (
            .O(N__37921),
            .I(N__37918));
    InMux I__7306 (
            .O(N__37918),
            .I(N__37915));
    LocalMux I__7305 (
            .O(N__37915),
            .I(N__37912));
    Odrv4 I__7304 (
            .O(N__37912),
            .I(n22341));
    InMux I__7303 (
            .O(N__37909),
            .I(N__37906));
    LocalMux I__7302 (
            .O(N__37906),
            .I(n2_adj_1675));
    InMux I__7301 (
            .O(N__37903),
            .I(N__37900));
    LocalMux I__7300 (
            .O(N__37900),
            .I(N__37896));
    CascadeMux I__7299 (
            .O(N__37899),
            .I(N__37893));
    Sp12to4 I__7298 (
            .O(N__37896),
            .I(N__37890));
    InMux I__7297 (
            .O(N__37893),
            .I(N__37887));
    Odrv12 I__7296 (
            .O(N__37890),
            .I(buf_adcdata_vdc_0));
    LocalMux I__7295 (
            .O(N__37887),
            .I(buf_adcdata_vdc_0));
    InMux I__7294 (
            .O(N__37882),
            .I(N__37879));
    LocalMux I__7293 (
            .O(N__37879),
            .I(N__37875));
    InMux I__7292 (
            .O(N__37878),
            .I(N__37871));
    Span12Mux_s10_h I__7291 (
            .O(N__37875),
            .I(N__37868));
    InMux I__7290 (
            .O(N__37874),
            .I(N__37865));
    LocalMux I__7289 (
            .O(N__37871),
            .I(buf_adcdata_vac_0));
    Odrv12 I__7288 (
            .O(N__37868),
            .I(buf_adcdata_vac_0));
    LocalMux I__7287 (
            .O(N__37865),
            .I(buf_adcdata_vac_0));
    CascadeMux I__7286 (
            .O(N__37858),
            .I(n19_adj_1590_cascade_));
    InMux I__7285 (
            .O(N__37855),
            .I(N__37852));
    LocalMux I__7284 (
            .O(N__37852),
            .I(N__37849));
    Span4Mux_v I__7283 (
            .O(N__37849),
            .I(N__37846));
    Odrv4 I__7282 (
            .O(N__37846),
            .I(n22_adj_1589));
    CascadeMux I__7281 (
            .O(N__37843),
            .I(n21965_cascade_));
    InMux I__7280 (
            .O(N__37840),
            .I(N__37833));
    InMux I__7279 (
            .O(N__37839),
            .I(N__37825));
    InMux I__7278 (
            .O(N__37838),
            .I(N__37825));
    InMux I__7277 (
            .O(N__37837),
            .I(N__37816));
    InMux I__7276 (
            .O(N__37836),
            .I(N__37816));
    LocalMux I__7275 (
            .O(N__37833),
            .I(N__37811));
    InMux I__7274 (
            .O(N__37832),
            .I(N__37807));
    InMux I__7273 (
            .O(N__37831),
            .I(N__37802));
    InMux I__7272 (
            .O(N__37830),
            .I(N__37802));
    LocalMux I__7271 (
            .O(N__37825),
            .I(N__37797));
    InMux I__7270 (
            .O(N__37824),
            .I(N__37786));
    InMux I__7269 (
            .O(N__37823),
            .I(N__37779));
    InMux I__7268 (
            .O(N__37822),
            .I(N__37779));
    InMux I__7267 (
            .O(N__37821),
            .I(N__37779));
    LocalMux I__7266 (
            .O(N__37816),
            .I(N__37776));
    InMux I__7265 (
            .O(N__37815),
            .I(N__37773));
    InMux I__7264 (
            .O(N__37814),
            .I(N__37769));
    Span4Mux_v I__7263 (
            .O(N__37811),
            .I(N__37766));
    InMux I__7262 (
            .O(N__37810),
            .I(N__37763));
    LocalMux I__7261 (
            .O(N__37807),
            .I(N__37758));
    LocalMux I__7260 (
            .O(N__37802),
            .I(N__37758));
    InMux I__7259 (
            .O(N__37801),
            .I(N__37755));
    InMux I__7258 (
            .O(N__37800),
            .I(N__37752));
    Span4Mux_v I__7257 (
            .O(N__37797),
            .I(N__37749));
    InMux I__7256 (
            .O(N__37796),
            .I(N__37740));
    InMux I__7255 (
            .O(N__37795),
            .I(N__37737));
    InMux I__7254 (
            .O(N__37794),
            .I(N__37732));
    InMux I__7253 (
            .O(N__37793),
            .I(N__37732));
    InMux I__7252 (
            .O(N__37792),
            .I(N__37723));
    InMux I__7251 (
            .O(N__37791),
            .I(N__37723));
    InMux I__7250 (
            .O(N__37790),
            .I(N__37723));
    InMux I__7249 (
            .O(N__37789),
            .I(N__37723));
    LocalMux I__7248 (
            .O(N__37786),
            .I(N__37718));
    LocalMux I__7247 (
            .O(N__37779),
            .I(N__37718));
    Span4Mux_h I__7246 (
            .O(N__37776),
            .I(N__37713));
    LocalMux I__7245 (
            .O(N__37773),
            .I(N__37713));
    InMux I__7244 (
            .O(N__37772),
            .I(N__37710));
    LocalMux I__7243 (
            .O(N__37769),
            .I(N__37707));
    Span4Mux_h I__7242 (
            .O(N__37766),
            .I(N__37700));
    LocalMux I__7241 (
            .O(N__37763),
            .I(N__37700));
    Span4Mux_v I__7240 (
            .O(N__37758),
            .I(N__37700));
    LocalMux I__7239 (
            .O(N__37755),
            .I(N__37697));
    LocalMux I__7238 (
            .O(N__37752),
            .I(N__37692));
    Sp12to4 I__7237 (
            .O(N__37749),
            .I(N__37692));
    InMux I__7236 (
            .O(N__37748),
            .I(N__37689));
    InMux I__7235 (
            .O(N__37747),
            .I(N__37678));
    InMux I__7234 (
            .O(N__37746),
            .I(N__37678));
    InMux I__7233 (
            .O(N__37745),
            .I(N__37678));
    InMux I__7232 (
            .O(N__37744),
            .I(N__37678));
    InMux I__7231 (
            .O(N__37743),
            .I(N__37678));
    LocalMux I__7230 (
            .O(N__37740),
            .I(N__37671));
    LocalMux I__7229 (
            .O(N__37737),
            .I(N__37671));
    LocalMux I__7228 (
            .O(N__37732),
            .I(N__37671));
    LocalMux I__7227 (
            .O(N__37723),
            .I(N__37668));
    Span4Mux_v I__7226 (
            .O(N__37718),
            .I(N__37665));
    Span4Mux_h I__7225 (
            .O(N__37713),
            .I(N__37662));
    LocalMux I__7224 (
            .O(N__37710),
            .I(N__37655));
    Span4Mux_h I__7223 (
            .O(N__37707),
            .I(N__37655));
    Span4Mux_h I__7222 (
            .O(N__37700),
            .I(N__37655));
    Sp12to4 I__7221 (
            .O(N__37697),
            .I(N__37650));
    Span12Mux_h I__7220 (
            .O(N__37692),
            .I(N__37650));
    LocalMux I__7219 (
            .O(N__37689),
            .I(n13746));
    LocalMux I__7218 (
            .O(N__37678),
            .I(n13746));
    Odrv12 I__7217 (
            .O(N__37671),
            .I(n13746));
    Odrv4 I__7216 (
            .O(N__37668),
            .I(n13746));
    Odrv4 I__7215 (
            .O(N__37665),
            .I(n13746));
    Odrv4 I__7214 (
            .O(N__37662),
            .I(n13746));
    Odrv4 I__7213 (
            .O(N__37655),
            .I(n13746));
    Odrv12 I__7212 (
            .O(N__37650),
            .I(n13746));
    InMux I__7211 (
            .O(N__37633),
            .I(N__37630));
    LocalMux I__7210 (
            .O(N__37630),
            .I(N__37627));
    Span4Mux_v I__7209 (
            .O(N__37627),
            .I(N__37623));
    InMux I__7208 (
            .O(N__37626),
            .I(N__37620));
    Sp12to4 I__7207 (
            .O(N__37623),
            .I(N__37615));
    LocalMux I__7206 (
            .O(N__37620),
            .I(N__37615));
    Odrv12 I__7205 (
            .O(N__37615),
            .I(\comm_spi.n15323 ));
    SRMux I__7204 (
            .O(N__37612),
            .I(N__37609));
    LocalMux I__7203 (
            .O(N__37609),
            .I(N__37606));
    Odrv4 I__7202 (
            .O(N__37606),
            .I(\comm_spi.data_tx_7__N_860 ));
    InMux I__7201 (
            .O(N__37603),
            .I(N__37600));
    LocalMux I__7200 (
            .O(N__37600),
            .I(N__37595));
    InMux I__7199 (
            .O(N__37599),
            .I(N__37592));
    InMux I__7198 (
            .O(N__37598),
            .I(N__37589));
    Odrv4 I__7197 (
            .O(N__37595),
            .I(\comm_spi.n24040 ));
    LocalMux I__7196 (
            .O(N__37592),
            .I(\comm_spi.n24040 ));
    LocalMux I__7195 (
            .O(N__37589),
            .I(\comm_spi.n24040 ));
    SRMux I__7194 (
            .O(N__37582),
            .I(N__37579));
    LocalMux I__7193 (
            .O(N__37579),
            .I(N__37576));
    Odrv12 I__7192 (
            .O(N__37576),
            .I(\comm_spi.data_tx_7__N_880 ));
    CascadeMux I__7191 (
            .O(N__37573),
            .I(N__37570));
    InMux I__7190 (
            .O(N__37570),
            .I(N__37567));
    LocalMux I__7189 (
            .O(N__37567),
            .I(N__37564));
    Span4Mux_v I__7188 (
            .O(N__37564),
            .I(N__37560));
    InMux I__7187 (
            .O(N__37563),
            .I(N__37557));
    Span4Mux_v I__7186 (
            .O(N__37560),
            .I(N__37553));
    LocalMux I__7185 (
            .O(N__37557),
            .I(N__37550));
    InMux I__7184 (
            .O(N__37556),
            .I(N__37547));
    Odrv4 I__7183 (
            .O(N__37553),
            .I(\comm_spi.n24037 ));
    Odrv4 I__7182 (
            .O(N__37550),
            .I(\comm_spi.n24037 ));
    LocalMux I__7181 (
            .O(N__37547),
            .I(\comm_spi.n24037 ));
    InMux I__7180 (
            .O(N__37540),
            .I(N__37537));
    LocalMux I__7179 (
            .O(N__37537),
            .I(N__37534));
    Span4Mux_v I__7178 (
            .O(N__37534),
            .I(N__37530));
    InMux I__7177 (
            .O(N__37533),
            .I(N__37527));
    Span4Mux_v I__7176 (
            .O(N__37530),
            .I(N__37522));
    LocalMux I__7175 (
            .O(N__37527),
            .I(N__37522));
    Odrv4 I__7174 (
            .O(N__37522),
            .I(\comm_spi.n15348 ));
    InMux I__7173 (
            .O(N__37519),
            .I(N__37516));
    LocalMux I__7172 (
            .O(N__37516),
            .I(N__37513));
    Span4Mux_v I__7171 (
            .O(N__37513),
            .I(N__37510));
    Span4Mux_v I__7170 (
            .O(N__37510),
            .I(N__37506));
    InMux I__7169 (
            .O(N__37509),
            .I(N__37503));
    Span4Mux_v I__7168 (
            .O(N__37506),
            .I(N__37500));
    LocalMux I__7167 (
            .O(N__37503),
            .I(N__37497));
    Odrv4 I__7166 (
            .O(N__37500),
            .I(\comm_spi.n15349 ));
    Odrv12 I__7165 (
            .O(N__37497),
            .I(\comm_spi.n15349 ));
    InMux I__7164 (
            .O(N__37492),
            .I(N__37489));
    LocalMux I__7163 (
            .O(N__37489),
            .I(\comm_spi.n15335 ));
    InMux I__7162 (
            .O(N__37486),
            .I(N__37480));
    InMux I__7161 (
            .O(N__37485),
            .I(N__37480));
    LocalMux I__7160 (
            .O(N__37480),
            .I(buf_control_6));
    InMux I__7159 (
            .O(N__37477),
            .I(N__37472));
    InMux I__7158 (
            .O(N__37476),
            .I(N__37467));
    InMux I__7157 (
            .O(N__37475),
            .I(N__37467));
    LocalMux I__7156 (
            .O(N__37472),
            .I(acadc_skipCount_14));
    LocalMux I__7155 (
            .O(N__37467),
            .I(acadc_skipCount_14));
    CascadeMux I__7154 (
            .O(N__37462),
            .I(N__37459));
    InMux I__7153 (
            .O(N__37459),
            .I(N__37456));
    LocalMux I__7152 (
            .O(N__37456),
            .I(N__37453));
    Span12Mux_h I__7151 (
            .O(N__37453),
            .I(N__37450));
    Odrv12 I__7150 (
            .O(N__37450),
            .I(n23_adj_1767));
    CascadeMux I__7149 (
            .O(N__37447),
            .I(N__37444));
    InMux I__7148 (
            .O(N__37444),
            .I(N__37441));
    LocalMux I__7147 (
            .O(N__37441),
            .I(\SIG_DDS.tmp_buf_0 ));
    CascadeMux I__7146 (
            .O(N__37438),
            .I(N__37435));
    InMux I__7145 (
            .O(N__37435),
            .I(N__37432));
    LocalMux I__7144 (
            .O(N__37432),
            .I(N__37429));
    Span4Mux_h I__7143 (
            .O(N__37429),
            .I(N__37426));
    Odrv4 I__7142 (
            .O(N__37426),
            .I(\SIG_DDS.tmp_buf_3 ));
    CascadeMux I__7141 (
            .O(N__37423),
            .I(N__37420));
    InMux I__7140 (
            .O(N__37420),
            .I(N__37417));
    LocalMux I__7139 (
            .O(N__37417),
            .I(\SIG_DDS.tmp_buf_1 ));
    CascadeMux I__7138 (
            .O(N__37414),
            .I(N__37411));
    InMux I__7137 (
            .O(N__37411),
            .I(N__37408));
    LocalMux I__7136 (
            .O(N__37408),
            .I(\SIG_DDS.tmp_buf_2 ));
    InMux I__7135 (
            .O(N__37405),
            .I(N__37398));
    InMux I__7134 (
            .O(N__37404),
            .I(N__37398));
    InMux I__7133 (
            .O(N__37403),
            .I(N__37395));
    LocalMux I__7132 (
            .O(N__37398),
            .I(N__37389));
    LocalMux I__7131 (
            .O(N__37395),
            .I(N__37386));
    InMux I__7130 (
            .O(N__37394),
            .I(N__37383));
    InMux I__7129 (
            .O(N__37393),
            .I(N__37376));
    InMux I__7128 (
            .O(N__37392),
            .I(N__37376));
    Span4Mux_h I__7127 (
            .O(N__37389),
            .I(N__37373));
    Span4Mux_v I__7126 (
            .O(N__37386),
            .I(N__37368));
    LocalMux I__7125 (
            .O(N__37383),
            .I(N__37368));
    InMux I__7124 (
            .O(N__37382),
            .I(N__37365));
    InMux I__7123 (
            .O(N__37381),
            .I(N__37362));
    LocalMux I__7122 (
            .O(N__37376),
            .I(n11979));
    Odrv4 I__7121 (
            .O(N__37373),
            .I(n11979));
    Odrv4 I__7120 (
            .O(N__37368),
            .I(n11979));
    LocalMux I__7119 (
            .O(N__37365),
            .I(n11979));
    LocalMux I__7118 (
            .O(N__37362),
            .I(n11979));
    InMux I__7117 (
            .O(N__37351),
            .I(N__37348));
    LocalMux I__7116 (
            .O(N__37348),
            .I(N__37344));
    InMux I__7115 (
            .O(N__37347),
            .I(N__37341));
    Span4Mux_h I__7114 (
            .O(N__37344),
            .I(N__37338));
    LocalMux I__7113 (
            .O(N__37341),
            .I(acadc_skipcnt_15));
    Odrv4 I__7112 (
            .O(N__37338),
            .I(acadc_skipcnt_15));
    InMux I__7111 (
            .O(N__37333),
            .I(N__37330));
    LocalMux I__7110 (
            .O(N__37330),
            .I(N__37326));
    InMux I__7109 (
            .O(N__37329),
            .I(N__37323));
    Span4Mux_h I__7108 (
            .O(N__37326),
            .I(N__37320));
    LocalMux I__7107 (
            .O(N__37323),
            .I(acadc_skipcnt_9));
    Odrv4 I__7106 (
            .O(N__37320),
            .I(acadc_skipcnt_9));
    InMux I__7105 (
            .O(N__37315),
            .I(N__37311));
    InMux I__7104 (
            .O(N__37314),
            .I(N__37308));
    LocalMux I__7103 (
            .O(N__37311),
            .I(N__37305));
    LocalMux I__7102 (
            .O(N__37308),
            .I(acadc_skipcnt_14));
    Odrv4 I__7101 (
            .O(N__37305),
            .I(acadc_skipcnt_14));
    InMux I__7100 (
            .O(N__37300),
            .I(N__37296));
    InMux I__7099 (
            .O(N__37299),
            .I(N__37293));
    LocalMux I__7098 (
            .O(N__37296),
            .I(N__37290));
    LocalMux I__7097 (
            .O(N__37293),
            .I(acadc_skipcnt_11));
    Odrv4 I__7096 (
            .O(N__37290),
            .I(acadc_skipcnt_11));
    CascadeMux I__7095 (
            .O(N__37285),
            .I(N__37281));
    InMux I__7094 (
            .O(N__37284),
            .I(N__37276));
    InMux I__7093 (
            .O(N__37281),
            .I(N__37276));
    LocalMux I__7092 (
            .O(N__37276),
            .I(N__37273));
    Span4Mux_h I__7091 (
            .O(N__37273),
            .I(N__37270));
    Span4Mux_h I__7090 (
            .O(N__37270),
            .I(N__37266));
    InMux I__7089 (
            .O(N__37269),
            .I(N__37263));
    Odrv4 I__7088 (
            .O(N__37266),
            .I(cmd_rdadctmp_19));
    LocalMux I__7087 (
            .O(N__37263),
            .I(cmd_rdadctmp_19));
    CascadeMux I__7086 (
            .O(N__37258),
            .I(N__37255));
    InMux I__7085 (
            .O(N__37255),
            .I(N__37251));
    CascadeMux I__7084 (
            .O(N__37254),
            .I(N__37248));
    LocalMux I__7083 (
            .O(N__37251),
            .I(N__37245));
    InMux I__7082 (
            .O(N__37248),
            .I(N__37241));
    Span4Mux_h I__7081 (
            .O(N__37245),
            .I(N__37238));
    InMux I__7080 (
            .O(N__37244),
            .I(N__37235));
    LocalMux I__7079 (
            .O(N__37241),
            .I(cmd_rdadctmp_20));
    Odrv4 I__7078 (
            .O(N__37238),
            .I(cmd_rdadctmp_20));
    LocalMux I__7077 (
            .O(N__37235),
            .I(cmd_rdadctmp_20));
    CascadeMux I__7076 (
            .O(N__37228),
            .I(N__37224));
    InMux I__7075 (
            .O(N__37227),
            .I(N__37221));
    InMux I__7074 (
            .O(N__37224),
            .I(N__37217));
    LocalMux I__7073 (
            .O(N__37221),
            .I(N__37214));
    InMux I__7072 (
            .O(N__37220),
            .I(N__37211));
    LocalMux I__7071 (
            .O(N__37217),
            .I(N__37208));
    Span4Mux_h I__7070 (
            .O(N__37214),
            .I(N__37205));
    LocalMux I__7069 (
            .O(N__37211),
            .I(buf_dds1_0));
    Odrv4 I__7068 (
            .O(N__37208),
            .I(buf_dds1_0));
    Odrv4 I__7067 (
            .O(N__37205),
            .I(buf_dds1_0));
    CascadeMux I__7066 (
            .O(N__37198),
            .I(N__37195));
    InMux I__7065 (
            .O(N__37195),
            .I(N__37192));
    LocalMux I__7064 (
            .O(N__37192),
            .I(N__37189));
    Span4Mux_h I__7063 (
            .O(N__37189),
            .I(N__37184));
    InMux I__7062 (
            .O(N__37188),
            .I(N__37181));
    InMux I__7061 (
            .O(N__37187),
            .I(N__37178));
    Odrv4 I__7060 (
            .O(N__37184),
            .I(cmd_rdadctmp_28));
    LocalMux I__7059 (
            .O(N__37181),
            .I(cmd_rdadctmp_28));
    LocalMux I__7058 (
            .O(N__37178),
            .I(cmd_rdadctmp_28));
    InMux I__7057 (
            .O(N__37171),
            .I(N__37168));
    LocalMux I__7056 (
            .O(N__37168),
            .I(N__37165));
    Span12Mux_s10_v I__7055 (
            .O(N__37165),
            .I(N__37160));
    InMux I__7054 (
            .O(N__37164),
            .I(N__37157));
    InMux I__7053 (
            .O(N__37163),
            .I(N__37154));
    Span12Mux_v I__7052 (
            .O(N__37160),
            .I(N__37151));
    LocalMux I__7051 (
            .O(N__37157),
            .I(N__37148));
    LocalMux I__7050 (
            .O(N__37154),
            .I(buf_adcdata_iac_20));
    Odrv12 I__7049 (
            .O(N__37151),
            .I(buf_adcdata_iac_20));
    Odrv4 I__7048 (
            .O(N__37148),
            .I(buf_adcdata_iac_20));
    SRMux I__7047 (
            .O(N__37141),
            .I(N__37138));
    LocalMux I__7046 (
            .O(N__37138),
            .I(N__37135));
    Span4Mux_h I__7045 (
            .O(N__37135),
            .I(N__37131));
    SRMux I__7044 (
            .O(N__37134),
            .I(N__37127));
    Span4Mux_v I__7043 (
            .O(N__37131),
            .I(N__37123));
    SRMux I__7042 (
            .O(N__37130),
            .I(N__37120));
    LocalMux I__7041 (
            .O(N__37127),
            .I(N__37117));
    SRMux I__7040 (
            .O(N__37126),
            .I(N__37114));
    Span4Mux_v I__7039 (
            .O(N__37123),
            .I(N__37109));
    LocalMux I__7038 (
            .O(N__37120),
            .I(N__37109));
    Span4Mux_v I__7037 (
            .O(N__37117),
            .I(N__37104));
    LocalMux I__7036 (
            .O(N__37114),
            .I(N__37104));
    Span4Mux_v I__7035 (
            .O(N__37109),
            .I(N__37101));
    Span4Mux_v I__7034 (
            .O(N__37104),
            .I(N__37098));
    Span4Mux_v I__7033 (
            .O(N__37101),
            .I(N__37095));
    Span4Mux_h I__7032 (
            .O(N__37098),
            .I(N__37092));
    Odrv4 I__7031 (
            .O(N__37095),
            .I(n15538));
    Odrv4 I__7030 (
            .O(N__37092),
            .I(n15538));
    IoInMux I__7029 (
            .O(N__37087),
            .I(N__37084));
    LocalMux I__7028 (
            .O(N__37084),
            .I(N__37080));
    CascadeMux I__7027 (
            .O(N__37083),
            .I(N__37076));
    Span12Mux_s11_v I__7026 (
            .O(N__37080),
            .I(N__37073));
    InMux I__7025 (
            .O(N__37079),
            .I(N__37070));
    InMux I__7024 (
            .O(N__37076),
            .I(N__37067));
    Odrv12 I__7023 (
            .O(N__37073),
            .I(IAC_OSR0));
    LocalMux I__7022 (
            .O(N__37070),
            .I(IAC_OSR0));
    LocalMux I__7021 (
            .O(N__37067),
            .I(IAC_OSR0));
    InMux I__7020 (
            .O(N__37060),
            .I(N__37057));
    LocalMux I__7019 (
            .O(N__37057),
            .I(n24_adj_1575));
    IoInMux I__7018 (
            .O(N__37054),
            .I(N__37051));
    LocalMux I__7017 (
            .O(N__37051),
            .I(N__37048));
    Span4Mux_s2_v I__7016 (
            .O(N__37048),
            .I(N__37044));
    InMux I__7015 (
            .O(N__37047),
            .I(N__37041));
    Span4Mux_h I__7014 (
            .O(N__37044),
            .I(N__37038));
    LocalMux I__7013 (
            .O(N__37041),
            .I(N__37034));
    Sp12to4 I__7012 (
            .O(N__37038),
            .I(N__37031));
    InMux I__7011 (
            .O(N__37037),
            .I(N__37028));
    Span4Mux_h I__7010 (
            .O(N__37034),
            .I(N__37025));
    Odrv12 I__7009 (
            .O(N__37031),
            .I(IAC_OSR1));
    LocalMux I__7008 (
            .O(N__37028),
            .I(IAC_OSR1));
    Odrv4 I__7007 (
            .O(N__37025),
            .I(IAC_OSR1));
    InMux I__7006 (
            .O(N__37018),
            .I(N__37015));
    LocalMux I__7005 (
            .O(N__37015),
            .I(n24_adj_1601));
    InMux I__7004 (
            .O(N__37012),
            .I(N__37009));
    LocalMux I__7003 (
            .O(N__37009),
            .I(n11984));
    InMux I__7002 (
            .O(N__37006),
            .I(N__37003));
    LocalMux I__7001 (
            .O(N__37003),
            .I(N__37000));
    Odrv4 I__7000 (
            .O(N__37000),
            .I(n16_adj_1733));
    InMux I__6999 (
            .O(N__36997),
            .I(N__36994));
    LocalMux I__6998 (
            .O(N__36994),
            .I(N__36991));
    Span12Mux_v I__6997 (
            .O(N__36991),
            .I(N__36988));
    Odrv12 I__6996 (
            .O(N__36988),
            .I(n23438));
    InMux I__6995 (
            .O(N__36985),
            .I(N__36982));
    LocalMux I__6994 (
            .O(N__36982),
            .I(N__36979));
    Span4Mux_v I__6993 (
            .O(N__36979),
            .I(N__36974));
    CascadeMux I__6992 (
            .O(N__36978),
            .I(N__36971));
    InMux I__6991 (
            .O(N__36977),
            .I(N__36968));
    Sp12to4 I__6990 (
            .O(N__36974),
            .I(N__36965));
    InMux I__6989 (
            .O(N__36971),
            .I(N__36962));
    LocalMux I__6988 (
            .O(N__36968),
            .I(buf_adcdata_iac_12));
    Odrv12 I__6987 (
            .O(N__36965),
            .I(buf_adcdata_iac_12));
    LocalMux I__6986 (
            .O(N__36962),
            .I(buf_adcdata_iac_12));
    CascadeMux I__6985 (
            .O(N__36955),
            .I(N__36952));
    InMux I__6984 (
            .O(N__36952),
            .I(N__36948));
    InMux I__6983 (
            .O(N__36951),
            .I(N__36945));
    LocalMux I__6982 (
            .O(N__36948),
            .I(comm_test_buf_24_21));
    LocalMux I__6981 (
            .O(N__36945),
            .I(comm_test_buf_24_21));
    InMux I__6980 (
            .O(N__36940),
            .I(N__36937));
    LocalMux I__6979 (
            .O(N__36937),
            .I(N__36934));
    Span4Mux_h I__6978 (
            .O(N__36934),
            .I(N__36930));
    InMux I__6977 (
            .O(N__36933),
            .I(N__36927));
    Span4Mux_v I__6976 (
            .O(N__36930),
            .I(N__36922));
    LocalMux I__6975 (
            .O(N__36927),
            .I(N__36922));
    Odrv4 I__6974 (
            .O(N__36922),
            .I(comm_test_buf_24_13));
    InMux I__6973 (
            .O(N__36919),
            .I(N__36915));
    InMux I__6972 (
            .O(N__36918),
            .I(N__36911));
    LocalMux I__6971 (
            .O(N__36915),
            .I(N__36908));
    InMux I__6970 (
            .O(N__36914),
            .I(N__36905));
    LocalMux I__6969 (
            .O(N__36911),
            .I(N__36902));
    Span4Mux_h I__6968 (
            .O(N__36908),
            .I(N__36899));
    LocalMux I__6967 (
            .O(N__36905),
            .I(N__36896));
    Span4Mux_h I__6966 (
            .O(N__36902),
            .I(N__36891));
    Span4Mux_h I__6965 (
            .O(N__36899),
            .I(N__36891));
    Span4Mux_v I__6964 (
            .O(N__36896),
            .I(N__36888));
    Odrv4 I__6963 (
            .O(N__36891),
            .I(comm_test_buf_24_5));
    Odrv4 I__6962 (
            .O(N__36888),
            .I(comm_test_buf_24_5));
    CascadeMux I__6961 (
            .O(N__36883),
            .I(n111_adj_1776_cascade_));
    InMux I__6960 (
            .O(N__36880),
            .I(N__36877));
    LocalMux I__6959 (
            .O(N__36877),
            .I(N__36874));
    Span4Mux_h I__6958 (
            .O(N__36874),
            .I(N__36871));
    Odrv4 I__6957 (
            .O(N__36871),
            .I(n111_adj_1761));
    InMux I__6956 (
            .O(N__36868),
            .I(N__36864));
    InMux I__6955 (
            .O(N__36867),
            .I(N__36861));
    LocalMux I__6954 (
            .O(N__36864),
            .I(N__36857));
    LocalMux I__6953 (
            .O(N__36861),
            .I(N__36854));
    InMux I__6952 (
            .O(N__36860),
            .I(N__36851));
    Span4Mux_h I__6951 (
            .O(N__36857),
            .I(N__36846));
    Span4Mux_h I__6950 (
            .O(N__36854),
            .I(N__36846));
    LocalMux I__6949 (
            .O(N__36851),
            .I(buf_dds1_3));
    Odrv4 I__6948 (
            .O(N__36846),
            .I(buf_dds1_3));
    InMux I__6947 (
            .O(N__36841),
            .I(N__36838));
    LocalMux I__6946 (
            .O(N__36838),
            .I(N__36835));
    Span4Mux_v I__6945 (
            .O(N__36835),
            .I(N__36830));
    InMux I__6944 (
            .O(N__36834),
            .I(N__36825));
    InMux I__6943 (
            .O(N__36833),
            .I(N__36825));
    Span4Mux_h I__6942 (
            .O(N__36830),
            .I(N__36820));
    LocalMux I__6941 (
            .O(N__36825),
            .I(N__36820));
    Odrv4 I__6940 (
            .O(N__36820),
            .I(comm_buf_2_4));
    CascadeMux I__6939 (
            .O(N__36817),
            .I(n11987_cascade_));
    InMux I__6938 (
            .O(N__36814),
            .I(N__36811));
    LocalMux I__6937 (
            .O(N__36811),
            .I(N__36808));
    Span4Mux_v I__6936 (
            .O(N__36808),
            .I(N__36805));
    Odrv4 I__6935 (
            .O(N__36805),
            .I(n17_adj_1779));
    CascadeMux I__6934 (
            .O(N__36802),
            .I(n11985_cascade_));
    CEMux I__6933 (
            .O(N__36799),
            .I(N__36795));
    CEMux I__6932 (
            .O(N__36798),
            .I(N__36791));
    LocalMux I__6931 (
            .O(N__36795),
            .I(N__36787));
    CEMux I__6930 (
            .O(N__36794),
            .I(N__36784));
    LocalMux I__6929 (
            .O(N__36791),
            .I(N__36781));
    CEMux I__6928 (
            .O(N__36790),
            .I(N__36778));
    Span4Mux_v I__6927 (
            .O(N__36787),
            .I(N__36774));
    LocalMux I__6926 (
            .O(N__36784),
            .I(N__36769));
    Span4Mux_h I__6925 (
            .O(N__36781),
            .I(N__36769));
    LocalMux I__6924 (
            .O(N__36778),
            .I(N__36766));
    InMux I__6923 (
            .O(N__36777),
            .I(N__36763));
    Span4Mux_v I__6922 (
            .O(N__36774),
            .I(N__36760));
    Span4Mux_v I__6921 (
            .O(N__36769),
            .I(N__36757));
    Span4Mux_v I__6920 (
            .O(N__36766),
            .I(N__36752));
    LocalMux I__6919 (
            .O(N__36763),
            .I(N__36752));
    Span4Mux_v I__6918 (
            .O(N__36760),
            .I(N__36749));
    Sp12to4 I__6917 (
            .O(N__36757),
            .I(N__36746));
    Span4Mux_v I__6916 (
            .O(N__36752),
            .I(N__36743));
    Span4Mux_h I__6915 (
            .O(N__36749),
            .I(N__36740));
    Span12Mux_v I__6914 (
            .O(N__36746),
            .I(N__36737));
    Span4Mux_h I__6913 (
            .O(N__36743),
            .I(N__36734));
    Odrv4 I__6912 (
            .O(N__36740),
            .I(n13117));
    Odrv12 I__6911 (
            .O(N__36737),
            .I(n13117));
    Odrv4 I__6910 (
            .O(N__36734),
            .I(n13117));
    InMux I__6909 (
            .O(N__36727),
            .I(N__36724));
    LocalMux I__6908 (
            .O(N__36724),
            .I(N__36721));
    Span4Mux_h I__6907 (
            .O(N__36721),
            .I(N__36718));
    Odrv4 I__6906 (
            .O(N__36718),
            .I(comm_buf_2_7_N_575_7));
    SRMux I__6905 (
            .O(N__36715),
            .I(N__36712));
    LocalMux I__6904 (
            .O(N__36712),
            .I(N__36709));
    Span4Mux_h I__6903 (
            .O(N__36709),
            .I(N__36706));
    Span4Mux_v I__6902 (
            .O(N__36706),
            .I(N__36703));
    Odrv4 I__6901 (
            .O(N__36703),
            .I(\comm_spi.data_tx_7__N_859 ));
    InMux I__6900 (
            .O(N__36700),
            .I(N__36675));
    InMux I__6899 (
            .O(N__36699),
            .I(N__36675));
    InMux I__6898 (
            .O(N__36698),
            .I(N__36675));
    InMux I__6897 (
            .O(N__36697),
            .I(N__36675));
    InMux I__6896 (
            .O(N__36696),
            .I(N__36675));
    InMux I__6895 (
            .O(N__36695),
            .I(N__36675));
    InMux I__6894 (
            .O(N__36694),
            .I(N__36675));
    InMux I__6893 (
            .O(N__36693),
            .I(N__36675));
    InMux I__6892 (
            .O(N__36692),
            .I(N__36672));
    LocalMux I__6891 (
            .O(N__36675),
            .I(N__36662));
    LocalMux I__6890 (
            .O(N__36672),
            .I(N__36659));
    InMux I__6889 (
            .O(N__36671),
            .I(N__36644));
    InMux I__6888 (
            .O(N__36670),
            .I(N__36644));
    InMux I__6887 (
            .O(N__36669),
            .I(N__36644));
    InMux I__6886 (
            .O(N__36668),
            .I(N__36644));
    InMux I__6885 (
            .O(N__36667),
            .I(N__36644));
    InMux I__6884 (
            .O(N__36666),
            .I(N__36644));
    InMux I__6883 (
            .O(N__36665),
            .I(N__36644));
    Sp12to4 I__6882 (
            .O(N__36662),
            .I(N__36641));
    Odrv4 I__6881 (
            .O(N__36659),
            .I(n6774));
    LocalMux I__6880 (
            .O(N__36644),
            .I(n6774));
    Odrv12 I__6879 (
            .O(N__36641),
            .I(n6774));
    CascadeMux I__6878 (
            .O(N__36634),
            .I(n111_adj_1796_cascade_));
    InMux I__6877 (
            .O(N__36631),
            .I(N__36625));
    InMux I__6876 (
            .O(N__36630),
            .I(N__36625));
    LocalMux I__6875 (
            .O(N__36625),
            .I(comm_test_buf_24_10));
    InMux I__6874 (
            .O(N__36622),
            .I(N__36619));
    LocalMux I__6873 (
            .O(N__36619),
            .I(N__36616));
    Span4Mux_v I__6872 (
            .O(N__36616),
            .I(N__36612));
    InMux I__6871 (
            .O(N__36615),
            .I(N__36609));
    Span4Mux_h I__6870 (
            .O(N__36612),
            .I(N__36606));
    LocalMux I__6869 (
            .O(N__36609),
            .I(N__36603));
    Odrv4 I__6868 (
            .O(N__36606),
            .I(\comm_spi.n15365 ));
    Odrv4 I__6867 (
            .O(N__36603),
            .I(\comm_spi.n15365 ));
    InMux I__6866 (
            .O(N__36598),
            .I(N__36595));
    LocalMux I__6865 (
            .O(N__36595),
            .I(N__36592));
    Span4Mux_v I__6864 (
            .O(N__36592),
            .I(N__36587));
    InMux I__6863 (
            .O(N__36591),
            .I(N__36584));
    InMux I__6862 (
            .O(N__36590),
            .I(N__36581));
    Odrv4 I__6861 (
            .O(N__36587),
            .I(\comm_spi.n24025 ));
    LocalMux I__6860 (
            .O(N__36584),
            .I(\comm_spi.n24025 ));
    LocalMux I__6859 (
            .O(N__36581),
            .I(\comm_spi.n24025 ));
    InMux I__6858 (
            .O(N__36574),
            .I(N__36571));
    LocalMux I__6857 (
            .O(N__36571),
            .I(N__36568));
    Span4Mux_v I__6856 (
            .O(N__36568),
            .I(N__36565));
    Span4Mux_v I__6855 (
            .O(N__36565),
            .I(N__36561));
    InMux I__6854 (
            .O(N__36564),
            .I(N__36558));
    Odrv4 I__6853 (
            .O(N__36561),
            .I(\comm_spi.n15364 ));
    LocalMux I__6852 (
            .O(N__36558),
            .I(\comm_spi.n15364 ));
    InMux I__6851 (
            .O(N__36553),
            .I(N__36549));
    InMux I__6850 (
            .O(N__36552),
            .I(N__36546));
    LocalMux I__6849 (
            .O(N__36549),
            .I(N__36543));
    LocalMux I__6848 (
            .O(N__36546),
            .I(N__36540));
    Span4Mux_v I__6847 (
            .O(N__36543),
            .I(N__36535));
    Span4Mux_v I__6846 (
            .O(N__36540),
            .I(N__36535));
    Span4Mux_v I__6845 (
            .O(N__36535),
            .I(N__36532));
    Odrv4 I__6844 (
            .O(N__36532),
            .I(\comm_spi.n15368 ));
    SRMux I__6843 (
            .O(N__36529),
            .I(N__36526));
    LocalMux I__6842 (
            .O(N__36526),
            .I(N__36523));
    Span4Mux_v I__6841 (
            .O(N__36523),
            .I(N__36520));
    Span4Mux_v I__6840 (
            .O(N__36520),
            .I(N__36517));
    Odrv4 I__6839 (
            .O(N__36517),
            .I(\comm_spi.data_tx_7__N_855 ));
    IoInMux I__6838 (
            .O(N__36514),
            .I(N__36511));
    LocalMux I__6837 (
            .O(N__36511),
            .I(N__36508));
    Span4Mux_s2_h I__6836 (
            .O(N__36508),
            .I(N__36505));
    Span4Mux_v I__6835 (
            .O(N__36505),
            .I(N__36502));
    Sp12to4 I__6834 (
            .O(N__36502),
            .I(N__36497));
    InMux I__6833 (
            .O(N__36501),
            .I(N__36494));
    InMux I__6832 (
            .O(N__36500),
            .I(N__36491));
    Span12Mux_h I__6831 (
            .O(N__36497),
            .I(N__36486));
    LocalMux I__6830 (
            .O(N__36494),
            .I(N__36486));
    LocalMux I__6829 (
            .O(N__36491),
            .I(AMPV_POW));
    Odrv12 I__6828 (
            .O(N__36486),
            .I(AMPV_POW));
    CascadeMux I__6827 (
            .O(N__36481),
            .I(N__36478));
    InMux I__6826 (
            .O(N__36478),
            .I(N__36475));
    LocalMux I__6825 (
            .O(N__36475),
            .I(N__36472));
    Span4Mux_h I__6824 (
            .O(N__36472),
            .I(N__36469));
    Odrv4 I__6823 (
            .O(N__36469),
            .I(comm_buf_0_7_N_543_7));
    InMux I__6822 (
            .O(N__36466),
            .I(N__36462));
    InMux I__6821 (
            .O(N__36465),
            .I(N__36459));
    LocalMux I__6820 (
            .O(N__36462),
            .I(N__36455));
    LocalMux I__6819 (
            .O(N__36459),
            .I(N__36452));
    InMux I__6818 (
            .O(N__36458),
            .I(N__36449));
    Span4Mux_v I__6817 (
            .O(N__36455),
            .I(N__36446));
    Odrv4 I__6816 (
            .O(N__36452),
            .I(clk_cnt_1));
    LocalMux I__6815 (
            .O(N__36449),
            .I(clk_cnt_1));
    Odrv4 I__6814 (
            .O(N__36446),
            .I(clk_cnt_1));
    InMux I__6813 (
            .O(N__36439),
            .I(N__36433));
    InMux I__6812 (
            .O(N__36438),
            .I(N__36430));
    InMux I__6811 (
            .O(N__36437),
            .I(N__36425));
    InMux I__6810 (
            .O(N__36436),
            .I(N__36425));
    LocalMux I__6809 (
            .O(N__36433),
            .I(N__36420));
    LocalMux I__6808 (
            .O(N__36430),
            .I(N__36420));
    LocalMux I__6807 (
            .O(N__36425),
            .I(clk_cnt_0));
    Odrv12 I__6806 (
            .O(N__36420),
            .I(clk_cnt_0));
    SRMux I__6805 (
            .O(N__36415),
            .I(N__36412));
    LocalMux I__6804 (
            .O(N__36412),
            .I(N__36409));
    Span4Mux_v I__6803 (
            .O(N__36409),
            .I(N__36406));
    Span4Mux_h I__6802 (
            .O(N__36406),
            .I(N__36403));
    Odrv4 I__6801 (
            .O(N__36403),
            .I(n18996));
    InMux I__6800 (
            .O(N__36400),
            .I(N__36397));
    LocalMux I__6799 (
            .O(N__36397),
            .I(comm_buf_2_7_N_575_0));
    CascadeMux I__6798 (
            .O(N__36394),
            .I(N__36391));
    InMux I__6797 (
            .O(N__36391),
            .I(N__36388));
    LocalMux I__6796 (
            .O(N__36388),
            .I(N__36385));
    Odrv4 I__6795 (
            .O(N__36385),
            .I(comm_buf_2_7_N_575_1));
    InMux I__6794 (
            .O(N__36382),
            .I(N__36379));
    LocalMux I__6793 (
            .O(N__36379),
            .I(N__36376));
    Odrv4 I__6792 (
            .O(N__36376),
            .I(comm_buf_2_7_N_575_3));
    InMux I__6791 (
            .O(N__36373),
            .I(N__36370));
    LocalMux I__6790 (
            .O(N__36370),
            .I(N__36367));
    Odrv12 I__6789 (
            .O(N__36367),
            .I(comm_buf_2_7_N_575_4));
    InMux I__6788 (
            .O(N__36364),
            .I(N__36361));
    LocalMux I__6787 (
            .O(N__36361),
            .I(N__36358));
    Odrv12 I__6786 (
            .O(N__36358),
            .I(comm_buf_2_7_N_575_5));
    InMux I__6785 (
            .O(N__36355),
            .I(N__36352));
    LocalMux I__6784 (
            .O(N__36352),
            .I(N__36349));
    Odrv12 I__6783 (
            .O(N__36349),
            .I(comm_buf_2_7_N_575_6));
    CascadeMux I__6782 (
            .O(N__36346),
            .I(N__36343));
    InMux I__6781 (
            .O(N__36343),
            .I(N__36338));
    InMux I__6780 (
            .O(N__36342),
            .I(N__36333));
    InMux I__6779 (
            .O(N__36341),
            .I(N__36333));
    LocalMux I__6778 (
            .O(N__36338),
            .I(N__36330));
    LocalMux I__6777 (
            .O(N__36333),
            .I(N__36327));
    Span4Mux_h I__6776 (
            .O(N__36330),
            .I(N__36324));
    Sp12to4 I__6775 (
            .O(N__36327),
            .I(N__36321));
    Odrv4 I__6774 (
            .O(N__36324),
            .I(comm_buf_2_6));
    Odrv12 I__6773 (
            .O(N__36321),
            .I(comm_buf_2_6));
    InMux I__6772 (
            .O(N__36316),
            .I(N__36313));
    LocalMux I__6771 (
            .O(N__36313),
            .I(n22669));
    InMux I__6770 (
            .O(N__36310),
            .I(N__36307));
    LocalMux I__6769 (
            .O(N__36307),
            .I(N__36304));
    Odrv4 I__6768 (
            .O(N__36304),
            .I(n1_adj_1668));
    InMux I__6767 (
            .O(N__36301),
            .I(N__36298));
    LocalMux I__6766 (
            .O(N__36298),
            .I(n13219));
    InMux I__6765 (
            .O(N__36295),
            .I(N__36289));
    InMux I__6764 (
            .O(N__36294),
            .I(N__36289));
    LocalMux I__6763 (
            .O(N__36289),
            .I(N__36286));
    Span4Mux_v I__6762 (
            .O(N__36286),
            .I(N__36282));
    InMux I__6761 (
            .O(N__36285),
            .I(N__36279));
    Odrv4 I__6760 (
            .O(N__36282),
            .I(comm_tx_buf_4));
    LocalMux I__6759 (
            .O(N__36279),
            .I(comm_tx_buf_4));
    SRMux I__6758 (
            .O(N__36274),
            .I(N__36271));
    LocalMux I__6757 (
            .O(N__36271),
            .I(N__36268));
    Span4Mux_v I__6756 (
            .O(N__36268),
            .I(N__36265));
    Odrv4 I__6755 (
            .O(N__36265),
            .I(\comm_spi.data_tx_7__N_871 ));
    InMux I__6754 (
            .O(N__36262),
            .I(N__36259));
    LocalMux I__6753 (
            .O(N__36259),
            .I(N__36256));
    Odrv12 I__6752 (
            .O(N__36256),
            .I(comm_buf_0_7_N_543_4));
    InMux I__6751 (
            .O(N__36253),
            .I(N__36250));
    LocalMux I__6750 (
            .O(N__36250),
            .I(N__36247));
    Span4Mux_h I__6749 (
            .O(N__36247),
            .I(N__36244));
    Odrv4 I__6748 (
            .O(N__36244),
            .I(comm_buf_0_7_N_543_6));
    CascadeMux I__6747 (
            .O(N__36241),
            .I(\comm_spi.n24034_cascade_ ));
    InMux I__6746 (
            .O(N__36238),
            .I(N__36235));
    LocalMux I__6745 (
            .O(N__36235),
            .I(N__36232));
    Span4Mux_h I__6744 (
            .O(N__36232),
            .I(N__36228));
    InMux I__6743 (
            .O(N__36231),
            .I(N__36225));
    Span4Mux_h I__6742 (
            .O(N__36228),
            .I(N__36222));
    LocalMux I__6741 (
            .O(N__36225),
            .I(N__36219));
    Odrv4 I__6740 (
            .O(N__36222),
            .I(\comm_spi.n15356 ));
    Odrv4 I__6739 (
            .O(N__36219),
            .I(\comm_spi.n15356 ));
    SRMux I__6738 (
            .O(N__36214),
            .I(N__36211));
    LocalMux I__6737 (
            .O(N__36211),
            .I(N__36208));
    Span4Mux_h I__6736 (
            .O(N__36208),
            .I(N__36205));
    Odrv4 I__6735 (
            .O(N__36205),
            .I(\comm_spi.data_tx_7__N_858 ));
    InMux I__6734 (
            .O(N__36202),
            .I(N__36195));
    InMux I__6733 (
            .O(N__36201),
            .I(N__36195));
    InMux I__6732 (
            .O(N__36200),
            .I(N__36192));
    LocalMux I__6731 (
            .O(N__36195),
            .I(comm_tx_buf_6));
    LocalMux I__6730 (
            .O(N__36192),
            .I(comm_tx_buf_6));
    CascadeMux I__6729 (
            .O(N__36187),
            .I(N__36184));
    InMux I__6728 (
            .O(N__36184),
            .I(N__36180));
    InMux I__6727 (
            .O(N__36183),
            .I(N__36177));
    LocalMux I__6726 (
            .O(N__36180),
            .I(N__36172));
    LocalMux I__6725 (
            .O(N__36177),
            .I(N__36172));
    Span4Mux_v I__6724 (
            .O(N__36172),
            .I(N__36169));
    Span4Mux_v I__6723 (
            .O(N__36169),
            .I(N__36165));
    InMux I__6722 (
            .O(N__36168),
            .I(N__36162));
    Odrv4 I__6721 (
            .O(N__36165),
            .I(\comm_spi.n24013 ));
    LocalMux I__6720 (
            .O(N__36162),
            .I(\comm_spi.n24013 ));
    SRMux I__6719 (
            .O(N__36157),
            .I(N__36154));
    LocalMux I__6718 (
            .O(N__36154),
            .I(N__36151));
    Span4Mux_v I__6717 (
            .O(N__36151),
            .I(N__36148));
    Span4Mux_h I__6716 (
            .O(N__36148),
            .I(N__36145));
    Odrv4 I__6715 (
            .O(N__36145),
            .I(\comm_spi.data_tx_7__N_856 ));
    CascadeMux I__6714 (
            .O(N__36142),
            .I(n2_adj_1669_cascade_));
    CascadeMux I__6713 (
            .O(N__36139),
            .I(n4_adj_1670_cascade_));
    InMux I__6712 (
            .O(N__36136),
            .I(N__36133));
    LocalMux I__6711 (
            .O(N__36133),
            .I(n23402));
    CascadeMux I__6710 (
            .O(N__36130),
            .I(n19_adj_1706_cascade_));
    CascadeMux I__6709 (
            .O(N__36127),
            .I(N__36123));
    CascadeMux I__6708 (
            .O(N__36126),
            .I(N__36120));
    InMux I__6707 (
            .O(N__36123),
            .I(N__36117));
    InMux I__6706 (
            .O(N__36120),
            .I(N__36114));
    LocalMux I__6705 (
            .O(N__36117),
            .I(N__36110));
    LocalMux I__6704 (
            .O(N__36114),
            .I(N__36107));
    InMux I__6703 (
            .O(N__36113),
            .I(N__36104));
    Span4Mux_v I__6702 (
            .O(N__36110),
            .I(N__36101));
    Odrv4 I__6701 (
            .O(N__36107),
            .I(cmd_rdadctmp_8_adj_1540));
    LocalMux I__6700 (
            .O(N__36104),
            .I(cmd_rdadctmp_8_adj_1540));
    Odrv4 I__6699 (
            .O(N__36101),
            .I(cmd_rdadctmp_8_adj_1540));
    InMux I__6698 (
            .O(N__36094),
            .I(N__36090));
    CascadeMux I__6697 (
            .O(N__36093),
            .I(N__36087));
    LocalMux I__6696 (
            .O(N__36090),
            .I(N__36083));
    InMux I__6695 (
            .O(N__36087),
            .I(N__36080));
    InMux I__6694 (
            .O(N__36086),
            .I(N__36077));
    Span12Mux_h I__6693 (
            .O(N__36083),
            .I(N__36074));
    LocalMux I__6692 (
            .O(N__36080),
            .I(buf_adcdata_iac_1));
    LocalMux I__6691 (
            .O(N__36077),
            .I(buf_adcdata_iac_1));
    Odrv12 I__6690 (
            .O(N__36074),
            .I(buf_adcdata_iac_1));
    InMux I__6689 (
            .O(N__36067),
            .I(N__36064));
    LocalMux I__6688 (
            .O(N__36064),
            .I(N__36061));
    Span4Mux_v I__6687 (
            .O(N__36061),
            .I(N__36058));
    Sp12to4 I__6686 (
            .O(N__36058),
            .I(N__36053));
    InMux I__6685 (
            .O(N__36057),
            .I(N__36048));
    InMux I__6684 (
            .O(N__36056),
            .I(N__36048));
    Odrv12 I__6683 (
            .O(N__36053),
            .I(buf_adcdata_iac_2));
    LocalMux I__6682 (
            .O(N__36048),
            .I(buf_adcdata_iac_2));
    CascadeMux I__6681 (
            .O(N__36043),
            .I(N__36040));
    InMux I__6680 (
            .O(N__36040),
            .I(N__36037));
    LocalMux I__6679 (
            .O(N__36037),
            .I(N__36034));
    Span4Mux_h I__6678 (
            .O(N__36034),
            .I(N__36030));
    InMux I__6677 (
            .O(N__36033),
            .I(N__36026));
    Span4Mux_h I__6676 (
            .O(N__36030),
            .I(N__36023));
    InMux I__6675 (
            .O(N__36029),
            .I(N__36020));
    LocalMux I__6674 (
            .O(N__36026),
            .I(cmd_rdadctmp_10_adj_1538));
    Odrv4 I__6673 (
            .O(N__36023),
            .I(cmd_rdadctmp_10_adj_1538));
    LocalMux I__6672 (
            .O(N__36020),
            .I(cmd_rdadctmp_10_adj_1538));
    InMux I__6671 (
            .O(N__36013),
            .I(N__35994));
    InMux I__6670 (
            .O(N__36012),
            .I(N__35977));
    InMux I__6669 (
            .O(N__36011),
            .I(N__35977));
    InMux I__6668 (
            .O(N__36010),
            .I(N__35977));
    InMux I__6667 (
            .O(N__36009),
            .I(N__35977));
    InMux I__6666 (
            .O(N__36008),
            .I(N__35977));
    InMux I__6665 (
            .O(N__36007),
            .I(N__35966));
    InMux I__6664 (
            .O(N__36006),
            .I(N__35966));
    InMux I__6663 (
            .O(N__36005),
            .I(N__35966));
    InMux I__6662 (
            .O(N__36004),
            .I(N__35966));
    InMux I__6661 (
            .O(N__36003),
            .I(N__35966));
    InMux I__6660 (
            .O(N__36002),
            .I(N__35959));
    InMux I__6659 (
            .O(N__36001),
            .I(N__35947));
    InMux I__6658 (
            .O(N__36000),
            .I(N__35947));
    InMux I__6657 (
            .O(N__35999),
            .I(N__35947));
    InMux I__6656 (
            .O(N__35998),
            .I(N__35947));
    InMux I__6655 (
            .O(N__35997),
            .I(N__35947));
    LocalMux I__6654 (
            .O(N__35994),
            .I(N__35943));
    InMux I__6653 (
            .O(N__35993),
            .I(N__35938));
    InMux I__6652 (
            .O(N__35992),
            .I(N__35938));
    InMux I__6651 (
            .O(N__35991),
            .I(N__35933));
    InMux I__6650 (
            .O(N__35990),
            .I(N__35933));
    CascadeMux I__6649 (
            .O(N__35989),
            .I(N__35930));
    InMux I__6648 (
            .O(N__35988),
            .I(N__35918));
    LocalMux I__6647 (
            .O(N__35977),
            .I(N__35904));
    LocalMux I__6646 (
            .O(N__35966),
            .I(N__35904));
    InMux I__6645 (
            .O(N__35965),
            .I(N__35899));
    InMux I__6644 (
            .O(N__35964),
            .I(N__35899));
    InMux I__6643 (
            .O(N__35963),
            .I(N__35891));
    InMux I__6642 (
            .O(N__35962),
            .I(N__35891));
    LocalMux I__6641 (
            .O(N__35959),
            .I(N__35888));
    InMux I__6640 (
            .O(N__35958),
            .I(N__35885));
    LocalMux I__6639 (
            .O(N__35947),
            .I(N__35882));
    InMux I__6638 (
            .O(N__35946),
            .I(N__35878));
    Span4Mux_v I__6637 (
            .O(N__35943),
            .I(N__35875));
    LocalMux I__6636 (
            .O(N__35938),
            .I(N__35872));
    LocalMux I__6635 (
            .O(N__35933),
            .I(N__35869));
    InMux I__6634 (
            .O(N__35930),
            .I(N__35860));
    InMux I__6633 (
            .O(N__35929),
            .I(N__35860));
    InMux I__6632 (
            .O(N__35928),
            .I(N__35855));
    InMux I__6631 (
            .O(N__35927),
            .I(N__35855));
    InMux I__6630 (
            .O(N__35926),
            .I(N__35851));
    InMux I__6629 (
            .O(N__35925),
            .I(N__35846));
    InMux I__6628 (
            .O(N__35924),
            .I(N__35846));
    InMux I__6627 (
            .O(N__35923),
            .I(N__35843));
    InMux I__6626 (
            .O(N__35922),
            .I(N__35838));
    InMux I__6625 (
            .O(N__35921),
            .I(N__35838));
    LocalMux I__6624 (
            .O(N__35918),
            .I(N__35835));
    InMux I__6623 (
            .O(N__35917),
            .I(N__35826));
    InMux I__6622 (
            .O(N__35916),
            .I(N__35826));
    InMux I__6621 (
            .O(N__35915),
            .I(N__35826));
    InMux I__6620 (
            .O(N__35914),
            .I(N__35826));
    InMux I__6619 (
            .O(N__35913),
            .I(N__35819));
    InMux I__6618 (
            .O(N__35912),
            .I(N__35819));
    InMux I__6617 (
            .O(N__35911),
            .I(N__35819));
    InMux I__6616 (
            .O(N__35910),
            .I(N__35814));
    InMux I__6615 (
            .O(N__35909),
            .I(N__35814));
    Span4Mux_v I__6614 (
            .O(N__35904),
            .I(N__35809));
    LocalMux I__6613 (
            .O(N__35899),
            .I(N__35809));
    InMux I__6612 (
            .O(N__35898),
            .I(N__35802));
    InMux I__6611 (
            .O(N__35897),
            .I(N__35802));
    InMux I__6610 (
            .O(N__35896),
            .I(N__35802));
    LocalMux I__6609 (
            .O(N__35891),
            .I(N__35799));
    Span4Mux_v I__6608 (
            .O(N__35888),
            .I(N__35792));
    LocalMux I__6607 (
            .O(N__35885),
            .I(N__35792));
    Span4Mux_h I__6606 (
            .O(N__35882),
            .I(N__35792));
    InMux I__6605 (
            .O(N__35881),
            .I(N__35789));
    LocalMux I__6604 (
            .O(N__35878),
            .I(N__35786));
    Span4Mux_h I__6603 (
            .O(N__35875),
            .I(N__35779));
    Span4Mux_v I__6602 (
            .O(N__35872),
            .I(N__35779));
    Span4Mux_h I__6601 (
            .O(N__35869),
            .I(N__35779));
    InMux I__6600 (
            .O(N__35868),
            .I(N__35771));
    InMux I__6599 (
            .O(N__35867),
            .I(N__35768));
    InMux I__6598 (
            .O(N__35866),
            .I(N__35763));
    InMux I__6597 (
            .O(N__35865),
            .I(N__35763));
    LocalMux I__6596 (
            .O(N__35860),
            .I(N__35758));
    LocalMux I__6595 (
            .O(N__35855),
            .I(N__35758));
    InMux I__6594 (
            .O(N__35854),
            .I(N__35755));
    LocalMux I__6593 (
            .O(N__35851),
            .I(N__35748));
    LocalMux I__6592 (
            .O(N__35846),
            .I(N__35748));
    LocalMux I__6591 (
            .O(N__35843),
            .I(N__35748));
    LocalMux I__6590 (
            .O(N__35838),
            .I(N__35745));
    Span4Mux_h I__6589 (
            .O(N__35835),
            .I(N__35740));
    LocalMux I__6588 (
            .O(N__35826),
            .I(N__35740));
    LocalMux I__6587 (
            .O(N__35819),
            .I(N__35737));
    LocalMux I__6586 (
            .O(N__35814),
            .I(N__35730));
    Span4Mux_h I__6585 (
            .O(N__35809),
            .I(N__35730));
    LocalMux I__6584 (
            .O(N__35802),
            .I(N__35730));
    Span4Mux_v I__6583 (
            .O(N__35799),
            .I(N__35727));
    Span4Mux_v I__6582 (
            .O(N__35792),
            .I(N__35724));
    LocalMux I__6581 (
            .O(N__35789),
            .I(N__35717));
    Span4Mux_h I__6580 (
            .O(N__35786),
            .I(N__35717));
    Span4Mux_h I__6579 (
            .O(N__35779),
            .I(N__35717));
    InMux I__6578 (
            .O(N__35778),
            .I(N__35702));
    InMux I__6577 (
            .O(N__35777),
            .I(N__35702));
    InMux I__6576 (
            .O(N__35776),
            .I(N__35702));
    InMux I__6575 (
            .O(N__35775),
            .I(N__35697));
    InMux I__6574 (
            .O(N__35774),
            .I(N__35697));
    LocalMux I__6573 (
            .O(N__35771),
            .I(N__35692));
    LocalMux I__6572 (
            .O(N__35768),
            .I(N__35692));
    LocalMux I__6571 (
            .O(N__35763),
            .I(N__35687));
    Span12Mux_h I__6570 (
            .O(N__35758),
            .I(N__35687));
    LocalMux I__6569 (
            .O(N__35755),
            .I(N__35670));
    Span4Mux_v I__6568 (
            .O(N__35748),
            .I(N__35670));
    Span4Mux_v I__6567 (
            .O(N__35745),
            .I(N__35670));
    Span4Mux_v I__6566 (
            .O(N__35740),
            .I(N__35670));
    Span4Mux_v I__6565 (
            .O(N__35737),
            .I(N__35670));
    Span4Mux_v I__6564 (
            .O(N__35730),
            .I(N__35670));
    Span4Mux_h I__6563 (
            .O(N__35727),
            .I(N__35670));
    Span4Mux_h I__6562 (
            .O(N__35724),
            .I(N__35670));
    Span4Mux_v I__6561 (
            .O(N__35717),
            .I(N__35667));
    InMux I__6560 (
            .O(N__35716),
            .I(N__35662));
    InMux I__6559 (
            .O(N__35715),
            .I(N__35662));
    InMux I__6558 (
            .O(N__35714),
            .I(N__35653));
    InMux I__6557 (
            .O(N__35713),
            .I(N__35653));
    InMux I__6556 (
            .O(N__35712),
            .I(N__35653));
    InMux I__6555 (
            .O(N__35711),
            .I(N__35653));
    InMux I__6554 (
            .O(N__35710),
            .I(N__35648));
    InMux I__6553 (
            .O(N__35709),
            .I(N__35648));
    LocalMux I__6552 (
            .O(N__35702),
            .I(adc_state_0_adj_1516));
    LocalMux I__6551 (
            .O(N__35697),
            .I(adc_state_0_adj_1516));
    Odrv4 I__6550 (
            .O(N__35692),
            .I(adc_state_0_adj_1516));
    Odrv12 I__6549 (
            .O(N__35687),
            .I(adc_state_0_adj_1516));
    Odrv4 I__6548 (
            .O(N__35670),
            .I(adc_state_0_adj_1516));
    Odrv4 I__6547 (
            .O(N__35667),
            .I(adc_state_0_adj_1516));
    LocalMux I__6546 (
            .O(N__35662),
            .I(adc_state_0_adj_1516));
    LocalMux I__6545 (
            .O(N__35653),
            .I(adc_state_0_adj_1516));
    LocalMux I__6544 (
            .O(N__35648),
            .I(adc_state_0_adj_1516));
    CascadeMux I__6543 (
            .O(N__35629),
            .I(N__35626));
    InMux I__6542 (
            .O(N__35626),
            .I(N__35618));
    InMux I__6541 (
            .O(N__35625),
            .I(N__35618));
    InMux I__6540 (
            .O(N__35624),
            .I(N__35611));
    InMux I__6539 (
            .O(N__35623),
            .I(N__35611));
    LocalMux I__6538 (
            .O(N__35618),
            .I(N__35604));
    InMux I__6537 (
            .O(N__35617),
            .I(N__35591));
    InMux I__6536 (
            .O(N__35616),
            .I(N__35591));
    LocalMux I__6535 (
            .O(N__35611),
            .I(N__35588));
    InMux I__6534 (
            .O(N__35610),
            .I(N__35584));
    InMux I__6533 (
            .O(N__35609),
            .I(N__35581));
    InMux I__6532 (
            .O(N__35608),
            .I(N__35578));
    InMux I__6531 (
            .O(N__35607),
            .I(N__35575));
    Span4Mux_v I__6530 (
            .O(N__35604),
            .I(N__35572));
    InMux I__6529 (
            .O(N__35603),
            .I(N__35568));
    InMux I__6528 (
            .O(N__35602),
            .I(N__35562));
    InMux I__6527 (
            .O(N__35601),
            .I(N__35559));
    InMux I__6526 (
            .O(N__35600),
            .I(N__35552));
    InMux I__6525 (
            .O(N__35599),
            .I(N__35552));
    InMux I__6524 (
            .O(N__35598),
            .I(N__35552));
    InMux I__6523 (
            .O(N__35597),
            .I(N__35547));
    InMux I__6522 (
            .O(N__35596),
            .I(N__35547));
    LocalMux I__6521 (
            .O(N__35591),
            .I(N__35542));
    Span4Mux_v I__6520 (
            .O(N__35588),
            .I(N__35542));
    InMux I__6519 (
            .O(N__35587),
            .I(N__35539));
    LocalMux I__6518 (
            .O(N__35584),
            .I(N__35534));
    LocalMux I__6517 (
            .O(N__35581),
            .I(N__35534));
    LocalMux I__6516 (
            .O(N__35578),
            .I(N__35531));
    LocalMux I__6515 (
            .O(N__35575),
            .I(N__35526));
    Span4Mux_h I__6514 (
            .O(N__35572),
            .I(N__35526));
    CascadeMux I__6513 (
            .O(N__35571),
            .I(N__35523));
    LocalMux I__6512 (
            .O(N__35568),
            .I(N__35520));
    InMux I__6511 (
            .O(N__35567),
            .I(N__35517));
    InMux I__6510 (
            .O(N__35566),
            .I(N__35512));
    InMux I__6509 (
            .O(N__35565),
            .I(N__35512));
    LocalMux I__6508 (
            .O(N__35562),
            .I(N__35507));
    LocalMux I__6507 (
            .O(N__35559),
            .I(N__35507));
    LocalMux I__6506 (
            .O(N__35552),
            .I(N__35504));
    LocalMux I__6505 (
            .O(N__35547),
            .I(N__35499));
    Span4Mux_h I__6504 (
            .O(N__35542),
            .I(N__35499));
    LocalMux I__6503 (
            .O(N__35539),
            .I(N__35494));
    Span4Mux_v I__6502 (
            .O(N__35534),
            .I(N__35494));
    Span4Mux_v I__6501 (
            .O(N__35531),
            .I(N__35489));
    Span4Mux_v I__6500 (
            .O(N__35526),
            .I(N__35489));
    InMux I__6499 (
            .O(N__35523),
            .I(N__35486));
    Span4Mux_h I__6498 (
            .O(N__35520),
            .I(N__35483));
    LocalMux I__6497 (
            .O(N__35517),
            .I(N__35472));
    LocalMux I__6496 (
            .O(N__35512),
            .I(N__35472));
    Span4Mux_h I__6495 (
            .O(N__35507),
            .I(N__35472));
    Span4Mux_v I__6494 (
            .O(N__35504),
            .I(N__35472));
    Span4Mux_h I__6493 (
            .O(N__35499),
            .I(N__35472));
    Span4Mux_v I__6492 (
            .O(N__35494),
            .I(N__35467));
    Span4Mux_h I__6491 (
            .O(N__35489),
            .I(N__35467));
    LocalMux I__6490 (
            .O(N__35486),
            .I(n21948));
    Odrv4 I__6489 (
            .O(N__35483),
            .I(n21948));
    Odrv4 I__6488 (
            .O(N__35472),
            .I(n21948));
    Odrv4 I__6487 (
            .O(N__35467),
            .I(n21948));
    InMux I__6486 (
            .O(N__35458),
            .I(N__35455));
    LocalMux I__6485 (
            .O(N__35455),
            .I(N__35452));
    Span4Mux_v I__6484 (
            .O(N__35452),
            .I(N__35449));
    Sp12to4 I__6483 (
            .O(N__35449),
            .I(N__35444));
    InMux I__6482 (
            .O(N__35448),
            .I(N__35439));
    InMux I__6481 (
            .O(N__35447),
            .I(N__35439));
    Odrv12 I__6480 (
            .O(N__35444),
            .I(buf_adcdata_vac_2));
    LocalMux I__6479 (
            .O(N__35439),
            .I(buf_adcdata_vac_2));
    CascadeMux I__6478 (
            .O(N__35434),
            .I(N__35430));
    InMux I__6477 (
            .O(N__35433),
            .I(N__35425));
    InMux I__6476 (
            .O(N__35430),
            .I(N__35425));
    LocalMux I__6475 (
            .O(N__35425),
            .I(N__35422));
    Span4Mux_v I__6474 (
            .O(N__35422),
            .I(N__35418));
    InMux I__6473 (
            .O(N__35421),
            .I(N__35415));
    Odrv4 I__6472 (
            .O(N__35418),
            .I(cmd_rdadctmp_9));
    LocalMux I__6471 (
            .O(N__35415),
            .I(cmd_rdadctmp_9));
    CascadeMux I__6470 (
            .O(N__35410),
            .I(N__35406));
    InMux I__6469 (
            .O(N__35409),
            .I(N__35398));
    InMux I__6468 (
            .O(N__35406),
            .I(N__35398));
    InMux I__6467 (
            .O(N__35405),
            .I(N__35398));
    LocalMux I__6466 (
            .O(N__35398),
            .I(cmd_rdadctmp_10));
    CascadeMux I__6465 (
            .O(N__35395),
            .I(N__35392));
    InMux I__6464 (
            .O(N__35392),
            .I(N__35389));
    LocalMux I__6463 (
            .O(N__35389),
            .I(N__35385));
    CascadeMux I__6462 (
            .O(N__35388),
            .I(N__35382));
    Span4Mux_v I__6461 (
            .O(N__35385),
            .I(N__35379));
    InMux I__6460 (
            .O(N__35382),
            .I(N__35375));
    Span4Mux_h I__6459 (
            .O(N__35379),
            .I(N__35372));
    InMux I__6458 (
            .O(N__35378),
            .I(N__35369));
    LocalMux I__6457 (
            .O(N__35375),
            .I(cmd_rdadctmp_11));
    Odrv4 I__6456 (
            .O(N__35372),
            .I(cmd_rdadctmp_11));
    LocalMux I__6455 (
            .O(N__35369),
            .I(cmd_rdadctmp_11));
    CascadeMux I__6454 (
            .O(N__35362),
            .I(N__35359));
    InMux I__6453 (
            .O(N__35359),
            .I(N__35356));
    LocalMux I__6452 (
            .O(N__35356),
            .I(N__35351));
    InMux I__6451 (
            .O(N__35355),
            .I(N__35348));
    CascadeMux I__6450 (
            .O(N__35354),
            .I(N__35345));
    Span4Mux_v I__6449 (
            .O(N__35351),
            .I(N__35341));
    LocalMux I__6448 (
            .O(N__35348),
            .I(N__35338));
    InMux I__6447 (
            .O(N__35345),
            .I(N__35334));
    InMux I__6446 (
            .O(N__35344),
            .I(N__35331));
    Span4Mux_h I__6445 (
            .O(N__35341),
            .I(N__35326));
    Span4Mux_v I__6444 (
            .O(N__35338),
            .I(N__35326));
    InMux I__6443 (
            .O(N__35337),
            .I(N__35323));
    LocalMux I__6442 (
            .O(N__35334),
            .I(N__35318));
    LocalMux I__6441 (
            .O(N__35331),
            .I(N__35318));
    Odrv4 I__6440 (
            .O(N__35326),
            .I(buf_cfgRTD_7));
    LocalMux I__6439 (
            .O(N__35323),
            .I(buf_cfgRTD_7));
    Odrv12 I__6438 (
            .O(N__35318),
            .I(buf_cfgRTD_7));
    CascadeMux I__6437 (
            .O(N__35311),
            .I(N__35308));
    InMux I__6436 (
            .O(N__35308),
            .I(N__35305));
    LocalMux I__6435 (
            .O(N__35305),
            .I(N__35302));
    Span4Mux_h I__6434 (
            .O(N__35302),
            .I(N__35299));
    Span4Mux_h I__6433 (
            .O(N__35299),
            .I(N__35295));
    InMux I__6432 (
            .O(N__35298),
            .I(N__35292));
    Odrv4 I__6431 (
            .O(N__35295),
            .I(buf_readRTD_15));
    LocalMux I__6430 (
            .O(N__35292),
            .I(buf_readRTD_15));
    InMux I__6429 (
            .O(N__35287),
            .I(N__35284));
    LocalMux I__6428 (
            .O(N__35284),
            .I(N__35281));
    Span4Mux_h I__6427 (
            .O(N__35281),
            .I(N__35278));
    Odrv4 I__6426 (
            .O(N__35278),
            .I(n23432));
    CascadeMux I__6425 (
            .O(N__35275),
            .I(n12610_cascade_));
    SRMux I__6424 (
            .O(N__35272),
            .I(N__35269));
    LocalMux I__6423 (
            .O(N__35269),
            .I(N__35266));
    Span4Mux_h I__6422 (
            .O(N__35266),
            .I(N__35263));
    Span4Mux_h I__6421 (
            .O(N__35263),
            .I(N__35260));
    Odrv4 I__6420 (
            .O(N__35260),
            .I(\comm_spi.data_tx_7__N_883 ));
    IoInMux I__6419 (
            .O(N__35257),
            .I(N__35254));
    LocalMux I__6418 (
            .O(N__35254),
            .I(N__35251));
    Span4Mux_s3_h I__6417 (
            .O(N__35251),
            .I(N__35248));
    Span4Mux_v I__6416 (
            .O(N__35248),
            .I(N__35245));
    Sp12to4 I__6415 (
            .O(N__35245),
            .I(N__35242));
    Span12Mux_h I__6414 (
            .O(N__35242),
            .I(N__35239));
    Odrv12 I__6413 (
            .O(N__35239),
            .I(ICE_SPI_MISO));
    SRMux I__6412 (
            .O(N__35236),
            .I(N__35233));
    LocalMux I__6411 (
            .O(N__35233),
            .I(N__35230));
    Span4Mux_h I__6410 (
            .O(N__35230),
            .I(N__35227));
    Span4Mux_h I__6409 (
            .O(N__35227),
            .I(N__35224));
    Odrv4 I__6408 (
            .O(N__35224),
            .I(\comm_spi.data_tx_7__N_868 ));
    InMux I__6407 (
            .O(N__35221),
            .I(N__35218));
    LocalMux I__6406 (
            .O(N__35218),
            .I(N__35215));
    Span4Mux_h I__6405 (
            .O(N__35215),
            .I(N__35211));
    CascadeMux I__6404 (
            .O(N__35214),
            .I(N__35208));
    Span4Mux_v I__6403 (
            .O(N__35211),
            .I(N__35205));
    InMux I__6402 (
            .O(N__35208),
            .I(N__35202));
    Odrv4 I__6401 (
            .O(N__35205),
            .I(buf_adcdata_vdc_2));
    LocalMux I__6400 (
            .O(N__35202),
            .I(buf_adcdata_vdc_2));
    InMux I__6399 (
            .O(N__35197),
            .I(n20649));
    InMux I__6398 (
            .O(N__35194),
            .I(n20650));
    InMux I__6397 (
            .O(N__35191),
            .I(n20651));
    CEMux I__6396 (
            .O(N__35188),
            .I(N__35184));
    CEMux I__6395 (
            .O(N__35187),
            .I(N__35181));
    LocalMux I__6394 (
            .O(N__35184),
            .I(N__35178));
    LocalMux I__6393 (
            .O(N__35181),
            .I(N__35175));
    Span4Mux_v I__6392 (
            .O(N__35178),
            .I(N__35172));
    Span4Mux_v I__6391 (
            .O(N__35175),
            .I(N__35168));
    Span4Mux_h I__6390 (
            .O(N__35172),
            .I(N__35165));
    CEMux I__6389 (
            .O(N__35171),
            .I(N__35162));
    Odrv4 I__6388 (
            .O(N__35168),
            .I(n12450));
    Odrv4 I__6387 (
            .O(N__35165),
            .I(n12450));
    LocalMux I__6386 (
            .O(N__35162),
            .I(n12450));
    SRMux I__6385 (
            .O(N__35155),
            .I(N__35151));
    SRMux I__6384 (
            .O(N__35154),
            .I(N__35148));
    LocalMux I__6383 (
            .O(N__35151),
            .I(N__35145));
    LocalMux I__6382 (
            .O(N__35148),
            .I(N__35142));
    Span4Mux_v I__6381 (
            .O(N__35145),
            .I(N__35139));
    Span4Mux_v I__6380 (
            .O(N__35142),
            .I(N__35136));
    Odrv4 I__6379 (
            .O(N__35139),
            .I(n15439));
    Odrv4 I__6378 (
            .O(N__35136),
            .I(n15439));
    InMux I__6377 (
            .O(N__35131),
            .I(N__35125));
    InMux I__6376 (
            .O(N__35130),
            .I(N__35118));
    InMux I__6375 (
            .O(N__35129),
            .I(N__35118));
    InMux I__6374 (
            .O(N__35128),
            .I(N__35118));
    LocalMux I__6373 (
            .O(N__35125),
            .I(N__35112));
    LocalMux I__6372 (
            .O(N__35118),
            .I(N__35112));
    InMux I__6371 (
            .O(N__35117),
            .I(N__35109));
    Span12Mux_s11_h I__6370 (
            .O(N__35112),
            .I(N__35106));
    LocalMux I__6369 (
            .O(N__35109),
            .I(\RTD.bit_cnt_3 ));
    Odrv12 I__6368 (
            .O(N__35106),
            .I(\RTD.bit_cnt_3 ));
    CascadeMux I__6367 (
            .O(N__35101),
            .I(N__35098));
    InMux I__6366 (
            .O(N__35098),
            .I(N__35091));
    InMux I__6365 (
            .O(N__35097),
            .I(N__35091));
    InMux I__6364 (
            .O(N__35096),
            .I(N__35088));
    LocalMux I__6363 (
            .O(N__35091),
            .I(\RTD.bit_cnt_2 ));
    LocalMux I__6362 (
            .O(N__35088),
            .I(\RTD.bit_cnt_2 ));
    InMux I__6361 (
            .O(N__35083),
            .I(N__35073));
    InMux I__6360 (
            .O(N__35082),
            .I(N__35073));
    InMux I__6359 (
            .O(N__35081),
            .I(N__35073));
    InMux I__6358 (
            .O(N__35080),
            .I(N__35070));
    LocalMux I__6357 (
            .O(N__35073),
            .I(\RTD.bit_cnt_1 ));
    LocalMux I__6356 (
            .O(N__35070),
            .I(\RTD.bit_cnt_1 ));
    InMux I__6355 (
            .O(N__35065),
            .I(N__35052));
    InMux I__6354 (
            .O(N__35064),
            .I(N__35052));
    InMux I__6353 (
            .O(N__35063),
            .I(N__35052));
    InMux I__6352 (
            .O(N__35062),
            .I(N__35052));
    InMux I__6351 (
            .O(N__35061),
            .I(N__35049));
    LocalMux I__6350 (
            .O(N__35052),
            .I(\RTD.bit_cnt_0 ));
    LocalMux I__6349 (
            .O(N__35049),
            .I(\RTD.bit_cnt_0 ));
    ClkMux I__6348 (
            .O(N__35044),
            .I(N__35039));
    ClkMux I__6347 (
            .O(N__35043),
            .I(N__35035));
    ClkMux I__6346 (
            .O(N__35042),
            .I(N__35031));
    LocalMux I__6345 (
            .O(N__35039),
            .I(N__35026));
    ClkMux I__6344 (
            .O(N__35038),
            .I(N__35023));
    LocalMux I__6343 (
            .O(N__35035),
            .I(N__35018));
    ClkMux I__6342 (
            .O(N__35034),
            .I(N__35015));
    LocalMux I__6341 (
            .O(N__35031),
            .I(N__35010));
    ClkMux I__6340 (
            .O(N__35030),
            .I(N__35007));
    ClkMux I__6339 (
            .O(N__35029),
            .I(N__35003));
    Span4Mux_h I__6338 (
            .O(N__35026),
            .I(N__34995));
    LocalMux I__6337 (
            .O(N__35023),
            .I(N__34995));
    ClkMux I__6336 (
            .O(N__35022),
            .I(N__34992));
    ClkMux I__6335 (
            .O(N__35021),
            .I(N__34989));
    Span4Mux_v I__6334 (
            .O(N__35018),
            .I(N__34984));
    LocalMux I__6333 (
            .O(N__35015),
            .I(N__34984));
    ClkMux I__6332 (
            .O(N__35014),
            .I(N__34981));
    ClkMux I__6331 (
            .O(N__35013),
            .I(N__34977));
    Span4Mux_h I__6330 (
            .O(N__35010),
            .I(N__34972));
    LocalMux I__6329 (
            .O(N__35007),
            .I(N__34972));
    ClkMux I__6328 (
            .O(N__35006),
            .I(N__34969));
    LocalMux I__6327 (
            .O(N__35003),
            .I(N__34966));
    ClkMux I__6326 (
            .O(N__35002),
            .I(N__34963));
    ClkMux I__6325 (
            .O(N__35001),
            .I(N__34960));
    ClkMux I__6324 (
            .O(N__35000),
            .I(N__34957));
    Span4Mux_v I__6323 (
            .O(N__34995),
            .I(N__34953));
    LocalMux I__6322 (
            .O(N__34992),
            .I(N__34948));
    LocalMux I__6321 (
            .O(N__34989),
            .I(N__34948));
    Span4Mux_v I__6320 (
            .O(N__34984),
            .I(N__34943));
    LocalMux I__6319 (
            .O(N__34981),
            .I(N__34943));
    ClkMux I__6318 (
            .O(N__34980),
            .I(N__34940));
    LocalMux I__6317 (
            .O(N__34977),
            .I(N__34937));
    Span4Mux_v I__6316 (
            .O(N__34972),
            .I(N__34932));
    LocalMux I__6315 (
            .O(N__34969),
            .I(N__34932));
    Span4Mux_h I__6314 (
            .O(N__34966),
            .I(N__34927));
    LocalMux I__6313 (
            .O(N__34963),
            .I(N__34927));
    LocalMux I__6312 (
            .O(N__34960),
            .I(N__34924));
    LocalMux I__6311 (
            .O(N__34957),
            .I(N__34921));
    ClkMux I__6310 (
            .O(N__34956),
            .I(N__34918));
    Span4Mux_h I__6309 (
            .O(N__34953),
            .I(N__34909));
    Span4Mux_v I__6308 (
            .O(N__34948),
            .I(N__34909));
    Span4Mux_v I__6307 (
            .O(N__34943),
            .I(N__34909));
    LocalMux I__6306 (
            .O(N__34940),
            .I(N__34909));
    Span4Mux_v I__6305 (
            .O(N__34937),
            .I(N__34902));
    Span4Mux_h I__6304 (
            .O(N__34932),
            .I(N__34902));
    Span4Mux_v I__6303 (
            .O(N__34927),
            .I(N__34902));
    Span4Mux_v I__6302 (
            .O(N__34924),
            .I(N__34895));
    Span4Mux_v I__6301 (
            .O(N__34921),
            .I(N__34895));
    LocalMux I__6300 (
            .O(N__34918),
            .I(N__34895));
    Span4Mux_h I__6299 (
            .O(N__34909),
            .I(N__34892));
    Span4Mux_h I__6298 (
            .O(N__34902),
            .I(N__34887));
    Span4Mux_v I__6297 (
            .O(N__34895),
            .I(N__34887));
    Span4Mux_h I__6296 (
            .O(N__34892),
            .I(N__34882));
    Span4Mux_h I__6295 (
            .O(N__34887),
            .I(N__34879));
    ClkMux I__6294 (
            .O(N__34886),
            .I(N__34876));
    InMux I__6293 (
            .O(N__34885),
            .I(N__34873));
    Odrv4 I__6292 (
            .O(N__34882),
            .I(clk_RTD));
    Odrv4 I__6291 (
            .O(N__34879),
            .I(clk_RTD));
    LocalMux I__6290 (
            .O(N__34876),
            .I(clk_RTD));
    LocalMux I__6289 (
            .O(N__34873),
            .I(clk_RTD));
    CEMux I__6288 (
            .O(N__34864),
            .I(N__34861));
    LocalMux I__6287 (
            .O(N__34861),
            .I(N__34858));
    Span4Mux_h I__6286 (
            .O(N__34858),
            .I(N__34855));
    Odrv4 I__6285 (
            .O(N__34855),
            .I(\RTD.n18274 ));
    SRMux I__6284 (
            .O(N__34852),
            .I(N__34849));
    LocalMux I__6283 (
            .O(N__34849),
            .I(N__34846));
    Span4Mux_h I__6282 (
            .O(N__34846),
            .I(N__34843));
    Odrv4 I__6281 (
            .O(N__34843),
            .I(\RTD.n18275 ));
    InMux I__6280 (
            .O(N__34840),
            .I(n20640));
    InMux I__6279 (
            .O(N__34837),
            .I(n20641));
    InMux I__6278 (
            .O(N__34834),
            .I(n20642));
    InMux I__6277 (
            .O(N__34831),
            .I(n20643));
    InMux I__6276 (
            .O(N__34828),
            .I(n20644));
    InMux I__6275 (
            .O(N__34825),
            .I(bfn_11_20_0_));
    InMux I__6274 (
            .O(N__34822),
            .I(n20646));
    InMux I__6273 (
            .O(N__34819),
            .I(n20647));
    InMux I__6272 (
            .O(N__34816),
            .I(n20648));
    InMux I__6271 (
            .O(N__34813),
            .I(bfn_11_19_0_));
    InMux I__6270 (
            .O(N__34810),
            .I(n20638));
    InMux I__6269 (
            .O(N__34807),
            .I(n20639));
    InMux I__6268 (
            .O(N__34804),
            .I(N__34801));
    LocalMux I__6267 (
            .O(N__34801),
            .I(n11980));
    CascadeMux I__6266 (
            .O(N__34798),
            .I(N__34792));
    CascadeMux I__6265 (
            .O(N__34797),
            .I(N__34788));
    CascadeMux I__6264 (
            .O(N__34796),
            .I(N__34778));
    CascadeMux I__6263 (
            .O(N__34795),
            .I(N__34775));
    InMux I__6262 (
            .O(N__34792),
            .I(N__34771));
    CascadeMux I__6261 (
            .O(N__34791),
            .I(N__34768));
    InMux I__6260 (
            .O(N__34788),
            .I(N__34765));
    CascadeMux I__6259 (
            .O(N__34787),
            .I(N__34762));
    CascadeMux I__6258 (
            .O(N__34786),
            .I(N__34759));
    CascadeMux I__6257 (
            .O(N__34785),
            .I(N__34756));
    InMux I__6256 (
            .O(N__34784),
            .I(N__34751));
    InMux I__6255 (
            .O(N__34783),
            .I(N__34751));
    InMux I__6254 (
            .O(N__34782),
            .I(N__34744));
    InMux I__6253 (
            .O(N__34781),
            .I(N__34744));
    InMux I__6252 (
            .O(N__34778),
            .I(N__34744));
    InMux I__6251 (
            .O(N__34775),
            .I(N__34739));
    InMux I__6250 (
            .O(N__34774),
            .I(N__34739));
    LocalMux I__6249 (
            .O(N__34771),
            .I(N__34736));
    InMux I__6248 (
            .O(N__34768),
            .I(N__34733));
    LocalMux I__6247 (
            .O(N__34765),
            .I(N__34730));
    InMux I__6246 (
            .O(N__34762),
            .I(N__34723));
    InMux I__6245 (
            .O(N__34759),
            .I(N__34723));
    InMux I__6244 (
            .O(N__34756),
            .I(N__34723));
    LocalMux I__6243 (
            .O(N__34751),
            .I(N__34718));
    LocalMux I__6242 (
            .O(N__34744),
            .I(N__34718));
    LocalMux I__6241 (
            .O(N__34739),
            .I(eis_state_0));
    Odrv12 I__6240 (
            .O(N__34736),
            .I(eis_state_0));
    LocalMux I__6239 (
            .O(N__34733),
            .I(eis_state_0));
    Odrv12 I__6238 (
            .O(N__34730),
            .I(eis_state_0));
    LocalMux I__6237 (
            .O(N__34723),
            .I(eis_state_0));
    Odrv4 I__6236 (
            .O(N__34718),
            .I(eis_state_0));
    CascadeMux I__6235 (
            .O(N__34705),
            .I(N__34702));
    InMux I__6234 (
            .O(N__34702),
            .I(N__34692));
    InMux I__6233 (
            .O(N__34701),
            .I(N__34687));
    InMux I__6232 (
            .O(N__34700),
            .I(N__34687));
    CascadeMux I__6231 (
            .O(N__34699),
            .I(N__34682));
    CascadeMux I__6230 (
            .O(N__34698),
            .I(N__34679));
    InMux I__6229 (
            .O(N__34697),
            .I(N__34673));
    InMux I__6228 (
            .O(N__34696),
            .I(N__34673));
    CascadeMux I__6227 (
            .O(N__34695),
            .I(N__34667));
    LocalMux I__6226 (
            .O(N__34692),
            .I(N__34663));
    LocalMux I__6225 (
            .O(N__34687),
            .I(N__34660));
    InMux I__6224 (
            .O(N__34686),
            .I(N__34655));
    InMux I__6223 (
            .O(N__34685),
            .I(N__34655));
    InMux I__6222 (
            .O(N__34682),
            .I(N__34648));
    InMux I__6221 (
            .O(N__34679),
            .I(N__34648));
    InMux I__6220 (
            .O(N__34678),
            .I(N__34648));
    LocalMux I__6219 (
            .O(N__34673),
            .I(N__34645));
    InMux I__6218 (
            .O(N__34672),
            .I(N__34640));
    InMux I__6217 (
            .O(N__34671),
            .I(N__34640));
    InMux I__6216 (
            .O(N__34670),
            .I(N__34633));
    InMux I__6215 (
            .O(N__34667),
            .I(N__34633));
    InMux I__6214 (
            .O(N__34666),
            .I(N__34633));
    Odrv4 I__6213 (
            .O(N__34663),
            .I(eis_state_2));
    Odrv4 I__6212 (
            .O(N__34660),
            .I(eis_state_2));
    LocalMux I__6211 (
            .O(N__34655),
            .I(eis_state_2));
    LocalMux I__6210 (
            .O(N__34648),
            .I(eis_state_2));
    Odrv4 I__6209 (
            .O(N__34645),
            .I(eis_state_2));
    LocalMux I__6208 (
            .O(N__34640),
            .I(eis_state_2));
    LocalMux I__6207 (
            .O(N__34633),
            .I(eis_state_2));
    CascadeMux I__6206 (
            .O(N__34618),
            .I(n12450_cascade_));
    CascadeMux I__6205 (
            .O(N__34615),
            .I(N__34611));
    CascadeMux I__6204 (
            .O(N__34614),
            .I(N__34608));
    InMux I__6203 (
            .O(N__34611),
            .I(N__34605));
    InMux I__6202 (
            .O(N__34608),
            .I(N__34602));
    LocalMux I__6201 (
            .O(N__34605),
            .I(N__34599));
    LocalMux I__6200 (
            .O(N__34602),
            .I(N__34596));
    Span4Mux_h I__6199 (
            .O(N__34599),
            .I(N__34593));
    Span4Mux_h I__6198 (
            .O(N__34596),
            .I(N__34590));
    Span4Mux_v I__6197 (
            .O(N__34593),
            .I(N__34586));
    Span4Mux_v I__6196 (
            .O(N__34590),
            .I(N__34583));
    InMux I__6195 (
            .O(N__34589),
            .I(N__34580));
    Odrv4 I__6194 (
            .O(N__34586),
            .I(cmd_rdadctmp_16));
    Odrv4 I__6193 (
            .O(N__34583),
            .I(cmd_rdadctmp_16));
    LocalMux I__6192 (
            .O(N__34580),
            .I(cmd_rdadctmp_16));
    SRMux I__6191 (
            .O(N__34573),
            .I(N__34570));
    LocalMux I__6190 (
            .O(N__34570),
            .I(N__34567));
    Span4Mux_h I__6189 (
            .O(N__34567),
            .I(N__34564));
    Odrv4 I__6188 (
            .O(N__34564),
            .I(n22120));
    InMux I__6187 (
            .O(N__34561),
            .I(N__34558));
    LocalMux I__6186 (
            .O(N__34558),
            .I(n22312));
    InMux I__6185 (
            .O(N__34555),
            .I(N__34552));
    LocalMux I__6184 (
            .O(N__34552),
            .I(n23330));
    InMux I__6183 (
            .O(N__34549),
            .I(N__34543));
    InMux I__6182 (
            .O(N__34548),
            .I(N__34543));
    LocalMux I__6181 (
            .O(N__34543),
            .I(n17633));
    SRMux I__6180 (
            .O(N__34540),
            .I(N__34537));
    LocalMux I__6179 (
            .O(N__34537),
            .I(N__34531));
    SRMux I__6178 (
            .O(N__34536),
            .I(N__34528));
    SRMux I__6177 (
            .O(N__34535),
            .I(N__34525));
    SRMux I__6176 (
            .O(N__34534),
            .I(N__34519));
    Span4Mux_v I__6175 (
            .O(N__34531),
            .I(N__34511));
    LocalMux I__6174 (
            .O(N__34528),
            .I(N__34511));
    LocalMux I__6173 (
            .O(N__34525),
            .I(N__34511));
    SRMux I__6172 (
            .O(N__34524),
            .I(N__34508));
    SRMux I__6171 (
            .O(N__34523),
            .I(N__34505));
    SRMux I__6170 (
            .O(N__34522),
            .I(N__34500));
    LocalMux I__6169 (
            .O(N__34519),
            .I(N__34495));
    SRMux I__6168 (
            .O(N__34518),
            .I(N__34492));
    Span4Mux_v I__6167 (
            .O(N__34511),
            .I(N__34485));
    LocalMux I__6166 (
            .O(N__34508),
            .I(N__34485));
    LocalMux I__6165 (
            .O(N__34505),
            .I(N__34485));
    SRMux I__6164 (
            .O(N__34504),
            .I(N__34482));
    SRMux I__6163 (
            .O(N__34503),
            .I(N__34479));
    LocalMux I__6162 (
            .O(N__34500),
            .I(N__34476));
    SRMux I__6161 (
            .O(N__34499),
            .I(N__34473));
    SRMux I__6160 (
            .O(N__34498),
            .I(N__34470));
    Span4Mux_v I__6159 (
            .O(N__34495),
            .I(N__34465));
    LocalMux I__6158 (
            .O(N__34492),
            .I(N__34465));
    Span4Mux_v I__6157 (
            .O(N__34485),
            .I(N__34458));
    LocalMux I__6156 (
            .O(N__34482),
            .I(N__34458));
    LocalMux I__6155 (
            .O(N__34479),
            .I(N__34458));
    Span4Mux_v I__6154 (
            .O(N__34476),
            .I(N__34451));
    LocalMux I__6153 (
            .O(N__34473),
            .I(N__34451));
    LocalMux I__6152 (
            .O(N__34470),
            .I(N__34451));
    Span4Mux_v I__6151 (
            .O(N__34465),
            .I(N__34448));
    Span4Mux_v I__6150 (
            .O(N__34458),
            .I(N__34443));
    Span4Mux_v I__6149 (
            .O(N__34451),
            .I(N__34443));
    Span4Mux_v I__6148 (
            .O(N__34448),
            .I(N__34440));
    Span4Mux_h I__6147 (
            .O(N__34443),
            .I(N__34437));
    Span4Mux_h I__6146 (
            .O(N__34440),
            .I(N__34432));
    Span4Mux_h I__6145 (
            .O(N__34437),
            .I(N__34432));
    Odrv4 I__6144 (
            .O(N__34432),
            .I(iac_raw_buf_N_821));
    InMux I__6143 (
            .O(N__34429),
            .I(N__34426));
    LocalMux I__6142 (
            .O(N__34426),
            .I(n17_adj_1742));
    CEMux I__6141 (
            .O(N__34423),
            .I(N__34420));
    LocalMux I__6140 (
            .O(N__34420),
            .I(N__34416));
    CEMux I__6139 (
            .O(N__34419),
            .I(N__34413));
    Span4Mux_h I__6138 (
            .O(N__34416),
            .I(N__34410));
    LocalMux I__6137 (
            .O(N__34413),
            .I(N__34405));
    Span4Mux_h I__6136 (
            .O(N__34410),
            .I(N__34405));
    Odrv4 I__6135 (
            .O(N__34405),
            .I(n12369));
    CascadeMux I__6134 (
            .O(N__34402),
            .I(N__34399));
    InMux I__6133 (
            .O(N__34399),
            .I(N__34396));
    LocalMux I__6132 (
            .O(N__34396),
            .I(N__34393));
    Odrv4 I__6131 (
            .O(N__34393),
            .I(n24_adj_1503));
    InMux I__6130 (
            .O(N__34390),
            .I(N__34387));
    LocalMux I__6129 (
            .O(N__34387),
            .I(N__34382));
    InMux I__6128 (
            .O(N__34386),
            .I(N__34379));
    CascadeMux I__6127 (
            .O(N__34385),
            .I(N__34376));
    Span12Mux_v I__6126 (
            .O(N__34382),
            .I(N__34373));
    LocalMux I__6125 (
            .O(N__34379),
            .I(N__34370));
    InMux I__6124 (
            .O(N__34376),
            .I(N__34367));
    Span12Mux_h I__6123 (
            .O(N__34373),
            .I(N__34364));
    Span4Mux_h I__6122 (
            .O(N__34370),
            .I(N__34361));
    LocalMux I__6121 (
            .O(N__34367),
            .I(buf_adcdata_iac_16));
    Odrv12 I__6120 (
            .O(N__34364),
            .I(buf_adcdata_iac_16));
    Odrv4 I__6119 (
            .O(N__34361),
            .I(buf_adcdata_iac_16));
    InMux I__6118 (
            .O(N__34354),
            .I(N__34351));
    LocalMux I__6117 (
            .O(N__34351),
            .I(N__34348));
    Odrv4 I__6116 (
            .O(N__34348),
            .I(n23324));
    CascadeMux I__6115 (
            .O(N__34345),
            .I(N__34340));
    InMux I__6114 (
            .O(N__34344),
            .I(N__34335));
    InMux I__6113 (
            .O(N__34343),
            .I(N__34335));
    InMux I__6112 (
            .O(N__34340),
            .I(N__34332));
    LocalMux I__6111 (
            .O(N__34335),
            .I(req_data_cnt_8));
    LocalMux I__6110 (
            .O(N__34332),
            .I(req_data_cnt_8));
    CascadeMux I__6109 (
            .O(N__34327),
            .I(n19_adj_1727_cascade_));
    CascadeMux I__6108 (
            .O(N__34324),
            .I(n29_adj_1770_cascade_));
    InMux I__6107 (
            .O(N__34321),
            .I(N__34317));
    CascadeMux I__6106 (
            .O(N__34320),
            .I(N__34314));
    LocalMux I__6105 (
            .O(N__34317),
            .I(N__34311));
    InMux I__6104 (
            .O(N__34314),
            .I(N__34308));
    Span4Mux_v I__6103 (
            .O(N__34311),
            .I(N__34305));
    LocalMux I__6102 (
            .O(N__34308),
            .I(comm_test_buf_24_14));
    Odrv4 I__6101 (
            .O(N__34305),
            .I(comm_test_buf_24_14));
    InMux I__6100 (
            .O(N__34300),
            .I(N__34294));
    InMux I__6099 (
            .O(N__34299),
            .I(N__34294));
    LocalMux I__6098 (
            .O(N__34294),
            .I(N__34290));
    InMux I__6097 (
            .O(N__34293),
            .I(N__34287));
    Span4Mux_v I__6096 (
            .O(N__34290),
            .I(N__34284));
    LocalMux I__6095 (
            .O(N__34287),
            .I(N__34281));
    Odrv4 I__6094 (
            .O(N__34284),
            .I(comm_test_buf_24_6));
    Odrv12 I__6093 (
            .O(N__34281),
            .I(comm_test_buf_24_6));
    InMux I__6092 (
            .O(N__34276),
            .I(N__34271));
    InMux I__6091 (
            .O(N__34275),
            .I(N__34266));
    InMux I__6090 (
            .O(N__34274),
            .I(N__34266));
    LocalMux I__6089 (
            .O(N__34271),
            .I(n16_adj_1683));
    LocalMux I__6088 (
            .O(N__34266),
            .I(n16_adj_1683));
    CascadeMux I__6087 (
            .O(N__34261),
            .I(n17642_cascade_));
    InMux I__6086 (
            .O(N__34258),
            .I(N__34254));
    InMux I__6085 (
            .O(N__34257),
            .I(N__34251));
    LocalMux I__6084 (
            .O(N__34254),
            .I(comm_test_buf_24_11));
    LocalMux I__6083 (
            .O(N__34251),
            .I(comm_test_buf_24_11));
    InMux I__6082 (
            .O(N__34246),
            .I(N__34240));
    InMux I__6081 (
            .O(N__34245),
            .I(N__34240));
    LocalMux I__6080 (
            .O(N__34240),
            .I(comm_test_buf_24_12));
    InMux I__6079 (
            .O(N__34237),
            .I(N__34234));
    LocalMux I__6078 (
            .O(N__34234),
            .I(N__34231));
    Odrv4 I__6077 (
            .O(N__34231),
            .I(n13237));
    InMux I__6076 (
            .O(N__34228),
            .I(N__34225));
    LocalMux I__6075 (
            .O(N__34225),
            .I(N__34222));
    Span4Mux_v I__6074 (
            .O(N__34222),
            .I(N__34219));
    Odrv4 I__6073 (
            .O(N__34219),
            .I(n22295));
    CascadeMux I__6072 (
            .O(N__34216),
            .I(N__34213));
    InMux I__6071 (
            .O(N__34213),
            .I(N__34210));
    LocalMux I__6070 (
            .O(N__34210),
            .I(N__34207));
    Odrv4 I__6069 (
            .O(N__34207),
            .I(n4_adj_1667));
    InMux I__6068 (
            .O(N__34204),
            .I(N__34201));
    LocalMux I__6067 (
            .O(N__34201),
            .I(N__34198));
    Odrv4 I__6066 (
            .O(N__34198),
            .I(n23294));
    InMux I__6065 (
            .O(N__34195),
            .I(N__34192));
    LocalMux I__6064 (
            .O(N__34192),
            .I(N__34189));
    Odrv4 I__6063 (
            .O(N__34189),
            .I(n30_adj_1588));
    InMux I__6062 (
            .O(N__34186),
            .I(N__34183));
    LocalMux I__6061 (
            .O(N__34183),
            .I(N__34180));
    Span4Mux_v I__6060 (
            .O(N__34180),
            .I(N__34175));
    InMux I__6059 (
            .O(N__34179),
            .I(N__34172));
    InMux I__6058 (
            .O(N__34178),
            .I(N__34169));
    Odrv4 I__6057 (
            .O(N__34175),
            .I(comm_test_buf_24_3));
    LocalMux I__6056 (
            .O(N__34172),
            .I(comm_test_buf_24_3));
    LocalMux I__6055 (
            .O(N__34169),
            .I(comm_test_buf_24_3));
    InMux I__6054 (
            .O(N__34162),
            .I(N__34159));
    LocalMux I__6053 (
            .O(N__34159),
            .I(n111_adj_1794));
    SRMux I__6052 (
            .O(N__34156),
            .I(N__34153));
    LocalMux I__6051 (
            .O(N__34153),
            .I(n15545));
    InMux I__6050 (
            .O(N__34150),
            .I(N__34147));
    LocalMux I__6049 (
            .O(N__34147),
            .I(N__34144));
    Span4Mux_h I__6048 (
            .O(N__34144),
            .I(N__34140));
    CascadeMux I__6047 (
            .O(N__34143),
            .I(N__34137));
    Span4Mux_h I__6046 (
            .O(N__34140),
            .I(N__34133));
    InMux I__6045 (
            .O(N__34137),
            .I(N__34128));
    InMux I__6044 (
            .O(N__34136),
            .I(N__34128));
    Odrv4 I__6043 (
            .O(N__34133),
            .I(buf_dds1_8));
    LocalMux I__6042 (
            .O(N__34128),
            .I(buf_dds1_8));
    InMux I__6041 (
            .O(N__34123),
            .I(N__34120));
    LocalMux I__6040 (
            .O(N__34120),
            .I(N__34117));
    Odrv4 I__6039 (
            .O(N__34117),
            .I(n1_adj_1665));
    SRMux I__6038 (
            .O(N__34114),
            .I(N__34111));
    LocalMux I__6037 (
            .O(N__34111),
            .I(N__34108));
    Span4Mux_h I__6036 (
            .O(N__34108),
            .I(N__34105));
    Odrv4 I__6035 (
            .O(N__34105),
            .I(\comm_spi.data_tx_7__N_865 ));
    InMux I__6034 (
            .O(N__34102),
            .I(N__34099));
    LocalMux I__6033 (
            .O(N__34099),
            .I(N__34095));
    InMux I__6032 (
            .O(N__34098),
            .I(N__34092));
    Span4Mux_v I__6031 (
            .O(N__34095),
            .I(N__34088));
    LocalMux I__6030 (
            .O(N__34092),
            .I(N__34085));
    InMux I__6029 (
            .O(N__34091),
            .I(N__34082));
    Span4Mux_v I__6028 (
            .O(N__34088),
            .I(N__34077));
    Span4Mux_h I__6027 (
            .O(N__34085),
            .I(N__34077));
    LocalMux I__6026 (
            .O(N__34082),
            .I(comm_test_buf_24_4));
    Odrv4 I__6025 (
            .O(N__34077),
            .I(comm_test_buf_24_4));
    InMux I__6024 (
            .O(N__34072),
            .I(N__34069));
    LocalMux I__6023 (
            .O(N__34069),
            .I(n13231));
    CascadeMux I__6022 (
            .O(N__34066),
            .I(n19_adj_1710_cascade_));
    InMux I__6021 (
            .O(N__34063),
            .I(N__34060));
    LocalMux I__6020 (
            .O(N__34060),
            .I(N__34057));
    Span12Mux_h I__6019 (
            .O(N__34057),
            .I(N__34054));
    Odrv12 I__6018 (
            .O(N__34054),
            .I(buf_data_iac_1));
    CascadeMux I__6017 (
            .O(N__34051),
            .I(n22_adj_1711_cascade_));
    CascadeMux I__6016 (
            .O(N__34048),
            .I(n30_adj_1712_cascade_));
    InMux I__6015 (
            .O(N__34045),
            .I(N__34042));
    LocalMux I__6014 (
            .O(N__34042),
            .I(N__34039));
    Span4Mux_v I__6013 (
            .O(N__34039),
            .I(N__34036));
    Span4Mux_v I__6012 (
            .O(N__34036),
            .I(N__34032));
    InMux I__6011 (
            .O(N__34035),
            .I(N__34029));
    Span4Mux_h I__6010 (
            .O(N__34032),
            .I(N__34024));
    LocalMux I__6009 (
            .O(N__34029),
            .I(N__34024));
    Span4Mux_h I__6008 (
            .O(N__34024),
            .I(N__34020));
    InMux I__6007 (
            .O(N__34023),
            .I(N__34017));
    Odrv4 I__6006 (
            .O(N__34020),
            .I(\comm_spi.n24031 ));
    LocalMux I__6005 (
            .O(N__34017),
            .I(\comm_spi.n24031 ));
    InMux I__6004 (
            .O(N__34012),
            .I(N__34009));
    LocalMux I__6003 (
            .O(N__34009),
            .I(n30_adj_1705));
    CascadeMux I__6002 (
            .O(N__34006),
            .I(N__34003));
    InMux I__6001 (
            .O(N__34003),
            .I(N__33997));
    InMux I__6000 (
            .O(N__34002),
            .I(N__33994));
    InMux I__5999 (
            .O(N__34001),
            .I(N__33982));
    CascadeMux I__5998 (
            .O(N__34000),
            .I(N__33975));
    LocalMux I__5997 (
            .O(N__33997),
            .I(N__33967));
    LocalMux I__5996 (
            .O(N__33994),
            .I(N__33967));
    InMux I__5995 (
            .O(N__33993),
            .I(N__33962));
    InMux I__5994 (
            .O(N__33992),
            .I(N__33962));
    InMux I__5993 (
            .O(N__33991),
            .I(N__33955));
    InMux I__5992 (
            .O(N__33990),
            .I(N__33955));
    InMux I__5991 (
            .O(N__33989),
            .I(N__33955));
    InMux I__5990 (
            .O(N__33988),
            .I(N__33945));
    InMux I__5989 (
            .O(N__33987),
            .I(N__33945));
    InMux I__5988 (
            .O(N__33986),
            .I(N__33940));
    InMux I__5987 (
            .O(N__33985),
            .I(N__33940));
    LocalMux I__5986 (
            .O(N__33982),
            .I(N__33931));
    InMux I__5985 (
            .O(N__33981),
            .I(N__33928));
    InMux I__5984 (
            .O(N__33980),
            .I(N__33921));
    InMux I__5983 (
            .O(N__33979),
            .I(N__33921));
    InMux I__5982 (
            .O(N__33978),
            .I(N__33921));
    InMux I__5981 (
            .O(N__33975),
            .I(N__33914));
    InMux I__5980 (
            .O(N__33974),
            .I(N__33914));
    InMux I__5979 (
            .O(N__33973),
            .I(N__33914));
    InMux I__5978 (
            .O(N__33972),
            .I(N__33911));
    Span4Mux_v I__5977 (
            .O(N__33967),
            .I(N__33908));
    LocalMux I__5976 (
            .O(N__33962),
            .I(N__33903));
    LocalMux I__5975 (
            .O(N__33955),
            .I(N__33903));
    InMux I__5974 (
            .O(N__33954),
            .I(N__33897));
    InMux I__5973 (
            .O(N__33953),
            .I(N__33897));
    InMux I__5972 (
            .O(N__33952),
            .I(N__33892));
    InMux I__5971 (
            .O(N__33951),
            .I(N__33892));
    InMux I__5970 (
            .O(N__33950),
            .I(N__33889));
    LocalMux I__5969 (
            .O(N__33945),
            .I(N__33886));
    LocalMux I__5968 (
            .O(N__33940),
            .I(N__33883));
    InMux I__5967 (
            .O(N__33939),
            .I(N__33880));
    InMux I__5966 (
            .O(N__33938),
            .I(N__33877));
    InMux I__5965 (
            .O(N__33937),
            .I(N__33868));
    InMux I__5964 (
            .O(N__33936),
            .I(N__33868));
    InMux I__5963 (
            .O(N__33935),
            .I(N__33868));
    InMux I__5962 (
            .O(N__33934),
            .I(N__33868));
    Span4Mux_h I__5961 (
            .O(N__33931),
            .I(N__33861));
    LocalMux I__5960 (
            .O(N__33928),
            .I(N__33861));
    LocalMux I__5959 (
            .O(N__33921),
            .I(N__33861));
    LocalMux I__5958 (
            .O(N__33914),
            .I(N__33858));
    LocalMux I__5957 (
            .O(N__33911),
            .I(N__33851));
    Span4Mux_h I__5956 (
            .O(N__33908),
            .I(N__33851));
    Span4Mux_v I__5955 (
            .O(N__33903),
            .I(N__33851));
    InMux I__5954 (
            .O(N__33902),
            .I(N__33848));
    LocalMux I__5953 (
            .O(N__33897),
            .I(N__33845));
    LocalMux I__5952 (
            .O(N__33892),
            .I(N__33836));
    LocalMux I__5951 (
            .O(N__33889),
            .I(N__33836));
    Span4Mux_h I__5950 (
            .O(N__33886),
            .I(N__33836));
    Span4Mux_v I__5949 (
            .O(N__33883),
            .I(N__33836));
    LocalMux I__5948 (
            .O(N__33880),
            .I(N__33823));
    LocalMux I__5947 (
            .O(N__33877),
            .I(N__33823));
    LocalMux I__5946 (
            .O(N__33868),
            .I(N__33823));
    Span4Mux_v I__5945 (
            .O(N__33861),
            .I(N__33823));
    Span4Mux_v I__5944 (
            .O(N__33858),
            .I(N__33823));
    Span4Mux_h I__5943 (
            .O(N__33851),
            .I(N__33823));
    LocalMux I__5942 (
            .O(N__33848),
            .I(N__33820));
    Span4Mux_v I__5941 (
            .O(N__33845),
            .I(N__33815));
    Span4Mux_v I__5940 (
            .O(N__33836),
            .I(N__33815));
    Span4Mux_h I__5939 (
            .O(N__33823),
            .I(N__33812));
    Odrv12 I__5938 (
            .O(N__33820),
            .I(n13847));
    Odrv4 I__5937 (
            .O(N__33815),
            .I(n13847));
    Odrv4 I__5936 (
            .O(N__33812),
            .I(n13847));
    CascadeMux I__5935 (
            .O(N__33805),
            .I(N__33801));
    CascadeMux I__5934 (
            .O(N__33804),
            .I(N__33798));
    InMux I__5933 (
            .O(N__33801),
            .I(N__33794));
    InMux I__5932 (
            .O(N__33798),
            .I(N__33789));
    InMux I__5931 (
            .O(N__33797),
            .I(N__33789));
    LocalMux I__5930 (
            .O(N__33794),
            .I(cmd_rdadctmp_9_adj_1539));
    LocalMux I__5929 (
            .O(N__33789),
            .I(cmd_rdadctmp_9_adj_1539));
    CascadeMux I__5928 (
            .O(N__33784),
            .I(n2_adj_1666_cascade_));
    SRMux I__5927 (
            .O(N__33781),
            .I(N__33778));
    LocalMux I__5926 (
            .O(N__33778),
            .I(N__33775));
    Odrv12 I__5925 (
            .O(N__33775),
            .I(\ADC_VDC.n17542 ));
    InMux I__5924 (
            .O(N__33772),
            .I(N__33768));
    InMux I__5923 (
            .O(N__33771),
            .I(N__33765));
    LocalMux I__5922 (
            .O(N__33768),
            .I(N__33762));
    LocalMux I__5921 (
            .O(N__33765),
            .I(N__33759));
    Span4Mux_v I__5920 (
            .O(N__33762),
            .I(N__33756));
    Span4Mux_h I__5919 (
            .O(N__33759),
            .I(N__33753));
    Odrv4 I__5918 (
            .O(N__33756),
            .I(\comm_spi.n15361 ));
    Odrv4 I__5917 (
            .O(N__33753),
            .I(\comm_spi.n15361 ));
    InMux I__5916 (
            .O(N__33748),
            .I(N__33745));
    LocalMux I__5915 (
            .O(N__33745),
            .I(N__33742));
    Span4Mux_v I__5914 (
            .O(N__33742),
            .I(N__33738));
    CascadeMux I__5913 (
            .O(N__33741),
            .I(N__33735));
    Span4Mux_h I__5912 (
            .O(N__33738),
            .I(N__33732));
    InMux I__5911 (
            .O(N__33735),
            .I(N__33729));
    Odrv4 I__5910 (
            .O(N__33732),
            .I(buf_adcdata_vdc_3));
    LocalMux I__5909 (
            .O(N__33729),
            .I(buf_adcdata_vdc_3));
    CascadeMux I__5908 (
            .O(N__33724),
            .I(n19_adj_1703_cascade_));
    InMux I__5907 (
            .O(N__33721),
            .I(N__33718));
    LocalMux I__5906 (
            .O(N__33718),
            .I(N__33715));
    Span4Mux_h I__5905 (
            .O(N__33715),
            .I(N__33712));
    Span4Mux_h I__5904 (
            .O(N__33712),
            .I(N__33709));
    Span4Mux_h I__5903 (
            .O(N__33709),
            .I(N__33706));
    Odrv4 I__5902 (
            .O(N__33706),
            .I(buf_data_iac_3));
    CascadeMux I__5901 (
            .O(N__33703),
            .I(n22_adj_1704_cascade_));
    InMux I__5900 (
            .O(N__33700),
            .I(N__33697));
    LocalMux I__5899 (
            .O(N__33697),
            .I(N__33694));
    Span4Mux_v I__5898 (
            .O(N__33694),
            .I(N__33691));
    Sp12to4 I__5897 (
            .O(N__33691),
            .I(N__33686));
    InMux I__5896 (
            .O(N__33690),
            .I(N__33681));
    InMux I__5895 (
            .O(N__33689),
            .I(N__33681));
    Odrv12 I__5894 (
            .O(N__33686),
            .I(buf_adcdata_iac_3));
    LocalMux I__5893 (
            .O(N__33681),
            .I(buf_adcdata_iac_3));
    InMux I__5892 (
            .O(N__33676),
            .I(N__33673));
    LocalMux I__5891 (
            .O(N__33673),
            .I(N__33670));
    Span12Mux_v I__5890 (
            .O(N__33670),
            .I(N__33665));
    InMux I__5889 (
            .O(N__33669),
            .I(N__33660));
    InMux I__5888 (
            .O(N__33668),
            .I(N__33660));
    Odrv12 I__5887 (
            .O(N__33665),
            .I(cmd_rdadctmp_11_adj_1537));
    LocalMux I__5886 (
            .O(N__33660),
            .I(cmd_rdadctmp_11_adj_1537));
    InMux I__5885 (
            .O(N__33655),
            .I(N__33652));
    LocalMux I__5884 (
            .O(N__33652),
            .I(N__33649));
    Span4Mux_v I__5883 (
            .O(N__33649),
            .I(N__33646));
    Sp12to4 I__5882 (
            .O(N__33646),
            .I(N__33641));
    InMux I__5881 (
            .O(N__33645),
            .I(N__33636));
    InMux I__5880 (
            .O(N__33644),
            .I(N__33636));
    Odrv12 I__5879 (
            .O(N__33641),
            .I(buf_adcdata_vac_3));
    LocalMux I__5878 (
            .O(N__33636),
            .I(buf_adcdata_vac_3));
    InMux I__5877 (
            .O(N__33631),
            .I(N__33628));
    LocalMux I__5876 (
            .O(N__33628),
            .I(N__33624));
    CascadeMux I__5875 (
            .O(N__33627),
            .I(N__33621));
    Span4Mux_h I__5874 (
            .O(N__33624),
            .I(N__33618));
    InMux I__5873 (
            .O(N__33621),
            .I(N__33615));
    Odrv4 I__5872 (
            .O(N__33618),
            .I(buf_adcdata_vdc_1));
    LocalMux I__5871 (
            .O(N__33615),
            .I(buf_adcdata_vdc_1));
    InMux I__5870 (
            .O(N__33610),
            .I(N__33607));
    LocalMux I__5869 (
            .O(N__33607),
            .I(N__33603));
    InMux I__5868 (
            .O(N__33606),
            .I(N__33599));
    Span12Mux_h I__5867 (
            .O(N__33603),
            .I(N__33596));
    InMux I__5866 (
            .O(N__33602),
            .I(N__33593));
    LocalMux I__5865 (
            .O(N__33599),
            .I(buf_adcdata_vac_1));
    Odrv12 I__5864 (
            .O(N__33596),
            .I(buf_adcdata_vac_1));
    LocalMux I__5863 (
            .O(N__33593),
            .I(buf_adcdata_vac_1));
    InMux I__5862 (
            .O(N__33586),
            .I(N__33583));
    LocalMux I__5861 (
            .O(N__33583),
            .I(N__33570));
    InMux I__5860 (
            .O(N__33582),
            .I(N__33567));
    InMux I__5859 (
            .O(N__33581),
            .I(N__33564));
    InMux I__5858 (
            .O(N__33580),
            .I(N__33561));
    InMux I__5857 (
            .O(N__33579),
            .I(N__33556));
    InMux I__5856 (
            .O(N__33578),
            .I(N__33556));
    InMux I__5855 (
            .O(N__33577),
            .I(N__33553));
    InMux I__5854 (
            .O(N__33576),
            .I(N__33545));
    InMux I__5853 (
            .O(N__33575),
            .I(N__33542));
    InMux I__5852 (
            .O(N__33574),
            .I(N__33537));
    InMux I__5851 (
            .O(N__33573),
            .I(N__33537));
    Span4Mux_v I__5850 (
            .O(N__33570),
            .I(N__33526));
    LocalMux I__5849 (
            .O(N__33567),
            .I(N__33526));
    LocalMux I__5848 (
            .O(N__33564),
            .I(N__33517));
    LocalMux I__5847 (
            .O(N__33561),
            .I(N__33517));
    LocalMux I__5846 (
            .O(N__33556),
            .I(N__33517));
    LocalMux I__5845 (
            .O(N__33553),
            .I(N__33517));
    InMux I__5844 (
            .O(N__33552),
            .I(N__33513));
    InMux I__5843 (
            .O(N__33551),
            .I(N__33510));
    InMux I__5842 (
            .O(N__33550),
            .I(N__33507));
    InMux I__5841 (
            .O(N__33549),
            .I(N__33504));
    InMux I__5840 (
            .O(N__33548),
            .I(N__33501));
    LocalMux I__5839 (
            .O(N__33545),
            .I(N__33494));
    LocalMux I__5838 (
            .O(N__33542),
            .I(N__33494));
    LocalMux I__5837 (
            .O(N__33537),
            .I(N__33494));
    InMux I__5836 (
            .O(N__33536),
            .I(N__33485));
    InMux I__5835 (
            .O(N__33535),
            .I(N__33485));
    InMux I__5834 (
            .O(N__33534),
            .I(N__33485));
    InMux I__5833 (
            .O(N__33533),
            .I(N__33485));
    InMux I__5832 (
            .O(N__33532),
            .I(N__33480));
    InMux I__5831 (
            .O(N__33531),
            .I(N__33480));
    Span4Mux_v I__5830 (
            .O(N__33526),
            .I(N__33475));
    Span4Mux_v I__5829 (
            .O(N__33517),
            .I(N__33475));
    InMux I__5828 (
            .O(N__33516),
            .I(N__33472));
    LocalMux I__5827 (
            .O(N__33513),
            .I(N__33467));
    LocalMux I__5826 (
            .O(N__33510),
            .I(N__33467));
    LocalMux I__5825 (
            .O(N__33507),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__5824 (
            .O(N__33504),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__5823 (
            .O(N__33501),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv12 I__5822 (
            .O(N__33494),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__5821 (
            .O(N__33485),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__5820 (
            .O(N__33480),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__5819 (
            .O(N__33475),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__5818 (
            .O(N__33472),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__5817 (
            .O(N__33467),
            .I(\ADC_VDC.adc_state_0 ));
    CascadeMux I__5816 (
            .O(N__33448),
            .I(N__33433));
    InMux I__5815 (
            .O(N__33447),
            .I(N__33426));
    InMux I__5814 (
            .O(N__33446),
            .I(N__33411));
    InMux I__5813 (
            .O(N__33445),
            .I(N__33411));
    InMux I__5812 (
            .O(N__33444),
            .I(N__33411));
    InMux I__5811 (
            .O(N__33443),
            .I(N__33411));
    InMux I__5810 (
            .O(N__33442),
            .I(N__33411));
    InMux I__5809 (
            .O(N__33441),
            .I(N__33411));
    InMux I__5808 (
            .O(N__33440),
            .I(N__33411));
    CascadeMux I__5807 (
            .O(N__33439),
            .I(N__33407));
    CascadeMux I__5806 (
            .O(N__33438),
            .I(N__33404));
    CascadeMux I__5805 (
            .O(N__33437),
            .I(N__33399));
    InMux I__5804 (
            .O(N__33436),
            .I(N__33388));
    InMux I__5803 (
            .O(N__33433),
            .I(N__33388));
    CascadeMux I__5802 (
            .O(N__33432),
            .I(N__33382));
    CascadeMux I__5801 (
            .O(N__33431),
            .I(N__33375));
    CascadeMux I__5800 (
            .O(N__33430),
            .I(N__33372));
    CascadeMux I__5799 (
            .O(N__33429),
            .I(N__33369));
    LocalMux I__5798 (
            .O(N__33426),
            .I(N__33363));
    LocalMux I__5797 (
            .O(N__33411),
            .I(N__33363));
    InMux I__5796 (
            .O(N__33410),
            .I(N__33356));
    InMux I__5795 (
            .O(N__33407),
            .I(N__33356));
    InMux I__5794 (
            .O(N__33404),
            .I(N__33356));
    CascadeMux I__5793 (
            .O(N__33403),
            .I(N__33349));
    InMux I__5792 (
            .O(N__33402),
            .I(N__33333));
    InMux I__5791 (
            .O(N__33399),
            .I(N__33333));
    InMux I__5790 (
            .O(N__33398),
            .I(N__33333));
    InMux I__5789 (
            .O(N__33397),
            .I(N__33333));
    InMux I__5788 (
            .O(N__33396),
            .I(N__33333));
    InMux I__5787 (
            .O(N__33395),
            .I(N__33333));
    InMux I__5786 (
            .O(N__33394),
            .I(N__33333));
    InMux I__5785 (
            .O(N__33393),
            .I(N__33330));
    LocalMux I__5784 (
            .O(N__33388),
            .I(N__33327));
    InMux I__5783 (
            .O(N__33387),
            .I(N__33320));
    InMux I__5782 (
            .O(N__33386),
            .I(N__33320));
    InMux I__5781 (
            .O(N__33385),
            .I(N__33320));
    InMux I__5780 (
            .O(N__33382),
            .I(N__33315));
    CascadeMux I__5779 (
            .O(N__33381),
            .I(N__33311));
    InMux I__5778 (
            .O(N__33380),
            .I(N__33308));
    InMux I__5777 (
            .O(N__33379),
            .I(N__33303));
    InMux I__5776 (
            .O(N__33378),
            .I(N__33303));
    InMux I__5775 (
            .O(N__33375),
            .I(N__33300));
    InMux I__5774 (
            .O(N__33372),
            .I(N__33295));
    InMux I__5773 (
            .O(N__33369),
            .I(N__33295));
    CascadeMux I__5772 (
            .O(N__33368),
            .I(N__33292));
    Span4Mux_h I__5771 (
            .O(N__33363),
            .I(N__33285));
    LocalMux I__5770 (
            .O(N__33356),
            .I(N__33285));
    InMux I__5769 (
            .O(N__33355),
            .I(N__33274));
    InMux I__5768 (
            .O(N__33354),
            .I(N__33274));
    InMux I__5767 (
            .O(N__33353),
            .I(N__33274));
    InMux I__5766 (
            .O(N__33352),
            .I(N__33274));
    InMux I__5765 (
            .O(N__33349),
            .I(N__33274));
    CascadeMux I__5764 (
            .O(N__33348),
            .I(N__33270));
    LocalMux I__5763 (
            .O(N__33333),
            .I(N__33267));
    LocalMux I__5762 (
            .O(N__33330),
            .I(N__33261));
    Span4Mux_h I__5761 (
            .O(N__33327),
            .I(N__33261));
    LocalMux I__5760 (
            .O(N__33320),
            .I(N__33258));
    InMux I__5759 (
            .O(N__33319),
            .I(N__33253));
    InMux I__5758 (
            .O(N__33318),
            .I(N__33253));
    LocalMux I__5757 (
            .O(N__33315),
            .I(N__33250));
    InMux I__5756 (
            .O(N__33314),
            .I(N__33246));
    InMux I__5755 (
            .O(N__33311),
            .I(N__33243));
    LocalMux I__5754 (
            .O(N__33308),
            .I(N__33240));
    LocalMux I__5753 (
            .O(N__33303),
            .I(N__33233));
    LocalMux I__5752 (
            .O(N__33300),
            .I(N__33233));
    LocalMux I__5751 (
            .O(N__33295),
            .I(N__33233));
    InMux I__5750 (
            .O(N__33292),
            .I(N__33226));
    InMux I__5749 (
            .O(N__33291),
            .I(N__33226));
    InMux I__5748 (
            .O(N__33290),
            .I(N__33226));
    Span4Mux_v I__5747 (
            .O(N__33285),
            .I(N__33221));
    LocalMux I__5746 (
            .O(N__33274),
            .I(N__33221));
    InMux I__5745 (
            .O(N__33273),
            .I(N__33218));
    InMux I__5744 (
            .O(N__33270),
            .I(N__33215));
    Span12Mux_v I__5743 (
            .O(N__33267),
            .I(N__33212));
    InMux I__5742 (
            .O(N__33266),
            .I(N__33209));
    Span4Mux_v I__5741 (
            .O(N__33261),
            .I(N__33206));
    Span4Mux_v I__5740 (
            .O(N__33258),
            .I(N__33201));
    LocalMux I__5739 (
            .O(N__33253),
            .I(N__33201));
    Span4Mux_h I__5738 (
            .O(N__33250),
            .I(N__33198));
    InMux I__5737 (
            .O(N__33249),
            .I(N__33195));
    LocalMux I__5736 (
            .O(N__33246),
            .I(N__33182));
    LocalMux I__5735 (
            .O(N__33243),
            .I(N__33182));
    Span4Mux_h I__5734 (
            .O(N__33240),
            .I(N__33182));
    Span4Mux_h I__5733 (
            .O(N__33233),
            .I(N__33182));
    LocalMux I__5732 (
            .O(N__33226),
            .I(N__33182));
    Span4Mux_v I__5731 (
            .O(N__33221),
            .I(N__33182));
    LocalMux I__5730 (
            .O(N__33218),
            .I(adc_state_2_adj_1550));
    LocalMux I__5729 (
            .O(N__33215),
            .I(adc_state_2_adj_1550));
    Odrv12 I__5728 (
            .O(N__33212),
            .I(adc_state_2_adj_1550));
    LocalMux I__5727 (
            .O(N__33209),
            .I(adc_state_2_adj_1550));
    Odrv4 I__5726 (
            .O(N__33206),
            .I(adc_state_2_adj_1550));
    Odrv4 I__5725 (
            .O(N__33201),
            .I(adc_state_2_adj_1550));
    Odrv4 I__5724 (
            .O(N__33198),
            .I(adc_state_2_adj_1550));
    LocalMux I__5723 (
            .O(N__33195),
            .I(adc_state_2_adj_1550));
    Odrv4 I__5722 (
            .O(N__33182),
            .I(adc_state_2_adj_1550));
    InMux I__5721 (
            .O(N__33163),
            .I(N__33160));
    LocalMux I__5720 (
            .O(N__33160),
            .I(\ADC_VDC.n11183 ));
    InMux I__5719 (
            .O(N__33157),
            .I(N__33154));
    LocalMux I__5718 (
            .O(N__33154),
            .I(\ADC_VDC.n23528 ));
    InMux I__5717 (
            .O(N__33151),
            .I(N__33147));
    InMux I__5716 (
            .O(N__33150),
            .I(N__33141));
    LocalMux I__5715 (
            .O(N__33147),
            .I(N__33138));
    InMux I__5714 (
            .O(N__33146),
            .I(N__33135));
    InMux I__5713 (
            .O(N__33145),
            .I(N__33130));
    InMux I__5712 (
            .O(N__33144),
            .I(N__33130));
    LocalMux I__5711 (
            .O(N__33141),
            .I(\ADC_VDC.bit_cnt_0 ));
    Odrv4 I__5710 (
            .O(N__33138),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__5709 (
            .O(N__33135),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__5708 (
            .O(N__33130),
            .I(\ADC_VDC.bit_cnt_0 ));
    InMux I__5707 (
            .O(N__33121),
            .I(bfn_11_6_0_));
    InMux I__5706 (
            .O(N__33118),
            .I(N__33112));
    InMux I__5705 (
            .O(N__33117),
            .I(N__33109));
    InMux I__5704 (
            .O(N__33116),
            .I(N__33106));
    InMux I__5703 (
            .O(N__33115),
            .I(N__33103));
    LocalMux I__5702 (
            .O(N__33112),
            .I(N__33096));
    LocalMux I__5701 (
            .O(N__33109),
            .I(N__33096));
    LocalMux I__5700 (
            .O(N__33106),
            .I(N__33096));
    LocalMux I__5699 (
            .O(N__33103),
            .I(\ADC_VDC.bit_cnt_1 ));
    Odrv4 I__5698 (
            .O(N__33096),
            .I(\ADC_VDC.bit_cnt_1 ));
    InMux I__5697 (
            .O(N__33091),
            .I(\ADC_VDC.n20812 ));
    CascadeMux I__5696 (
            .O(N__33088),
            .I(N__33083));
    CascadeMux I__5695 (
            .O(N__33087),
            .I(N__33080));
    InMux I__5694 (
            .O(N__33086),
            .I(N__33077));
    InMux I__5693 (
            .O(N__33083),
            .I(N__33073));
    InMux I__5692 (
            .O(N__33080),
            .I(N__33070));
    LocalMux I__5691 (
            .O(N__33077),
            .I(N__33067));
    InMux I__5690 (
            .O(N__33076),
            .I(N__33063));
    LocalMux I__5689 (
            .O(N__33073),
            .I(N__33056));
    LocalMux I__5688 (
            .O(N__33070),
            .I(N__33056));
    Span4Mux_v I__5687 (
            .O(N__33067),
            .I(N__33056));
    InMux I__5686 (
            .O(N__33066),
            .I(N__33053));
    LocalMux I__5685 (
            .O(N__33063),
            .I(\ADC_VDC.bit_cnt_2 ));
    Odrv4 I__5684 (
            .O(N__33056),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__5683 (
            .O(N__33053),
            .I(\ADC_VDC.bit_cnt_2 ));
    InMux I__5682 (
            .O(N__33046),
            .I(\ADC_VDC.n20813 ));
    InMux I__5681 (
            .O(N__33043),
            .I(N__33036));
    InMux I__5680 (
            .O(N__33042),
            .I(N__33033));
    InMux I__5679 (
            .O(N__33041),
            .I(N__33028));
    InMux I__5678 (
            .O(N__33040),
            .I(N__33028));
    InMux I__5677 (
            .O(N__33039),
            .I(N__33025));
    LocalMux I__5676 (
            .O(N__33036),
            .I(N__33022));
    LocalMux I__5675 (
            .O(N__33033),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__5674 (
            .O(N__33028),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__5673 (
            .O(N__33025),
            .I(\ADC_VDC.bit_cnt_3 ));
    Odrv4 I__5672 (
            .O(N__33022),
            .I(\ADC_VDC.bit_cnt_3 ));
    InMux I__5671 (
            .O(N__33013),
            .I(\ADC_VDC.n20814 ));
    InMux I__5670 (
            .O(N__33010),
            .I(N__33003));
    InMux I__5669 (
            .O(N__33009),
            .I(N__33000));
    InMux I__5668 (
            .O(N__33008),
            .I(N__32997));
    InMux I__5667 (
            .O(N__33007),
            .I(N__32992));
    InMux I__5666 (
            .O(N__33006),
            .I(N__32992));
    LocalMux I__5665 (
            .O(N__33003),
            .I(N__32989));
    LocalMux I__5664 (
            .O(N__33000),
            .I(\ADC_VDC.bit_cnt_4 ));
    LocalMux I__5663 (
            .O(N__32997),
            .I(\ADC_VDC.bit_cnt_4 ));
    LocalMux I__5662 (
            .O(N__32992),
            .I(\ADC_VDC.bit_cnt_4 ));
    Odrv4 I__5661 (
            .O(N__32989),
            .I(\ADC_VDC.bit_cnt_4 ));
    InMux I__5660 (
            .O(N__32980),
            .I(\ADC_VDC.n20815 ));
    InMux I__5659 (
            .O(N__32977),
            .I(N__32973));
    InMux I__5658 (
            .O(N__32976),
            .I(N__32970));
    LocalMux I__5657 (
            .O(N__32973),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__5656 (
            .O(N__32970),
            .I(\ADC_VDC.bit_cnt_5 ));
    InMux I__5655 (
            .O(N__32965),
            .I(\ADC_VDC.n20816 ));
    InMux I__5654 (
            .O(N__32962),
            .I(N__32958));
    InMux I__5653 (
            .O(N__32961),
            .I(N__32955));
    LocalMux I__5652 (
            .O(N__32958),
            .I(\ADC_VDC.bit_cnt_6 ));
    LocalMux I__5651 (
            .O(N__32955),
            .I(\ADC_VDC.bit_cnt_6 ));
    InMux I__5650 (
            .O(N__32950),
            .I(\ADC_VDC.n20817 ));
    InMux I__5649 (
            .O(N__32947),
            .I(\ADC_VDC.n20818 ));
    InMux I__5648 (
            .O(N__32944),
            .I(N__32940));
    InMux I__5647 (
            .O(N__32943),
            .I(N__32937));
    LocalMux I__5646 (
            .O(N__32940),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__5645 (
            .O(N__32937),
            .I(\ADC_VDC.bit_cnt_7 ));
    CEMux I__5644 (
            .O(N__32932),
            .I(N__32929));
    LocalMux I__5643 (
            .O(N__32929),
            .I(N__32926));
    Odrv12 I__5642 (
            .O(N__32926),
            .I(\ADC_VDC.n17565 ));
    CascadeMux I__5641 (
            .O(N__32923),
            .I(N__32920));
    InMux I__5640 (
            .O(N__32920),
            .I(N__32917));
    LocalMux I__5639 (
            .O(N__32917),
            .I(N__32914));
    Odrv4 I__5638 (
            .O(N__32914),
            .I(\SIG_DDS.tmp_buf_10 ));
    InMux I__5637 (
            .O(N__32911),
            .I(N__32908));
    LocalMux I__5636 (
            .O(N__32908),
            .I(N__32905));
    Span12Mux_v I__5635 (
            .O(N__32905),
            .I(N__32900));
    InMux I__5634 (
            .O(N__32904),
            .I(N__32897));
    InMux I__5633 (
            .O(N__32903),
            .I(N__32894));
    Odrv12 I__5632 (
            .O(N__32900),
            .I(buf_dds0_11));
    LocalMux I__5631 (
            .O(N__32897),
            .I(buf_dds0_11));
    LocalMux I__5630 (
            .O(N__32894),
            .I(buf_dds0_11));
    InMux I__5629 (
            .O(N__32887),
            .I(N__32884));
    LocalMux I__5628 (
            .O(N__32884),
            .I(\SIG_DDS.tmp_buf_11 ));
    InMux I__5627 (
            .O(N__32881),
            .I(N__32878));
    LocalMux I__5626 (
            .O(N__32878),
            .I(\ADC_VDC.n22063 ));
    InMux I__5625 (
            .O(N__32875),
            .I(N__32869));
    InMux I__5624 (
            .O(N__32874),
            .I(N__32862));
    InMux I__5623 (
            .O(N__32873),
            .I(N__32862));
    InMux I__5622 (
            .O(N__32872),
            .I(N__32862));
    LocalMux I__5621 (
            .O(N__32869),
            .I(N__32857));
    LocalMux I__5620 (
            .O(N__32862),
            .I(N__32857));
    Odrv12 I__5619 (
            .O(N__32857),
            .I(\RTD.n20050 ));
    InMux I__5618 (
            .O(N__32854),
            .I(N__32845));
    InMux I__5617 (
            .O(N__32853),
            .I(N__32840));
    InMux I__5616 (
            .O(N__32852),
            .I(N__32840));
    InMux I__5615 (
            .O(N__32851),
            .I(N__32837));
    InMux I__5614 (
            .O(N__32850),
            .I(N__32834));
    InMux I__5613 (
            .O(N__32849),
            .I(N__32830));
    CascadeMux I__5612 (
            .O(N__32848),
            .I(N__32825));
    LocalMux I__5611 (
            .O(N__32845),
            .I(N__32820));
    LocalMux I__5610 (
            .O(N__32840),
            .I(N__32820));
    LocalMux I__5609 (
            .O(N__32837),
            .I(N__32815));
    LocalMux I__5608 (
            .O(N__32834),
            .I(N__32815));
    InMux I__5607 (
            .O(N__32833),
            .I(N__32812));
    LocalMux I__5606 (
            .O(N__32830),
            .I(N__32809));
    InMux I__5605 (
            .O(N__32829),
            .I(N__32804));
    InMux I__5604 (
            .O(N__32828),
            .I(N__32804));
    InMux I__5603 (
            .O(N__32825),
            .I(N__32801));
    Span4Mux_v I__5602 (
            .O(N__32820),
            .I(N__32795));
    Span4Mux_v I__5601 (
            .O(N__32815),
            .I(N__32795));
    LocalMux I__5600 (
            .O(N__32812),
            .I(N__32792));
    Span4Mux_h I__5599 (
            .O(N__32809),
            .I(N__32785));
    LocalMux I__5598 (
            .O(N__32804),
            .I(N__32785));
    LocalMux I__5597 (
            .O(N__32801),
            .I(N__32785));
    CascadeMux I__5596 (
            .O(N__32800),
            .I(N__32782));
    Span4Mux_v I__5595 (
            .O(N__32795),
            .I(N__32779));
    Span4Mux_v I__5594 (
            .O(N__32792),
            .I(N__32774));
    Span4Mux_v I__5593 (
            .O(N__32785),
            .I(N__32774));
    InMux I__5592 (
            .O(N__32782),
            .I(N__32771));
    Sp12to4 I__5591 (
            .O(N__32779),
            .I(N__32768));
    Span4Mux_v I__5590 (
            .O(N__32774),
            .I(N__32765));
    LocalMux I__5589 (
            .O(N__32771),
            .I(N__32762));
    Span12Mux_h I__5588 (
            .O(N__32768),
            .I(N__32755));
    Sp12to4 I__5587 (
            .O(N__32765),
            .I(N__32755));
    Span12Mux_v I__5586 (
            .O(N__32762),
            .I(N__32755));
    Odrv12 I__5585 (
            .O(N__32755),
            .I(VDC_SDO));
    CascadeMux I__5584 (
            .O(N__32752),
            .I(\ADC_VDC.n35_cascade_ ));
    InMux I__5583 (
            .O(N__32749),
            .I(N__32746));
    LocalMux I__5582 (
            .O(N__32746),
            .I(\ADC_VDC.n45 ));
    CascadeMux I__5581 (
            .O(N__32743),
            .I(N__32740));
    InMux I__5580 (
            .O(N__32740),
            .I(N__32737));
    LocalMux I__5579 (
            .O(N__32737),
            .I(\ADC_VDC.n22067 ));
    CascadeMux I__5578 (
            .O(N__32734),
            .I(N__32719));
    CascadeMux I__5577 (
            .O(N__32733),
            .I(N__32716));
    InMux I__5576 (
            .O(N__32732),
            .I(N__32704));
    InMux I__5575 (
            .O(N__32731),
            .I(N__32697));
    InMux I__5574 (
            .O(N__32730),
            .I(N__32689));
    InMux I__5573 (
            .O(N__32729),
            .I(N__32689));
    InMux I__5572 (
            .O(N__32728),
            .I(N__32689));
    InMux I__5571 (
            .O(N__32727),
            .I(N__32679));
    InMux I__5570 (
            .O(N__32726),
            .I(N__32679));
    InMux I__5569 (
            .O(N__32725),
            .I(N__32679));
    InMux I__5568 (
            .O(N__32724),
            .I(N__32679));
    InMux I__5567 (
            .O(N__32723),
            .I(N__32674));
    InMux I__5566 (
            .O(N__32722),
            .I(N__32674));
    InMux I__5565 (
            .O(N__32719),
            .I(N__32665));
    InMux I__5564 (
            .O(N__32716),
            .I(N__32665));
    InMux I__5563 (
            .O(N__32715),
            .I(N__32665));
    InMux I__5562 (
            .O(N__32714),
            .I(N__32665));
    InMux I__5561 (
            .O(N__32713),
            .I(N__32650));
    InMux I__5560 (
            .O(N__32712),
            .I(N__32650));
    InMux I__5559 (
            .O(N__32711),
            .I(N__32650));
    InMux I__5558 (
            .O(N__32710),
            .I(N__32650));
    InMux I__5557 (
            .O(N__32709),
            .I(N__32650));
    InMux I__5556 (
            .O(N__32708),
            .I(N__32650));
    InMux I__5555 (
            .O(N__32707),
            .I(N__32650));
    LocalMux I__5554 (
            .O(N__32704),
            .I(N__32647));
    InMux I__5553 (
            .O(N__32703),
            .I(N__32642));
    InMux I__5552 (
            .O(N__32702),
            .I(N__32642));
    InMux I__5551 (
            .O(N__32701),
            .I(N__32638));
    InMux I__5550 (
            .O(N__32700),
            .I(N__32635));
    LocalMux I__5549 (
            .O(N__32697),
            .I(N__32632));
    InMux I__5548 (
            .O(N__32696),
            .I(N__32629));
    LocalMux I__5547 (
            .O(N__32689),
            .I(N__32626));
    InMux I__5546 (
            .O(N__32688),
            .I(N__32623));
    LocalMux I__5545 (
            .O(N__32679),
            .I(N__32608));
    LocalMux I__5544 (
            .O(N__32674),
            .I(N__32608));
    LocalMux I__5543 (
            .O(N__32665),
            .I(N__32608));
    LocalMux I__5542 (
            .O(N__32650),
            .I(N__32608));
    Span4Mux_h I__5541 (
            .O(N__32647),
            .I(N__32600));
    LocalMux I__5540 (
            .O(N__32642),
            .I(N__32600));
    CascadeMux I__5539 (
            .O(N__32641),
            .I(N__32592));
    LocalMux I__5538 (
            .O(N__32638),
            .I(N__32577));
    LocalMux I__5537 (
            .O(N__32635),
            .I(N__32577));
    Span4Mux_h I__5536 (
            .O(N__32632),
            .I(N__32577));
    LocalMux I__5535 (
            .O(N__32629),
            .I(N__32577));
    Span4Mux_v I__5534 (
            .O(N__32626),
            .I(N__32577));
    LocalMux I__5533 (
            .O(N__32623),
            .I(N__32577));
    InMux I__5532 (
            .O(N__32622),
            .I(N__32564));
    InMux I__5531 (
            .O(N__32621),
            .I(N__32564));
    InMux I__5530 (
            .O(N__32620),
            .I(N__32564));
    InMux I__5529 (
            .O(N__32619),
            .I(N__32564));
    InMux I__5528 (
            .O(N__32618),
            .I(N__32564));
    InMux I__5527 (
            .O(N__32617),
            .I(N__32564));
    Span4Mux_v I__5526 (
            .O(N__32608),
            .I(N__32561));
    InMux I__5525 (
            .O(N__32607),
            .I(N__32556));
    InMux I__5524 (
            .O(N__32606),
            .I(N__32556));
    InMux I__5523 (
            .O(N__32605),
            .I(N__32553));
    Span4Mux_h I__5522 (
            .O(N__32600),
            .I(N__32550));
    InMux I__5521 (
            .O(N__32599),
            .I(N__32543));
    InMux I__5520 (
            .O(N__32598),
            .I(N__32543));
    InMux I__5519 (
            .O(N__32597),
            .I(N__32543));
    InMux I__5518 (
            .O(N__32596),
            .I(N__32536));
    InMux I__5517 (
            .O(N__32595),
            .I(N__32536));
    InMux I__5516 (
            .O(N__32592),
            .I(N__32536));
    InMux I__5515 (
            .O(N__32591),
            .I(N__32531));
    InMux I__5514 (
            .O(N__32590),
            .I(N__32531));
    Span4Mux_v I__5513 (
            .O(N__32577),
            .I(N__32528));
    LocalMux I__5512 (
            .O(N__32564),
            .I(adc_state_3));
    Odrv4 I__5511 (
            .O(N__32561),
            .I(adc_state_3));
    LocalMux I__5510 (
            .O(N__32556),
            .I(adc_state_3));
    LocalMux I__5509 (
            .O(N__32553),
            .I(adc_state_3));
    Odrv4 I__5508 (
            .O(N__32550),
            .I(adc_state_3));
    LocalMux I__5507 (
            .O(N__32543),
            .I(adc_state_3));
    LocalMux I__5506 (
            .O(N__32536),
            .I(adc_state_3));
    LocalMux I__5505 (
            .O(N__32531),
            .I(adc_state_3));
    Odrv4 I__5504 (
            .O(N__32528),
            .I(adc_state_3));
    InMux I__5503 (
            .O(N__32509),
            .I(N__32498));
    InMux I__5502 (
            .O(N__32508),
            .I(N__32498));
    InMux I__5501 (
            .O(N__32507),
            .I(N__32498));
    InMux I__5500 (
            .O(N__32506),
            .I(N__32491));
    InMux I__5499 (
            .O(N__32505),
            .I(N__32487));
    LocalMux I__5498 (
            .O(N__32498),
            .I(N__32481));
    InMux I__5497 (
            .O(N__32497),
            .I(N__32478));
    InMux I__5496 (
            .O(N__32496),
            .I(N__32473));
    InMux I__5495 (
            .O(N__32495),
            .I(N__32473));
    InMux I__5494 (
            .O(N__32494),
            .I(N__32467));
    LocalMux I__5493 (
            .O(N__32491),
            .I(N__32464));
    InMux I__5492 (
            .O(N__32490),
            .I(N__32461));
    LocalMux I__5491 (
            .O(N__32487),
            .I(N__32454));
    InMux I__5490 (
            .O(N__32486),
            .I(N__32451));
    InMux I__5489 (
            .O(N__32485),
            .I(N__32447));
    InMux I__5488 (
            .O(N__32484),
            .I(N__32444));
    Sp12to4 I__5487 (
            .O(N__32481),
            .I(N__32441));
    LocalMux I__5486 (
            .O(N__32478),
            .I(N__32438));
    LocalMux I__5485 (
            .O(N__32473),
            .I(N__32435));
    InMux I__5484 (
            .O(N__32472),
            .I(N__32428));
    InMux I__5483 (
            .O(N__32471),
            .I(N__32428));
    InMux I__5482 (
            .O(N__32470),
            .I(N__32428));
    LocalMux I__5481 (
            .O(N__32467),
            .I(N__32421));
    Span4Mux_h I__5480 (
            .O(N__32464),
            .I(N__32421));
    LocalMux I__5479 (
            .O(N__32461),
            .I(N__32421));
    InMux I__5478 (
            .O(N__32460),
            .I(N__32414));
    InMux I__5477 (
            .O(N__32459),
            .I(N__32414));
    InMux I__5476 (
            .O(N__32458),
            .I(N__32414));
    InMux I__5475 (
            .O(N__32457),
            .I(N__32411));
    Span4Mux_v I__5474 (
            .O(N__32454),
            .I(N__32406));
    LocalMux I__5473 (
            .O(N__32451),
            .I(N__32406));
    InMux I__5472 (
            .O(N__32450),
            .I(N__32403));
    LocalMux I__5471 (
            .O(N__32447),
            .I(adc_state_1_adj_1551));
    LocalMux I__5470 (
            .O(N__32444),
            .I(adc_state_1_adj_1551));
    Odrv12 I__5469 (
            .O(N__32441),
            .I(adc_state_1_adj_1551));
    Odrv4 I__5468 (
            .O(N__32438),
            .I(adc_state_1_adj_1551));
    Odrv4 I__5467 (
            .O(N__32435),
            .I(adc_state_1_adj_1551));
    LocalMux I__5466 (
            .O(N__32428),
            .I(adc_state_1_adj_1551));
    Odrv4 I__5465 (
            .O(N__32421),
            .I(adc_state_1_adj_1551));
    LocalMux I__5464 (
            .O(N__32414),
            .I(adc_state_1_adj_1551));
    LocalMux I__5463 (
            .O(N__32411),
            .I(adc_state_1_adj_1551));
    Odrv4 I__5462 (
            .O(N__32406),
            .I(adc_state_1_adj_1551));
    LocalMux I__5461 (
            .O(N__32403),
            .I(adc_state_1_adj_1551));
    CascadeMux I__5460 (
            .O(N__32380),
            .I(N__32377));
    InMux I__5459 (
            .O(N__32377),
            .I(N__32373));
    CascadeMux I__5458 (
            .O(N__32376),
            .I(N__32369));
    LocalMux I__5457 (
            .O(N__32373),
            .I(N__32366));
    InMux I__5456 (
            .O(N__32372),
            .I(N__32363));
    InMux I__5455 (
            .O(N__32369),
            .I(N__32360));
    Span4Mux_v I__5454 (
            .O(N__32366),
            .I(N__32357));
    LocalMux I__5453 (
            .O(N__32363),
            .I(N__32354));
    LocalMux I__5452 (
            .O(N__32360),
            .I(buf_dds0_5));
    Odrv4 I__5451 (
            .O(N__32357),
            .I(buf_dds0_5));
    Odrv12 I__5450 (
            .O(N__32354),
            .I(buf_dds0_5));
    InMux I__5449 (
            .O(N__32347),
            .I(N__32344));
    LocalMux I__5448 (
            .O(N__32344),
            .I(\SIG_DDS.tmp_buf_4 ));
    CascadeMux I__5447 (
            .O(N__32341),
            .I(N__32338));
    InMux I__5446 (
            .O(N__32338),
            .I(N__32335));
    LocalMux I__5445 (
            .O(N__32335),
            .I(\SIG_DDS.tmp_buf_5 ));
    CascadeMux I__5444 (
            .O(N__32332),
            .I(N__32329));
    InMux I__5443 (
            .O(N__32329),
            .I(N__32326));
    LocalMux I__5442 (
            .O(N__32326),
            .I(\SIG_DDS.tmp_buf_9 ));
    CascadeMux I__5441 (
            .O(N__32323),
            .I(N__32320));
    InMux I__5440 (
            .O(N__32320),
            .I(N__32317));
    LocalMux I__5439 (
            .O(N__32317),
            .I(\SIG_DDS.tmp_buf_6 ));
    InMux I__5438 (
            .O(N__32314),
            .I(N__32309));
    InMux I__5437 (
            .O(N__32313),
            .I(N__32306));
    InMux I__5436 (
            .O(N__32312),
            .I(N__32303));
    LocalMux I__5435 (
            .O(N__32309),
            .I(N__32300));
    LocalMux I__5434 (
            .O(N__32306),
            .I(buf_dds0_7));
    LocalMux I__5433 (
            .O(N__32303),
            .I(buf_dds0_7));
    Odrv4 I__5432 (
            .O(N__32300),
            .I(buf_dds0_7));
    CascadeMux I__5431 (
            .O(N__32293),
            .I(N__32290));
    InMux I__5430 (
            .O(N__32290),
            .I(N__32287));
    LocalMux I__5429 (
            .O(N__32287),
            .I(N__32284));
    Span4Mux_v I__5428 (
            .O(N__32284),
            .I(N__32279));
    InMux I__5427 (
            .O(N__32283),
            .I(N__32276));
    InMux I__5426 (
            .O(N__32282),
            .I(N__32273));
    Span4Mux_h I__5425 (
            .O(N__32279),
            .I(N__32270));
    LocalMux I__5424 (
            .O(N__32276),
            .I(N__32267));
    LocalMux I__5423 (
            .O(N__32273),
            .I(buf_dds0_12));
    Odrv4 I__5422 (
            .O(N__32270),
            .I(buf_dds0_12));
    Odrv4 I__5421 (
            .O(N__32267),
            .I(buf_dds0_12));
    CascadeMux I__5420 (
            .O(N__32260),
            .I(N__32257));
    InMux I__5419 (
            .O(N__32257),
            .I(N__32254));
    LocalMux I__5418 (
            .O(N__32254),
            .I(\SIG_DDS.tmp_buf_12 ));
    CascadeMux I__5417 (
            .O(N__32251),
            .I(N__32248));
    InMux I__5416 (
            .O(N__32248),
            .I(N__32245));
    LocalMux I__5415 (
            .O(N__32245),
            .I(\SIG_DDS.tmp_buf_13 ));
    InMux I__5414 (
            .O(N__32242),
            .I(N__32239));
    LocalMux I__5413 (
            .O(N__32239),
            .I(N__32236));
    Span4Mux_h I__5412 (
            .O(N__32236),
            .I(N__32232));
    InMux I__5411 (
            .O(N__32235),
            .I(N__32228));
    Span4Mux_v I__5410 (
            .O(N__32232),
            .I(N__32225));
    InMux I__5409 (
            .O(N__32231),
            .I(N__32222));
    LocalMux I__5408 (
            .O(N__32228),
            .I(N__32219));
    Odrv4 I__5407 (
            .O(N__32225),
            .I(buf_dds0_14));
    LocalMux I__5406 (
            .O(N__32222),
            .I(buf_dds0_14));
    Odrv4 I__5405 (
            .O(N__32219),
            .I(buf_dds0_14));
    CascadeMux I__5404 (
            .O(N__32212),
            .I(N__32209));
    InMux I__5403 (
            .O(N__32209),
            .I(N__32206));
    LocalMux I__5402 (
            .O(N__32206),
            .I(\SIG_DDS.tmp_buf_14 ));
    CascadeMux I__5401 (
            .O(N__32203),
            .I(N__32200));
    InMux I__5400 (
            .O(N__32200),
            .I(N__32197));
    LocalMux I__5399 (
            .O(N__32197),
            .I(N__32192));
    InMux I__5398 (
            .O(N__32196),
            .I(N__32189));
    InMux I__5397 (
            .O(N__32195),
            .I(N__32186));
    Span4Mux_h I__5396 (
            .O(N__32192),
            .I(N__32183));
    LocalMux I__5395 (
            .O(N__32189),
            .I(buf_dds0_15));
    LocalMux I__5394 (
            .O(N__32186),
            .I(buf_dds0_15));
    Odrv4 I__5393 (
            .O(N__32183),
            .I(buf_dds0_15));
    InMux I__5392 (
            .O(N__32176),
            .I(N__32173));
    LocalMux I__5391 (
            .O(N__32173),
            .I(\SIG_DDS.tmp_buf_7 ));
    CascadeMux I__5390 (
            .O(N__32170),
            .I(N__32167));
    InMux I__5389 (
            .O(N__32167),
            .I(N__32164));
    LocalMux I__5388 (
            .O(N__32164),
            .I(\SIG_DDS.tmp_buf_8 ));
    InMux I__5387 (
            .O(N__32161),
            .I(N__32157));
    InMux I__5386 (
            .O(N__32160),
            .I(N__32154));
    LocalMux I__5385 (
            .O(N__32157),
            .I(cmd_rdadctmp_6));
    LocalMux I__5384 (
            .O(N__32154),
            .I(cmd_rdadctmp_6));
    CascadeMux I__5383 (
            .O(N__32149),
            .I(N__32143));
    InMux I__5382 (
            .O(N__32148),
            .I(N__32137));
    InMux I__5381 (
            .O(N__32147),
            .I(N__32137));
    InMux I__5380 (
            .O(N__32146),
            .I(N__32132));
    InMux I__5379 (
            .O(N__32143),
            .I(N__32132));
    InMux I__5378 (
            .O(N__32142),
            .I(N__32129));
    LocalMux I__5377 (
            .O(N__32137),
            .I(acadc_dtrig_i));
    LocalMux I__5376 (
            .O(N__32132),
            .I(acadc_dtrig_i));
    LocalMux I__5375 (
            .O(N__32129),
            .I(acadc_dtrig_i));
    CascadeMux I__5374 (
            .O(N__32122),
            .I(N__32118));
    CascadeMux I__5373 (
            .O(N__32121),
            .I(N__32115));
    InMux I__5372 (
            .O(N__32118),
            .I(N__32109));
    InMux I__5371 (
            .O(N__32115),
            .I(N__32109));
    InMux I__5370 (
            .O(N__32114),
            .I(N__32106));
    LocalMux I__5369 (
            .O(N__32109),
            .I(cmd_rdadctmp_29));
    LocalMux I__5368 (
            .O(N__32106),
            .I(cmd_rdadctmp_29));
    InMux I__5367 (
            .O(N__32101),
            .I(N__32096));
    CascadeMux I__5366 (
            .O(N__32100),
            .I(N__32086));
    InMux I__5365 (
            .O(N__32099),
            .I(N__32083));
    LocalMux I__5364 (
            .O(N__32096),
            .I(N__32080));
    InMux I__5363 (
            .O(N__32095),
            .I(N__32073));
    InMux I__5362 (
            .O(N__32094),
            .I(N__32073));
    InMux I__5361 (
            .O(N__32093),
            .I(N__32073));
    CascadeMux I__5360 (
            .O(N__32092),
            .I(N__32068));
    InMux I__5359 (
            .O(N__32091),
            .I(N__32061));
    InMux I__5358 (
            .O(N__32090),
            .I(N__32061));
    InMux I__5357 (
            .O(N__32089),
            .I(N__32056));
    InMux I__5356 (
            .O(N__32086),
            .I(N__32056));
    LocalMux I__5355 (
            .O(N__32083),
            .I(N__32053));
    Span4Mux_v I__5354 (
            .O(N__32080),
            .I(N__32050));
    LocalMux I__5353 (
            .O(N__32073),
            .I(N__32047));
    InMux I__5352 (
            .O(N__32072),
            .I(N__32044));
    InMux I__5351 (
            .O(N__32071),
            .I(N__32039));
    InMux I__5350 (
            .O(N__32068),
            .I(N__32039));
    InMux I__5349 (
            .O(N__32067),
            .I(N__32034));
    InMux I__5348 (
            .O(N__32066),
            .I(N__32034));
    LocalMux I__5347 (
            .O(N__32061),
            .I(N__32029));
    LocalMux I__5346 (
            .O(N__32056),
            .I(N__32029));
    Span4Mux_v I__5345 (
            .O(N__32053),
            .I(N__32020));
    Span4Mux_h I__5344 (
            .O(N__32050),
            .I(N__32020));
    Span4Mux_h I__5343 (
            .O(N__32047),
            .I(N__32020));
    LocalMux I__5342 (
            .O(N__32044),
            .I(N__32020));
    LocalMux I__5341 (
            .O(N__32039),
            .I(DTRIG_N_1182_adj_1549));
    LocalMux I__5340 (
            .O(N__32034),
            .I(DTRIG_N_1182_adj_1549));
    Odrv4 I__5339 (
            .O(N__32029),
            .I(DTRIG_N_1182_adj_1549));
    Odrv4 I__5338 (
            .O(N__32020),
            .I(DTRIG_N_1182_adj_1549));
    CascadeMux I__5337 (
            .O(N__32011),
            .I(N__32008));
    InMux I__5336 (
            .O(N__32008),
            .I(N__32005));
    LocalMux I__5335 (
            .O(N__32005),
            .I(N__32001));
    InMux I__5334 (
            .O(N__32004),
            .I(N__31993));
    Span4Mux_v I__5333 (
            .O(N__32001),
            .I(N__31988));
    InMux I__5332 (
            .O(N__32000),
            .I(N__31981));
    InMux I__5331 (
            .O(N__31999),
            .I(N__31981));
    InMux I__5330 (
            .O(N__31998),
            .I(N__31981));
    InMux I__5329 (
            .O(N__31997),
            .I(N__31976));
    InMux I__5328 (
            .O(N__31996),
            .I(N__31976));
    LocalMux I__5327 (
            .O(N__31993),
            .I(N__31973));
    InMux I__5326 (
            .O(N__31992),
            .I(N__31967));
    InMux I__5325 (
            .O(N__31991),
            .I(N__31964));
    Span4Mux_h I__5324 (
            .O(N__31988),
            .I(N__31958));
    LocalMux I__5323 (
            .O(N__31981),
            .I(N__31958));
    LocalMux I__5322 (
            .O(N__31976),
            .I(N__31953));
    Span4Mux_h I__5321 (
            .O(N__31973),
            .I(N__31953));
    InMux I__5320 (
            .O(N__31972),
            .I(N__31948));
    InMux I__5319 (
            .O(N__31971),
            .I(N__31948));
    InMux I__5318 (
            .O(N__31970),
            .I(N__31945));
    LocalMux I__5317 (
            .O(N__31967),
            .I(N__31940));
    LocalMux I__5316 (
            .O(N__31964),
            .I(N__31940));
    InMux I__5315 (
            .O(N__31963),
            .I(N__31937));
    Span4Mux_h I__5314 (
            .O(N__31958),
            .I(N__31934));
    Span4Mux_h I__5313 (
            .O(N__31953),
            .I(N__31931));
    LocalMux I__5312 (
            .O(N__31948),
            .I(adc_state_1_adj_1515));
    LocalMux I__5311 (
            .O(N__31945),
            .I(adc_state_1_adj_1515));
    Odrv4 I__5310 (
            .O(N__31940),
            .I(adc_state_1_adj_1515));
    LocalMux I__5309 (
            .O(N__31937),
            .I(adc_state_1_adj_1515));
    Odrv4 I__5308 (
            .O(N__31934),
            .I(adc_state_1_adj_1515));
    Odrv4 I__5307 (
            .O(N__31931),
            .I(adc_state_1_adj_1515));
    CascadeMux I__5306 (
            .O(N__31918),
            .I(N__31915));
    InMux I__5305 (
            .O(N__31915),
            .I(N__31906));
    InMux I__5304 (
            .O(N__31914),
            .I(N__31906));
    InMux I__5303 (
            .O(N__31913),
            .I(N__31901));
    InMux I__5302 (
            .O(N__31912),
            .I(N__31901));
    InMux I__5301 (
            .O(N__31911),
            .I(N__31898));
    LocalMux I__5300 (
            .O(N__31906),
            .I(acadc_dtrig_v));
    LocalMux I__5299 (
            .O(N__31901),
            .I(acadc_dtrig_v));
    LocalMux I__5298 (
            .O(N__31898),
            .I(acadc_dtrig_v));
    InMux I__5297 (
            .O(N__31891),
            .I(N__31887));
    InMux I__5296 (
            .O(N__31890),
            .I(N__31884));
    LocalMux I__5295 (
            .O(N__31887),
            .I(N__31881));
    LocalMux I__5294 (
            .O(N__31884),
            .I(N__31878));
    Span4Mux_h I__5293 (
            .O(N__31881),
            .I(N__31872));
    Span4Mux_h I__5292 (
            .O(N__31878),
            .I(N__31872));
    InMux I__5291 (
            .O(N__31877),
            .I(N__31869));
    Span4Mux_v I__5290 (
            .O(N__31872),
            .I(N__31866));
    LocalMux I__5289 (
            .O(N__31869),
            .I(buf_dds1_9));
    Odrv4 I__5288 (
            .O(N__31866),
            .I(buf_dds1_9));
    InMux I__5287 (
            .O(N__31861),
            .I(N__31858));
    LocalMux I__5286 (
            .O(N__31858),
            .I(n23534));
    InMux I__5285 (
            .O(N__31855),
            .I(N__31850));
    InMux I__5284 (
            .O(N__31854),
            .I(N__31845));
    InMux I__5283 (
            .O(N__31853),
            .I(N__31845));
    LocalMux I__5282 (
            .O(N__31850),
            .I(buf_dds0_10));
    LocalMux I__5281 (
            .O(N__31845),
            .I(buf_dds0_10));
    InMux I__5280 (
            .O(N__31840),
            .I(N__31836));
    InMux I__5279 (
            .O(N__31839),
            .I(N__31833));
    LocalMux I__5278 (
            .O(N__31836),
            .I(N__31830));
    LocalMux I__5277 (
            .O(N__31833),
            .I(N__31826));
    Span4Mux_v I__5276 (
            .O(N__31830),
            .I(N__31823));
    InMux I__5275 (
            .O(N__31829),
            .I(N__31820));
    Span4Mux_v I__5274 (
            .O(N__31826),
            .I(N__31817));
    Odrv4 I__5273 (
            .O(N__31823),
            .I(buf_dds0_6));
    LocalMux I__5272 (
            .O(N__31820),
            .I(buf_dds0_6));
    Odrv4 I__5271 (
            .O(N__31817),
            .I(buf_dds0_6));
    CascadeMux I__5270 (
            .O(N__31810),
            .I(n13_cascade_));
    InMux I__5269 (
            .O(N__31807),
            .I(N__31804));
    LocalMux I__5268 (
            .O(N__31804),
            .I(n22395));
    CascadeMux I__5267 (
            .O(N__31801),
            .I(N__31798));
    InMux I__5266 (
            .O(N__31798),
            .I(N__31794));
    InMux I__5265 (
            .O(N__31797),
            .I(N__31791));
    LocalMux I__5264 (
            .O(N__31794),
            .I(N__31788));
    LocalMux I__5263 (
            .O(N__31791),
            .I(N__31785));
    Span4Mux_v I__5262 (
            .O(N__31788),
            .I(N__31782));
    Span4Mux_v I__5261 (
            .O(N__31785),
            .I(N__31779));
    Span4Mux_h I__5260 (
            .O(N__31782),
            .I(N__31775));
    Span4Mux_h I__5259 (
            .O(N__31779),
            .I(N__31772));
    InMux I__5258 (
            .O(N__31778),
            .I(N__31769));
    Odrv4 I__5257 (
            .O(N__31775),
            .I(cmd_rdadctmp_30));
    Odrv4 I__5256 (
            .O(N__31772),
            .I(cmd_rdadctmp_30));
    LocalMux I__5255 (
            .O(N__31769),
            .I(cmd_rdadctmp_30));
    InMux I__5254 (
            .O(N__31762),
            .I(N__31758));
    InMux I__5253 (
            .O(N__31761),
            .I(N__31755));
    LocalMux I__5252 (
            .O(N__31758),
            .I(N__31752));
    LocalMux I__5251 (
            .O(N__31755),
            .I(n13_adj_1591));
    Odrv4 I__5250 (
            .O(N__31752),
            .I(n13_adj_1591));
    InMux I__5249 (
            .O(N__31747),
            .I(N__31744));
    LocalMux I__5248 (
            .O(N__31744),
            .I(n11_adj_1592));
    CascadeMux I__5247 (
            .O(N__31741),
            .I(n23510_cascade_));
    InMux I__5246 (
            .O(N__31738),
            .I(N__31735));
    LocalMux I__5245 (
            .O(N__31735),
            .I(N__31732));
    Odrv12 I__5244 (
            .O(N__31732),
            .I(n22276));
    CascadeMux I__5243 (
            .O(N__31729),
            .I(n23513_cascade_));
    CascadeMux I__5242 (
            .O(N__31726),
            .I(n30_adj_1759_cascade_));
    InMux I__5241 (
            .O(N__31723),
            .I(N__31720));
    LocalMux I__5240 (
            .O(N__31720),
            .I(n26_adj_1758));
    InMux I__5239 (
            .O(N__31717),
            .I(N__31711));
    InMux I__5238 (
            .O(N__31716),
            .I(N__31711));
    LocalMux I__5237 (
            .O(N__31711),
            .I(eis_end));
    InMux I__5236 (
            .O(N__31708),
            .I(N__31705));
    LocalMux I__5235 (
            .O(N__31705),
            .I(n112_adj_1762));
    CascadeMux I__5234 (
            .O(N__31702),
            .I(n21946_cascade_));
    InMux I__5233 (
            .O(N__31699),
            .I(N__31696));
    LocalMux I__5232 (
            .O(N__31696),
            .I(n21880));
    CascadeMux I__5231 (
            .O(N__31693),
            .I(n24_cascade_));
    InMux I__5230 (
            .O(N__31690),
            .I(N__31687));
    LocalMux I__5229 (
            .O(N__31687),
            .I(N__31684));
    Span12Mux_s8_v I__5228 (
            .O(N__31684),
            .I(N__31680));
    InMux I__5227 (
            .O(N__31683),
            .I(N__31677));
    Span12Mux_h I__5226 (
            .O(N__31680),
            .I(N__31673));
    LocalMux I__5225 (
            .O(N__31677),
            .I(N__31670));
    InMux I__5224 (
            .O(N__31676),
            .I(N__31667));
    Span12Mux_v I__5223 (
            .O(N__31673),
            .I(N__31664));
    Span4Mux_h I__5222 (
            .O(N__31670),
            .I(N__31661));
    LocalMux I__5221 (
            .O(N__31667),
            .I(buf_adcdata_iac_22));
    Odrv12 I__5220 (
            .O(N__31664),
            .I(buf_adcdata_iac_22));
    Odrv4 I__5219 (
            .O(N__31661),
            .I(buf_adcdata_iac_22));
    IoInMux I__5218 (
            .O(N__31654),
            .I(N__31651));
    LocalMux I__5217 (
            .O(N__31651),
            .I(N__31648));
    Span12Mux_s1_h I__5216 (
            .O(N__31648),
            .I(N__31645));
    Span12Mux_h I__5215 (
            .O(N__31645),
            .I(N__31640));
    InMux I__5214 (
            .O(N__31644),
            .I(N__31635));
    InMux I__5213 (
            .O(N__31643),
            .I(N__31635));
    Odrv12 I__5212 (
            .O(N__31640),
            .I(VAC_FLT0));
    LocalMux I__5211 (
            .O(N__31635),
            .I(VAC_FLT0));
    InMux I__5210 (
            .O(N__31630),
            .I(N__31627));
    LocalMux I__5209 (
            .O(N__31627),
            .I(N__31624));
    Odrv4 I__5208 (
            .O(N__31624),
            .I(n17_adj_1764));
    CascadeMux I__5207 (
            .O(N__31621),
            .I(n11981_cascade_));
    IoInMux I__5206 (
            .O(N__31618),
            .I(N__31615));
    LocalMux I__5205 (
            .O(N__31615),
            .I(N__31612));
    IoSpan4Mux I__5204 (
            .O(N__31612),
            .I(N__31609));
    Span4Mux_s3_h I__5203 (
            .O(N__31609),
            .I(N__31606));
    Span4Mux_h I__5202 (
            .O(N__31606),
            .I(N__31603));
    Span4Mux_h I__5201 (
            .O(N__31603),
            .I(N__31599));
    InMux I__5200 (
            .O(N__31602),
            .I(N__31596));
    Span4Mux_v I__5199 (
            .O(N__31599),
            .I(N__31590));
    LocalMux I__5198 (
            .O(N__31596),
            .I(N__31590));
    InMux I__5197 (
            .O(N__31595),
            .I(N__31587));
    Span4Mux_v I__5196 (
            .O(N__31590),
            .I(N__31584));
    LocalMux I__5195 (
            .O(N__31587),
            .I(VAC_FLT1));
    Odrv4 I__5194 (
            .O(N__31584),
            .I(VAC_FLT1));
    InMux I__5193 (
            .O(N__31579),
            .I(N__31576));
    LocalMux I__5192 (
            .O(N__31576),
            .I(n24_adj_1576));
    InMux I__5191 (
            .O(N__31573),
            .I(N__31570));
    LocalMux I__5190 (
            .O(N__31570),
            .I(n11986));
    InMux I__5189 (
            .O(N__31567),
            .I(N__31564));
    LocalMux I__5188 (
            .O(N__31564),
            .I(N__31561));
    Span4Mux_h I__5187 (
            .O(N__31561),
            .I(N__31558));
    Odrv4 I__5186 (
            .O(N__31558),
            .I(n30_adj_1692));
    CascadeMux I__5185 (
            .O(N__31555),
            .I(N__31552));
    InMux I__5184 (
            .O(N__31552),
            .I(N__31548));
    CascadeMux I__5183 (
            .O(N__31551),
            .I(N__31544));
    LocalMux I__5182 (
            .O(N__31548),
            .I(N__31541));
    CascadeMux I__5181 (
            .O(N__31547),
            .I(N__31538));
    InMux I__5180 (
            .O(N__31544),
            .I(N__31535));
    Span4Mux_h I__5179 (
            .O(N__31541),
            .I(N__31532));
    InMux I__5178 (
            .O(N__31538),
            .I(N__31529));
    LocalMux I__5177 (
            .O(N__31535),
            .I(N__31526));
    Span4Mux_h I__5176 (
            .O(N__31532),
            .I(N__31523));
    LocalMux I__5175 (
            .O(N__31529),
            .I(cmd_rdadctmp_25_adj_1523));
    Odrv12 I__5174 (
            .O(N__31526),
            .I(cmd_rdadctmp_25_adj_1523));
    Odrv4 I__5173 (
            .O(N__31523),
            .I(cmd_rdadctmp_25_adj_1523));
    InMux I__5172 (
            .O(N__31516),
            .I(N__31513));
    LocalMux I__5171 (
            .O(N__31513),
            .I(N__31509));
    CascadeMux I__5170 (
            .O(N__31512),
            .I(N__31506));
    Span4Mux_h I__5169 (
            .O(N__31509),
            .I(N__31503));
    InMux I__5168 (
            .O(N__31506),
            .I(N__31500));
    Odrv4 I__5167 (
            .O(N__31503),
            .I(buf_adcdata_vdc_18));
    LocalMux I__5166 (
            .O(N__31500),
            .I(buf_adcdata_vdc_18));
    InMux I__5165 (
            .O(N__31495),
            .I(N__31492));
    LocalMux I__5164 (
            .O(N__31492),
            .I(N__31489));
    Span4Mux_v I__5163 (
            .O(N__31489),
            .I(N__31486));
    Sp12to4 I__5162 (
            .O(N__31486),
            .I(N__31481));
    InMux I__5161 (
            .O(N__31485),
            .I(N__31478));
    InMux I__5160 (
            .O(N__31484),
            .I(N__31475));
    Span12Mux_h I__5159 (
            .O(N__31481),
            .I(N__31472));
    LocalMux I__5158 (
            .O(N__31478),
            .I(N__31469));
    LocalMux I__5157 (
            .O(N__31475),
            .I(buf_adcdata_vac_18));
    Odrv12 I__5156 (
            .O(N__31472),
            .I(buf_adcdata_vac_18));
    Odrv4 I__5155 (
            .O(N__31469),
            .I(buf_adcdata_vac_18));
    InMux I__5154 (
            .O(N__31462),
            .I(N__31459));
    LocalMux I__5153 (
            .O(N__31459),
            .I(n22163));
    InMux I__5152 (
            .O(N__31456),
            .I(N__31453));
    LocalMux I__5151 (
            .O(N__31453),
            .I(N__31449));
    InMux I__5150 (
            .O(N__31452),
            .I(N__31446));
    Odrv4 I__5149 (
            .O(N__31449),
            .I(\comm_spi.n15360 ));
    LocalMux I__5148 (
            .O(N__31446),
            .I(\comm_spi.n15360 ));
    SRMux I__5147 (
            .O(N__31441),
            .I(N__31438));
    LocalMux I__5146 (
            .O(N__31438),
            .I(N__31435));
    Odrv4 I__5145 (
            .O(N__31435),
            .I(\comm_spi.data_tx_7__N_857 ));
    InMux I__5144 (
            .O(N__31432),
            .I(N__31428));
    InMux I__5143 (
            .O(N__31431),
            .I(N__31425));
    LocalMux I__5142 (
            .O(N__31428),
            .I(N__31422));
    LocalMux I__5141 (
            .O(N__31425),
            .I(comm_test_buf_24_19));
    Odrv4 I__5140 (
            .O(N__31422),
            .I(comm_test_buf_24_19));
    InMux I__5139 (
            .O(N__31417),
            .I(N__31413));
    InMux I__5138 (
            .O(N__31416),
            .I(N__31410));
    LocalMux I__5137 (
            .O(N__31413),
            .I(comm_test_buf_24_20));
    LocalMux I__5136 (
            .O(N__31410),
            .I(comm_test_buf_24_20));
    InMux I__5135 (
            .O(N__31405),
            .I(N__31402));
    LocalMux I__5134 (
            .O(N__31402),
            .I(N__31399));
    Span4Mux_v I__5133 (
            .O(N__31399),
            .I(N__31396));
    Odrv4 I__5132 (
            .O(N__31396),
            .I(n111_adj_1785));
    CascadeMux I__5131 (
            .O(N__31393),
            .I(N__31390));
    InMux I__5130 (
            .O(N__31390),
            .I(N__31384));
    InMux I__5129 (
            .O(N__31389),
            .I(N__31384));
    LocalMux I__5128 (
            .O(N__31384),
            .I(cmd_rdadctmp_7_adj_1541));
    CascadeMux I__5127 (
            .O(N__31381),
            .I(N__31378));
    InMux I__5126 (
            .O(N__31378),
            .I(N__31372));
    InMux I__5125 (
            .O(N__31377),
            .I(N__31372));
    LocalMux I__5124 (
            .O(N__31372),
            .I(cmd_rdadctmp_6_adj_1542));
    CascadeMux I__5123 (
            .O(N__31369),
            .I(N__31366));
    InMux I__5122 (
            .O(N__31366),
            .I(N__31360));
    InMux I__5121 (
            .O(N__31365),
            .I(N__31360));
    LocalMux I__5120 (
            .O(N__31360),
            .I(cmd_rdadctmp_5_adj_1543));
    CascadeMux I__5119 (
            .O(N__31357),
            .I(N__31353));
    InMux I__5118 (
            .O(N__31356),
            .I(N__31350));
    InMux I__5117 (
            .O(N__31353),
            .I(N__31347));
    LocalMux I__5116 (
            .O(N__31350),
            .I(N__31344));
    LocalMux I__5115 (
            .O(N__31347),
            .I(cmd_rdadctmp_3_adj_1545));
    Odrv12 I__5114 (
            .O(N__31344),
            .I(cmd_rdadctmp_3_adj_1545));
    CascadeMux I__5113 (
            .O(N__31339),
            .I(N__31336));
    InMux I__5112 (
            .O(N__31336),
            .I(N__31330));
    InMux I__5111 (
            .O(N__31335),
            .I(N__31330));
    LocalMux I__5110 (
            .O(N__31330),
            .I(cmd_rdadctmp_4_adj_1544));
    InMux I__5109 (
            .O(N__31327),
            .I(N__31324));
    LocalMux I__5108 (
            .O(N__31324),
            .I(N__31319));
    InMux I__5107 (
            .O(N__31323),
            .I(N__31316));
    InMux I__5106 (
            .O(N__31322),
            .I(N__31313));
    Span4Mux_v I__5105 (
            .O(N__31319),
            .I(N__31310));
    LocalMux I__5104 (
            .O(N__31316),
            .I(N__31307));
    LocalMux I__5103 (
            .O(N__31313),
            .I(buf_dds1_6));
    Odrv4 I__5102 (
            .O(N__31310),
            .I(buf_dds1_6));
    Odrv4 I__5101 (
            .O(N__31307),
            .I(buf_dds1_6));
    InMux I__5100 (
            .O(N__31300),
            .I(N__31297));
    LocalMux I__5099 (
            .O(N__31297),
            .I(N__31294));
    Span4Mux_v I__5098 (
            .O(N__31294),
            .I(N__31291));
    Span4Mux_h I__5097 (
            .O(N__31291),
            .I(N__31288));
    Span4Mux_h I__5096 (
            .O(N__31288),
            .I(N__31285));
    Odrv4 I__5095 (
            .O(N__31285),
            .I(buf_data_iac_0));
    CascadeMux I__5094 (
            .O(N__31282),
            .I(N__31279));
    InMux I__5093 (
            .O(N__31279),
            .I(N__31276));
    LocalMux I__5092 (
            .O(N__31276),
            .I(N__31272));
    CascadeMux I__5091 (
            .O(N__31275),
            .I(N__31269));
    Span12Mux_v I__5090 (
            .O(N__31272),
            .I(N__31265));
    InMux I__5089 (
            .O(N__31269),
            .I(N__31262));
    InMux I__5088 (
            .O(N__31268),
            .I(N__31259));
    Odrv12 I__5087 (
            .O(N__31265),
            .I(cmd_rdadctmp_21_adj_1527));
    LocalMux I__5086 (
            .O(N__31262),
            .I(cmd_rdadctmp_21_adj_1527));
    LocalMux I__5085 (
            .O(N__31259),
            .I(cmd_rdadctmp_21_adj_1527));
    InMux I__5084 (
            .O(N__31252),
            .I(N__31248));
    InMux I__5083 (
            .O(N__31251),
            .I(N__31245));
    LocalMux I__5082 (
            .O(N__31248),
            .I(N__31240));
    LocalMux I__5081 (
            .O(N__31245),
            .I(N__31240));
    Span4Mux_h I__5080 (
            .O(N__31240),
            .I(N__31237));
    Odrv4 I__5079 (
            .O(N__31237),
            .I(\comm_spi.n15369 ));
    InMux I__5078 (
            .O(N__31234),
            .I(N__31231));
    LocalMux I__5077 (
            .O(N__31231),
            .I(N__31228));
    Span4Mux_v I__5076 (
            .O(N__31228),
            .I(N__31224));
    CascadeMux I__5075 (
            .O(N__31227),
            .I(N__31221));
    Span4Mux_h I__5074 (
            .O(N__31224),
            .I(N__31218));
    InMux I__5073 (
            .O(N__31221),
            .I(N__31215));
    Odrv4 I__5072 (
            .O(N__31218),
            .I(buf_readRTD_13));
    LocalMux I__5071 (
            .O(N__31215),
            .I(buf_readRTD_13));
    InMux I__5070 (
            .O(N__31210),
            .I(N__31207));
    LocalMux I__5069 (
            .O(N__31207),
            .I(N__31204));
    Span4Mux_v I__5068 (
            .O(N__31204),
            .I(N__31201));
    Span4Mux_v I__5067 (
            .O(N__31201),
            .I(N__31198));
    Sp12to4 I__5066 (
            .O(N__31198),
            .I(N__31193));
    InMux I__5065 (
            .O(N__31197),
            .I(N__31190));
    InMux I__5064 (
            .O(N__31196),
            .I(N__31187));
    Span12Mux_h I__5063 (
            .O(N__31193),
            .I(N__31182));
    LocalMux I__5062 (
            .O(N__31190),
            .I(N__31182));
    LocalMux I__5061 (
            .O(N__31187),
            .I(buf_adcdata_vac_21));
    Odrv12 I__5060 (
            .O(N__31182),
            .I(buf_adcdata_vac_21));
    CascadeMux I__5059 (
            .O(N__31177),
            .I(N__31174));
    InMux I__5058 (
            .O(N__31174),
            .I(N__31171));
    LocalMux I__5057 (
            .O(N__31171),
            .I(N__31166));
    InMux I__5056 (
            .O(N__31170),
            .I(N__31163));
    CascadeMux I__5055 (
            .O(N__31169),
            .I(N__31160));
    Span4Mux_h I__5054 (
            .O(N__31166),
            .I(N__31153));
    LocalMux I__5053 (
            .O(N__31163),
            .I(N__31153));
    InMux I__5052 (
            .O(N__31160),
            .I(N__31148));
    InMux I__5051 (
            .O(N__31159),
            .I(N__31148));
    InMux I__5050 (
            .O(N__31158),
            .I(N__31145));
    Span4Mux_h I__5049 (
            .O(N__31153),
            .I(N__31142));
    LocalMux I__5048 (
            .O(N__31148),
            .I(buf_cfgRTD_5));
    LocalMux I__5047 (
            .O(N__31145),
            .I(buf_cfgRTD_5));
    Odrv4 I__5046 (
            .O(N__31142),
            .I(buf_cfgRTD_5));
    CascadeMux I__5045 (
            .O(N__31135),
            .I(n23384_cascade_));
    InMux I__5044 (
            .O(N__31132),
            .I(N__31129));
    LocalMux I__5043 (
            .O(N__31129),
            .I(N__31126));
    Span4Mux_v I__5042 (
            .O(N__31126),
            .I(N__31122));
    InMux I__5041 (
            .O(N__31125),
            .I(N__31119));
    Odrv4 I__5040 (
            .O(N__31122),
            .I(cmd_rdadcbuf_32));
    LocalMux I__5039 (
            .O(N__31119),
            .I(cmd_rdadcbuf_32));
    CascadeMux I__5038 (
            .O(N__31114),
            .I(N__31110));
    CascadeMux I__5037 (
            .O(N__31113),
            .I(N__31107));
    InMux I__5036 (
            .O(N__31110),
            .I(N__31102));
    InMux I__5035 (
            .O(N__31107),
            .I(N__31102));
    LocalMux I__5034 (
            .O(N__31102),
            .I(buf_adcdata_vdc_21));
    InMux I__5033 (
            .O(N__31099),
            .I(N__31096));
    LocalMux I__5032 (
            .O(N__31096),
            .I(N__31092));
    InMux I__5031 (
            .O(N__31095),
            .I(N__31089));
    Odrv12 I__5030 (
            .O(N__31092),
            .I(cmd_rdadcbuf_24));
    LocalMux I__5029 (
            .O(N__31089),
            .I(cmd_rdadcbuf_24));
    CascadeMux I__5028 (
            .O(N__31084),
            .I(N__31069));
    InMux I__5027 (
            .O(N__31083),
            .I(N__31057));
    InMux I__5026 (
            .O(N__31082),
            .I(N__31054));
    InMux I__5025 (
            .O(N__31081),
            .I(N__31037));
    InMux I__5024 (
            .O(N__31080),
            .I(N__31037));
    InMux I__5023 (
            .O(N__31079),
            .I(N__31037));
    InMux I__5022 (
            .O(N__31078),
            .I(N__31037));
    InMux I__5021 (
            .O(N__31077),
            .I(N__31037));
    InMux I__5020 (
            .O(N__31076),
            .I(N__31037));
    InMux I__5019 (
            .O(N__31075),
            .I(N__31037));
    InMux I__5018 (
            .O(N__31074),
            .I(N__31037));
    CascadeMux I__5017 (
            .O(N__31073),
            .I(N__31034));
    InMux I__5016 (
            .O(N__31072),
            .I(N__31017));
    InMux I__5015 (
            .O(N__31069),
            .I(N__31017));
    InMux I__5014 (
            .O(N__31068),
            .I(N__31017));
    InMux I__5013 (
            .O(N__31067),
            .I(N__31017));
    InMux I__5012 (
            .O(N__31066),
            .I(N__31017));
    InMux I__5011 (
            .O(N__31065),
            .I(N__31017));
    InMux I__5010 (
            .O(N__31064),
            .I(N__31017));
    InMux I__5009 (
            .O(N__31063),
            .I(N__31008));
    InMux I__5008 (
            .O(N__31062),
            .I(N__31008));
    InMux I__5007 (
            .O(N__31061),
            .I(N__31008));
    InMux I__5006 (
            .O(N__31060),
            .I(N__31008));
    LocalMux I__5005 (
            .O(N__31057),
            .I(N__31005));
    LocalMux I__5004 (
            .O(N__31054),
            .I(N__31002));
    LocalMux I__5003 (
            .O(N__31037),
            .I(N__30999));
    InMux I__5002 (
            .O(N__31034),
            .I(N__30996));
    InMux I__5001 (
            .O(N__31033),
            .I(N__30991));
    InMux I__5000 (
            .O(N__31032),
            .I(N__30991));
    LocalMux I__4999 (
            .O(N__31017),
            .I(N__30988));
    LocalMux I__4998 (
            .O(N__31008),
            .I(N__30985));
    Span4Mux_h I__4997 (
            .O(N__31005),
            .I(N__30982));
    Span4Mux_v I__4996 (
            .O(N__31002),
            .I(N__30977));
    Span4Mux_h I__4995 (
            .O(N__30999),
            .I(N__30977));
    LocalMux I__4994 (
            .O(N__30996),
            .I(n12352));
    LocalMux I__4993 (
            .O(N__30991),
            .I(n12352));
    Odrv4 I__4992 (
            .O(N__30988),
            .I(n12352));
    Odrv12 I__4991 (
            .O(N__30985),
            .I(n12352));
    Odrv4 I__4990 (
            .O(N__30982),
            .I(n12352));
    Odrv4 I__4989 (
            .O(N__30977),
            .I(n12352));
    InMux I__4988 (
            .O(N__30964),
            .I(N__30961));
    LocalMux I__4987 (
            .O(N__30961),
            .I(N__30958));
    Span4Mux_v I__4986 (
            .O(N__30958),
            .I(N__30954));
    InMux I__4985 (
            .O(N__30957),
            .I(N__30951));
    Odrv4 I__4984 (
            .O(N__30954),
            .I(cmd_rdadcbuf_11));
    LocalMux I__4983 (
            .O(N__30951),
            .I(cmd_rdadcbuf_11));
    InMux I__4982 (
            .O(N__30946),
            .I(N__30942));
    CascadeMux I__4981 (
            .O(N__30945),
            .I(N__30939));
    LocalMux I__4980 (
            .O(N__30942),
            .I(N__30936));
    InMux I__4979 (
            .O(N__30939),
            .I(N__30933));
    Odrv4 I__4978 (
            .O(N__30936),
            .I(buf_adcdata_vdc_12));
    LocalMux I__4977 (
            .O(N__30933),
            .I(buf_adcdata_vdc_12));
    InMux I__4976 (
            .O(N__30928),
            .I(N__30925));
    LocalMux I__4975 (
            .O(N__30925),
            .I(N__30922));
    Span4Mux_h I__4974 (
            .O(N__30922),
            .I(N__30919));
    Span4Mux_h I__4973 (
            .O(N__30919),
            .I(N__30915));
    InMux I__4972 (
            .O(N__30918),
            .I(N__30912));
    Span4Mux_h I__4971 (
            .O(N__30915),
            .I(N__30908));
    LocalMux I__4970 (
            .O(N__30912),
            .I(N__30905));
    InMux I__4969 (
            .O(N__30911),
            .I(N__30902));
    Span4Mux_v I__4968 (
            .O(N__30908),
            .I(N__30899));
    Span4Mux_h I__4967 (
            .O(N__30905),
            .I(N__30896));
    LocalMux I__4966 (
            .O(N__30902),
            .I(buf_adcdata_vac_12));
    Odrv4 I__4965 (
            .O(N__30899),
            .I(buf_adcdata_vac_12));
    Odrv4 I__4964 (
            .O(N__30896),
            .I(buf_adcdata_vac_12));
    InMux I__4963 (
            .O(N__30889),
            .I(N__30886));
    LocalMux I__4962 (
            .O(N__30886),
            .I(N__30883));
    Span4Mux_v I__4961 (
            .O(N__30883),
            .I(N__30879));
    CascadeMux I__4960 (
            .O(N__30882),
            .I(N__30876));
    Span4Mux_h I__4959 (
            .O(N__30879),
            .I(N__30873));
    InMux I__4958 (
            .O(N__30876),
            .I(N__30870));
    Odrv4 I__4957 (
            .O(N__30873),
            .I(buf_readRTD_4));
    LocalMux I__4956 (
            .O(N__30870),
            .I(buf_readRTD_4));
    CascadeMux I__4955 (
            .O(N__30865),
            .I(n19_adj_1734_cascade_));
    InMux I__4954 (
            .O(N__30862),
            .I(N__30859));
    LocalMux I__4953 (
            .O(N__30859),
            .I(N__30856));
    Span4Mux_v I__4952 (
            .O(N__30856),
            .I(N__30853));
    Odrv4 I__4951 (
            .O(N__30853),
            .I(\ADC_VDC.n21991 ));
    CascadeMux I__4950 (
            .O(N__30850),
            .I(\ADC_VDC.n22075_cascade_ ));
    InMux I__4949 (
            .O(N__30847),
            .I(N__30844));
    LocalMux I__4948 (
            .O(N__30844),
            .I(\ADC_VDC.n44_adj_1487 ));
    CEMux I__4947 (
            .O(N__30841),
            .I(N__30838));
    LocalMux I__4946 (
            .O(N__30838),
            .I(N__30835));
    Odrv12 I__4945 (
            .O(N__30835),
            .I(\ADC_VDC.n39_adj_1488 ));
    InMux I__4944 (
            .O(N__30832),
            .I(N__30829));
    LocalMux I__4943 (
            .O(N__30829),
            .I(\ADC_VDC.n6_adj_1485 ));
    CascadeMux I__4942 (
            .O(N__30826),
            .I(\ADC_VDC.n21859_cascade_ ));
    CascadeMux I__4941 (
            .O(N__30823),
            .I(\ADC_VDC.n22628_cascade_ ));
    InMux I__4940 (
            .O(N__30820),
            .I(N__30816));
    InMux I__4939 (
            .O(N__30819),
            .I(N__30813));
    LocalMux I__4938 (
            .O(N__30816),
            .I(\ADC_VDC.n21859 ));
    LocalMux I__4937 (
            .O(N__30813),
            .I(\ADC_VDC.n21859 ));
    InMux I__4936 (
            .O(N__30808),
            .I(N__30805));
    LocalMux I__4935 (
            .O(N__30805),
            .I(\ADC_VDC.n22625 ));
    InMux I__4934 (
            .O(N__30802),
            .I(N__30799));
    LocalMux I__4933 (
            .O(N__30799),
            .I(\ADC_VDC.n6 ));
    InMux I__4932 (
            .O(N__30796),
            .I(N__30791));
    CascadeMux I__4931 (
            .O(N__30795),
            .I(N__30788));
    CascadeMux I__4930 (
            .O(N__30794),
            .I(N__30785));
    LocalMux I__4929 (
            .O(N__30791),
            .I(N__30782));
    InMux I__4928 (
            .O(N__30788),
            .I(N__30779));
    InMux I__4927 (
            .O(N__30785),
            .I(N__30776));
    Span4Mux_h I__4926 (
            .O(N__30782),
            .I(N__30773));
    LocalMux I__4925 (
            .O(N__30779),
            .I(N__30768));
    LocalMux I__4924 (
            .O(N__30776),
            .I(N__30768));
    Odrv4 I__4923 (
            .O(N__30773),
            .I(cmd_rdadctmp_22_adj_1552));
    Odrv4 I__4922 (
            .O(N__30768),
            .I(cmd_rdadctmp_22_adj_1552));
    CascadeMux I__4921 (
            .O(N__30763),
            .I(\ADC_VDC.n11183_cascade_ ));
    CascadeMux I__4920 (
            .O(N__30760),
            .I(N__30757));
    InMux I__4919 (
            .O(N__30757),
            .I(N__30754));
    LocalMux I__4918 (
            .O(N__30754),
            .I(N__30750));
    InMux I__4917 (
            .O(N__30753),
            .I(N__30747));
    Span4Mux_h I__4916 (
            .O(N__30750),
            .I(N__30744));
    LocalMux I__4915 (
            .O(N__30747),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    Odrv4 I__4914 (
            .O(N__30744),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    CEMux I__4913 (
            .O(N__30739),
            .I(N__30736));
    LocalMux I__4912 (
            .O(N__30736),
            .I(N__30733));
    Span4Mux_v I__4911 (
            .O(N__30733),
            .I(N__30730));
    Span4Mux_h I__4910 (
            .O(N__30730),
            .I(N__30727));
    Odrv4 I__4909 (
            .O(N__30727),
            .I(\ADC_VDC.n13957 ));
    SRMux I__4908 (
            .O(N__30724),
            .I(N__30721));
    LocalMux I__4907 (
            .O(N__30721),
            .I(N__30718));
    Odrv4 I__4906 (
            .O(N__30718),
            .I(\ADC_VDC.n21707 ));
    CascadeMux I__4905 (
            .O(N__30715),
            .I(\ADC_VDC.n17_cascade_ ));
    InMux I__4904 (
            .O(N__30712),
            .I(N__30709));
    LocalMux I__4903 (
            .O(N__30709),
            .I(N__30706));
    Odrv4 I__4902 (
            .O(N__30706),
            .I(\ADC_VDC.n22055 ));
    CascadeMux I__4901 (
            .O(N__30703),
            .I(\ADC_VDC.n27_cascade_ ));
    InMux I__4900 (
            .O(N__30700),
            .I(N__30697));
    LocalMux I__4899 (
            .O(N__30697),
            .I(\ADC_VDC.n10 ));
    CEMux I__4898 (
            .O(N__30694),
            .I(N__30691));
    LocalMux I__4897 (
            .O(N__30691),
            .I(N__30688));
    Odrv4 I__4896 (
            .O(N__30688),
            .I(\ADC_VDC.n21869 ));
    InMux I__4895 (
            .O(N__30685),
            .I(N__30682));
    LocalMux I__4894 (
            .O(N__30682),
            .I(\ADC_VDC.n11923 ));
    CascadeMux I__4893 (
            .O(N__30679),
            .I(\ADC_VDC.n11923_cascade_ ));
    CascadeMux I__4892 (
            .O(N__30676),
            .I(\ADC_VDC.n20869_cascade_ ));
    InMux I__4891 (
            .O(N__30673),
            .I(N__30670));
    LocalMux I__4890 (
            .O(N__30670),
            .I(N__30667));
    Span4Mux_h I__4889 (
            .O(N__30667),
            .I(N__30664));
    Odrv4 I__4888 (
            .O(N__30664),
            .I(\ADC_VDC.n8031 ));
    CascadeMux I__4887 (
            .O(N__30661),
            .I(N__30658));
    InMux I__4886 (
            .O(N__30658),
            .I(N__30655));
    LocalMux I__4885 (
            .O(N__30655),
            .I(N__30652));
    Odrv12 I__4884 (
            .O(N__30652),
            .I(\ADC_VDC.n23531 ));
    InMux I__4883 (
            .O(N__30649),
            .I(N__30646));
    LocalMux I__4882 (
            .O(N__30646),
            .I(\ADC_VDC.n20869 ));
    InMux I__4881 (
            .O(N__30643),
            .I(N__30640));
    LocalMux I__4880 (
            .O(N__30640),
            .I(N__30635));
    InMux I__4879 (
            .O(N__30639),
            .I(N__30632));
    InMux I__4878 (
            .O(N__30638),
            .I(N__30629));
    Span4Mux_v I__4877 (
            .O(N__30635),
            .I(N__30626));
    LocalMux I__4876 (
            .O(N__30632),
            .I(buf_dds1_10));
    LocalMux I__4875 (
            .O(N__30629),
            .I(buf_dds1_10));
    Odrv4 I__4874 (
            .O(N__30626),
            .I(buf_dds1_10));
    CascadeMux I__4873 (
            .O(N__30619),
            .I(N__30616));
    InMux I__4872 (
            .O(N__30616),
            .I(N__30613));
    LocalMux I__4871 (
            .O(N__30613),
            .I(n22160));
    InMux I__4870 (
            .O(N__30610),
            .I(N__30607));
    LocalMux I__4869 (
            .O(N__30607),
            .I(N__30604));
    Span4Mux_v I__4868 (
            .O(N__30604),
            .I(N__30600));
    CascadeMux I__4867 (
            .O(N__30603),
            .I(N__30596));
    Span4Mux_v I__4866 (
            .O(N__30600),
            .I(N__30593));
    InMux I__4865 (
            .O(N__30599),
            .I(N__30590));
    InMux I__4864 (
            .O(N__30596),
            .I(N__30587));
    Sp12to4 I__4863 (
            .O(N__30593),
            .I(N__30584));
    LocalMux I__4862 (
            .O(N__30590),
            .I(N__30581));
    LocalMux I__4861 (
            .O(N__30587),
            .I(buf_adcdata_iac_18));
    Odrv12 I__4860 (
            .O(N__30584),
            .I(buf_adcdata_iac_18));
    Odrv4 I__4859 (
            .O(N__30581),
            .I(buf_adcdata_iac_18));
    IoInMux I__4858 (
            .O(N__30574),
            .I(N__30571));
    LocalMux I__4857 (
            .O(N__30571),
            .I(N__30568));
    Span4Mux_s2_v I__4856 (
            .O(N__30568),
            .I(N__30565));
    Span4Mux_v I__4855 (
            .O(N__30565),
            .I(N__30561));
    InMux I__4854 (
            .O(N__30564),
            .I(N__30557));
    Span4Mux_v I__4853 (
            .O(N__30561),
            .I(N__30554));
    InMux I__4852 (
            .O(N__30560),
            .I(N__30551));
    LocalMux I__4851 (
            .O(N__30557),
            .I(N__30548));
    Odrv4 I__4850 (
            .O(N__30554),
            .I(IAC_FLT0));
    LocalMux I__4849 (
            .O(N__30551),
            .I(IAC_FLT0));
    Odrv4 I__4848 (
            .O(N__30548),
            .I(IAC_FLT0));
    InMux I__4847 (
            .O(N__30541),
            .I(N__30538));
    LocalMux I__4846 (
            .O(N__30538),
            .I(n22161));
    InMux I__4845 (
            .O(N__30535),
            .I(N__30532));
    LocalMux I__4844 (
            .O(N__30532),
            .I(N__30528));
    InMux I__4843 (
            .O(N__30531),
            .I(N__30525));
    Odrv12 I__4842 (
            .O(N__30528),
            .I(\ADC_VDC.adc_state_3_N_1316_1 ));
    LocalMux I__4841 (
            .O(N__30525),
            .I(\ADC_VDC.adc_state_3_N_1316_1 ));
    CascadeMux I__4840 (
            .O(N__30520),
            .I(\ADC_VDC.n22404_cascade_ ));
    InMux I__4839 (
            .O(N__30517),
            .I(N__30514));
    LocalMux I__4838 (
            .O(N__30514),
            .I(\ADC_VDC.n17 ));
    CascadeMux I__4837 (
            .O(N__30511),
            .I(N__30507));
    InMux I__4836 (
            .O(N__30510),
            .I(N__30503));
    InMux I__4835 (
            .O(N__30507),
            .I(N__30500));
    InMux I__4834 (
            .O(N__30506),
            .I(N__30497));
    LocalMux I__4833 (
            .O(N__30503),
            .I(cmd_rdadctmp_24));
    LocalMux I__4832 (
            .O(N__30500),
            .I(cmd_rdadctmp_24));
    LocalMux I__4831 (
            .O(N__30497),
            .I(cmd_rdadctmp_24));
    CascadeMux I__4830 (
            .O(N__30490),
            .I(N__30487));
    InMux I__4829 (
            .O(N__30487),
            .I(N__30484));
    LocalMux I__4828 (
            .O(N__30484),
            .I(N__30481));
    Span4Mux_h I__4827 (
            .O(N__30481),
            .I(N__30477));
    InMux I__4826 (
            .O(N__30480),
            .I(N__30474));
    Odrv4 I__4825 (
            .O(N__30477),
            .I(cmd_rdadctmp_5));
    LocalMux I__4824 (
            .O(N__30474),
            .I(cmd_rdadctmp_5));
    InMux I__4823 (
            .O(N__30469),
            .I(N__30466));
    LocalMux I__4822 (
            .O(N__30466),
            .I(N__30463));
    Odrv12 I__4821 (
            .O(N__30463),
            .I(n23468));
    CascadeMux I__4820 (
            .O(N__30460),
            .I(N__30457));
    InMux I__4819 (
            .O(N__30457),
            .I(N__30453));
    InMux I__4818 (
            .O(N__30456),
            .I(N__30449));
    LocalMux I__4817 (
            .O(N__30453),
            .I(N__30446));
    InMux I__4816 (
            .O(N__30452),
            .I(N__30443));
    LocalMux I__4815 (
            .O(N__30449),
            .I(cmd_rdadctmp_25));
    Odrv4 I__4814 (
            .O(N__30446),
            .I(cmd_rdadctmp_25));
    LocalMux I__4813 (
            .O(N__30443),
            .I(cmd_rdadctmp_25));
    InMux I__4812 (
            .O(N__30436),
            .I(N__30429));
    InMux I__4811 (
            .O(N__30435),
            .I(N__30426));
    CascadeMux I__4810 (
            .O(N__30434),
            .I(N__30419));
    CascadeMux I__4809 (
            .O(N__30433),
            .I(N__30415));
    CascadeMux I__4808 (
            .O(N__30432),
            .I(N__30412));
    LocalMux I__4807 (
            .O(N__30429),
            .I(N__30405));
    LocalMux I__4806 (
            .O(N__30426),
            .I(N__30405));
    InMux I__4805 (
            .O(N__30425),
            .I(N__30402));
    InMux I__4804 (
            .O(N__30424),
            .I(N__30395));
    InMux I__4803 (
            .O(N__30423),
            .I(N__30395));
    InMux I__4802 (
            .O(N__30422),
            .I(N__30395));
    InMux I__4801 (
            .O(N__30419),
            .I(N__30382));
    InMux I__4800 (
            .O(N__30418),
            .I(N__30382));
    InMux I__4799 (
            .O(N__30415),
            .I(N__30382));
    InMux I__4798 (
            .O(N__30412),
            .I(N__30382));
    InMux I__4797 (
            .O(N__30411),
            .I(N__30382));
    InMux I__4796 (
            .O(N__30410),
            .I(N__30382));
    Odrv12 I__4795 (
            .O(N__30405),
            .I(DTRIG_N_1182));
    LocalMux I__4794 (
            .O(N__30402),
            .I(DTRIG_N_1182));
    LocalMux I__4793 (
            .O(N__30395),
            .I(DTRIG_N_1182));
    LocalMux I__4792 (
            .O(N__30382),
            .I(DTRIG_N_1182));
    CascadeMux I__4791 (
            .O(N__30373),
            .I(N__30368));
    CascadeMux I__4790 (
            .O(N__30372),
            .I(N__30362));
    InMux I__4789 (
            .O(N__30371),
            .I(N__30359));
    InMux I__4788 (
            .O(N__30368),
            .I(N__30356));
    InMux I__4787 (
            .O(N__30367),
            .I(N__30353));
    InMux I__4786 (
            .O(N__30366),
            .I(N__30346));
    InMux I__4785 (
            .O(N__30365),
            .I(N__30346));
    InMux I__4784 (
            .O(N__30362),
            .I(N__30346));
    LocalMux I__4783 (
            .O(N__30359),
            .I(N__30337));
    LocalMux I__4782 (
            .O(N__30356),
            .I(N__30334));
    LocalMux I__4781 (
            .O(N__30353),
            .I(N__30331));
    LocalMux I__4780 (
            .O(N__30346),
            .I(N__30328));
    InMux I__4779 (
            .O(N__30345),
            .I(N__30315));
    InMux I__4778 (
            .O(N__30344),
            .I(N__30315));
    InMux I__4777 (
            .O(N__30343),
            .I(N__30315));
    InMux I__4776 (
            .O(N__30342),
            .I(N__30315));
    InMux I__4775 (
            .O(N__30341),
            .I(N__30315));
    InMux I__4774 (
            .O(N__30340),
            .I(N__30315));
    Odrv4 I__4773 (
            .O(N__30337),
            .I(adc_state_1));
    Odrv12 I__4772 (
            .O(N__30334),
            .I(adc_state_1));
    Odrv4 I__4771 (
            .O(N__30331),
            .I(adc_state_1));
    Odrv4 I__4770 (
            .O(N__30328),
            .I(adc_state_1));
    LocalMux I__4769 (
            .O(N__30315),
            .I(adc_state_1));
    CascadeMux I__4768 (
            .O(N__30304),
            .I(N__30300));
    CascadeMux I__4767 (
            .O(N__30303),
            .I(N__30297));
    InMux I__4766 (
            .O(N__30300),
            .I(N__30294));
    InMux I__4765 (
            .O(N__30297),
            .I(N__30291));
    LocalMux I__4764 (
            .O(N__30294),
            .I(N__30288));
    LocalMux I__4763 (
            .O(N__30291),
            .I(N__30284));
    Span4Mux_v I__4762 (
            .O(N__30288),
            .I(N__30281));
    InMux I__4761 (
            .O(N__30287),
            .I(N__30278));
    Odrv12 I__4760 (
            .O(N__30284),
            .I(cmd_rdadctmp_27));
    Odrv4 I__4759 (
            .O(N__30281),
            .I(cmd_rdadctmp_27));
    LocalMux I__4758 (
            .O(N__30278),
            .I(cmd_rdadctmp_27));
    InMux I__4757 (
            .O(N__30271),
            .I(N__30268));
    LocalMux I__4756 (
            .O(N__30268),
            .I(N__30264));
    CascadeMux I__4755 (
            .O(N__30267),
            .I(N__30260));
    Span12Mux_v I__4754 (
            .O(N__30264),
            .I(N__30257));
    CascadeMux I__4753 (
            .O(N__30263),
            .I(N__30254));
    InMux I__4752 (
            .O(N__30260),
            .I(N__30251));
    Span12Mux_h I__4751 (
            .O(N__30257),
            .I(N__30248));
    InMux I__4750 (
            .O(N__30254),
            .I(N__30245));
    LocalMux I__4749 (
            .O(N__30251),
            .I(buf_adcdata_iac_17));
    Odrv12 I__4748 (
            .O(N__30248),
            .I(buf_adcdata_iac_17));
    LocalMux I__4747 (
            .O(N__30245),
            .I(buf_adcdata_iac_17));
    CascadeMux I__4746 (
            .O(N__30238),
            .I(N__30235));
    CascadeBuf I__4745 (
            .O(N__30235),
            .I(N__30232));
    CascadeMux I__4744 (
            .O(N__30232),
            .I(N__30229));
    CascadeBuf I__4743 (
            .O(N__30229),
            .I(N__30226));
    CascadeMux I__4742 (
            .O(N__30226),
            .I(N__30223));
    CascadeBuf I__4741 (
            .O(N__30223),
            .I(N__30220));
    CascadeMux I__4740 (
            .O(N__30220),
            .I(N__30217));
    CascadeBuf I__4739 (
            .O(N__30217),
            .I(N__30214));
    CascadeMux I__4738 (
            .O(N__30214),
            .I(N__30211));
    CascadeBuf I__4737 (
            .O(N__30211),
            .I(N__30208));
    CascadeMux I__4736 (
            .O(N__30208),
            .I(N__30205));
    CascadeBuf I__4735 (
            .O(N__30205),
            .I(N__30202));
    CascadeMux I__4734 (
            .O(N__30202),
            .I(N__30199));
    CascadeBuf I__4733 (
            .O(N__30199),
            .I(N__30196));
    CascadeMux I__4732 (
            .O(N__30196),
            .I(N__30193));
    CascadeBuf I__4731 (
            .O(N__30193),
            .I(N__30190));
    CascadeMux I__4730 (
            .O(N__30190),
            .I(N__30186));
    CascadeMux I__4729 (
            .O(N__30189),
            .I(N__30183));
    CascadeBuf I__4728 (
            .O(N__30186),
            .I(N__30180));
    CascadeBuf I__4727 (
            .O(N__30183),
            .I(N__30177));
    CascadeMux I__4726 (
            .O(N__30180),
            .I(N__30174));
    CascadeMux I__4725 (
            .O(N__30177),
            .I(N__30171));
    InMux I__4724 (
            .O(N__30174),
            .I(N__30168));
    InMux I__4723 (
            .O(N__30171),
            .I(N__30165));
    LocalMux I__4722 (
            .O(N__30168),
            .I(N__30162));
    LocalMux I__4721 (
            .O(N__30165),
            .I(N__30158));
    Span12Mux_s7_h I__4720 (
            .O(N__30162),
            .I(N__30155));
    InMux I__4719 (
            .O(N__30161),
            .I(N__30152));
    Span12Mux_h I__4718 (
            .O(N__30158),
            .I(N__30147));
    Span12Mux_h I__4717 (
            .O(N__30155),
            .I(N__30147));
    LocalMux I__4716 (
            .O(N__30152),
            .I(data_count_6));
    Odrv12 I__4715 (
            .O(N__30147),
            .I(data_count_6));
    InMux I__4714 (
            .O(N__30142),
            .I(n20618));
    CascadeMux I__4713 (
            .O(N__30139),
            .I(N__30136));
    CascadeBuf I__4712 (
            .O(N__30136),
            .I(N__30133));
    CascadeMux I__4711 (
            .O(N__30133),
            .I(N__30130));
    CascadeBuf I__4710 (
            .O(N__30130),
            .I(N__30127));
    CascadeMux I__4709 (
            .O(N__30127),
            .I(N__30124));
    CascadeBuf I__4708 (
            .O(N__30124),
            .I(N__30121));
    CascadeMux I__4707 (
            .O(N__30121),
            .I(N__30118));
    CascadeBuf I__4706 (
            .O(N__30118),
            .I(N__30115));
    CascadeMux I__4705 (
            .O(N__30115),
            .I(N__30112));
    CascadeBuf I__4704 (
            .O(N__30112),
            .I(N__30109));
    CascadeMux I__4703 (
            .O(N__30109),
            .I(N__30106));
    CascadeBuf I__4702 (
            .O(N__30106),
            .I(N__30103));
    CascadeMux I__4701 (
            .O(N__30103),
            .I(N__30100));
    CascadeBuf I__4700 (
            .O(N__30100),
            .I(N__30097));
    CascadeMux I__4699 (
            .O(N__30097),
            .I(N__30094));
    CascadeBuf I__4698 (
            .O(N__30094),
            .I(N__30090));
    CascadeMux I__4697 (
            .O(N__30093),
            .I(N__30087));
    CascadeMux I__4696 (
            .O(N__30090),
            .I(N__30084));
    CascadeBuf I__4695 (
            .O(N__30087),
            .I(N__30081));
    CascadeBuf I__4694 (
            .O(N__30084),
            .I(N__30078));
    CascadeMux I__4693 (
            .O(N__30081),
            .I(N__30075));
    CascadeMux I__4692 (
            .O(N__30078),
            .I(N__30072));
    InMux I__4691 (
            .O(N__30075),
            .I(N__30069));
    InMux I__4690 (
            .O(N__30072),
            .I(N__30066));
    LocalMux I__4689 (
            .O(N__30069),
            .I(N__30063));
    LocalMux I__4688 (
            .O(N__30066),
            .I(N__30060));
    Span4Mux_h I__4687 (
            .O(N__30063),
            .I(N__30057));
    Span4Mux_v I__4686 (
            .O(N__30060),
            .I(N__30054));
    Span4Mux_h I__4685 (
            .O(N__30057),
            .I(N__30050));
    Sp12to4 I__4684 (
            .O(N__30054),
            .I(N__30047));
    InMux I__4683 (
            .O(N__30053),
            .I(N__30044));
    Sp12to4 I__4682 (
            .O(N__30050),
            .I(N__30039));
    Span12Mux_h I__4681 (
            .O(N__30047),
            .I(N__30039));
    LocalMux I__4680 (
            .O(N__30044),
            .I(data_count_7));
    Odrv12 I__4679 (
            .O(N__30039),
            .I(data_count_7));
    InMux I__4678 (
            .O(N__30034),
            .I(n20619));
    CascadeMux I__4677 (
            .O(N__30031),
            .I(N__30028));
    CascadeBuf I__4676 (
            .O(N__30028),
            .I(N__30025));
    CascadeMux I__4675 (
            .O(N__30025),
            .I(N__30022));
    CascadeBuf I__4674 (
            .O(N__30022),
            .I(N__30019));
    CascadeMux I__4673 (
            .O(N__30019),
            .I(N__30016));
    CascadeBuf I__4672 (
            .O(N__30016),
            .I(N__30013));
    CascadeMux I__4671 (
            .O(N__30013),
            .I(N__30010));
    CascadeBuf I__4670 (
            .O(N__30010),
            .I(N__30007));
    CascadeMux I__4669 (
            .O(N__30007),
            .I(N__30004));
    CascadeBuf I__4668 (
            .O(N__30004),
            .I(N__30001));
    CascadeMux I__4667 (
            .O(N__30001),
            .I(N__29998));
    CascadeBuf I__4666 (
            .O(N__29998),
            .I(N__29995));
    CascadeMux I__4665 (
            .O(N__29995),
            .I(N__29992));
    CascadeBuf I__4664 (
            .O(N__29992),
            .I(N__29989));
    CascadeMux I__4663 (
            .O(N__29989),
            .I(N__29986));
    CascadeBuf I__4662 (
            .O(N__29986),
            .I(N__29982));
    CascadeMux I__4661 (
            .O(N__29985),
            .I(N__29979));
    CascadeMux I__4660 (
            .O(N__29982),
            .I(N__29976));
    CascadeBuf I__4659 (
            .O(N__29979),
            .I(N__29973));
    CascadeBuf I__4658 (
            .O(N__29976),
            .I(N__29970));
    CascadeMux I__4657 (
            .O(N__29973),
            .I(N__29967));
    CascadeMux I__4656 (
            .O(N__29970),
            .I(N__29964));
    InMux I__4655 (
            .O(N__29967),
            .I(N__29961));
    InMux I__4654 (
            .O(N__29964),
            .I(N__29958));
    LocalMux I__4653 (
            .O(N__29961),
            .I(N__29955));
    LocalMux I__4652 (
            .O(N__29958),
            .I(N__29952));
    Span4Mux_v I__4651 (
            .O(N__29955),
            .I(N__29948));
    Span12Mux_v I__4650 (
            .O(N__29952),
            .I(N__29945));
    InMux I__4649 (
            .O(N__29951),
            .I(N__29942));
    Span4Mux_h I__4648 (
            .O(N__29948),
            .I(N__29939));
    Span12Mux_h I__4647 (
            .O(N__29945),
            .I(N__29936));
    LocalMux I__4646 (
            .O(N__29942),
            .I(data_count_8));
    Odrv4 I__4645 (
            .O(N__29939),
            .I(data_count_8));
    Odrv12 I__4644 (
            .O(N__29936),
            .I(data_count_8));
    InMux I__4643 (
            .O(N__29929),
            .I(bfn_9_15_0_));
    InMux I__4642 (
            .O(N__29926),
            .I(n20621));
    CascadeMux I__4641 (
            .O(N__29923),
            .I(N__29920));
    CascadeBuf I__4640 (
            .O(N__29920),
            .I(N__29917));
    CascadeMux I__4639 (
            .O(N__29917),
            .I(N__29914));
    CascadeBuf I__4638 (
            .O(N__29914),
            .I(N__29911));
    CascadeMux I__4637 (
            .O(N__29911),
            .I(N__29908));
    CascadeBuf I__4636 (
            .O(N__29908),
            .I(N__29905));
    CascadeMux I__4635 (
            .O(N__29905),
            .I(N__29902));
    CascadeBuf I__4634 (
            .O(N__29902),
            .I(N__29899));
    CascadeMux I__4633 (
            .O(N__29899),
            .I(N__29896));
    CascadeBuf I__4632 (
            .O(N__29896),
            .I(N__29893));
    CascadeMux I__4631 (
            .O(N__29893),
            .I(N__29890));
    CascadeBuf I__4630 (
            .O(N__29890),
            .I(N__29887));
    CascadeMux I__4629 (
            .O(N__29887),
            .I(N__29884));
    CascadeBuf I__4628 (
            .O(N__29884),
            .I(N__29881));
    CascadeMux I__4627 (
            .O(N__29881),
            .I(N__29878));
    CascadeBuf I__4626 (
            .O(N__29878),
            .I(N__29875));
    CascadeMux I__4625 (
            .O(N__29875),
            .I(N__29871));
    CascadeMux I__4624 (
            .O(N__29874),
            .I(N__29868));
    CascadeBuf I__4623 (
            .O(N__29871),
            .I(N__29865));
    CascadeBuf I__4622 (
            .O(N__29868),
            .I(N__29862));
    CascadeMux I__4621 (
            .O(N__29865),
            .I(N__29859));
    CascadeMux I__4620 (
            .O(N__29862),
            .I(N__29856));
    InMux I__4619 (
            .O(N__29859),
            .I(N__29853));
    InMux I__4618 (
            .O(N__29856),
            .I(N__29850));
    LocalMux I__4617 (
            .O(N__29853),
            .I(N__29847));
    LocalMux I__4616 (
            .O(N__29850),
            .I(N__29843));
    Span12Mux_v I__4615 (
            .O(N__29847),
            .I(N__29840));
    InMux I__4614 (
            .O(N__29846),
            .I(N__29837));
    Span12Mux_v I__4613 (
            .O(N__29843),
            .I(N__29834));
    Span12Mux_h I__4612 (
            .O(N__29840),
            .I(N__29831));
    LocalMux I__4611 (
            .O(N__29837),
            .I(data_count_9));
    Odrv12 I__4610 (
            .O(N__29834),
            .I(data_count_9));
    Odrv12 I__4609 (
            .O(N__29831),
            .I(data_count_9));
    InMux I__4608 (
            .O(N__29824),
            .I(N__29821));
    LocalMux I__4607 (
            .O(N__29821),
            .I(N__29818));
    Odrv4 I__4606 (
            .O(N__29818),
            .I(n11983));
    CascadeMux I__4605 (
            .O(N__29815),
            .I(n24_adj_1598_cascade_));
    CascadeMux I__4604 (
            .O(N__29812),
            .I(n24_adj_1506_cascade_));
    IoInMux I__4603 (
            .O(N__29809),
            .I(N__29806));
    LocalMux I__4602 (
            .O(N__29806),
            .I(N__29803));
    Span4Mux_s2_v I__4601 (
            .O(N__29803),
            .I(N__29800));
    Span4Mux_h I__4600 (
            .O(N__29800),
            .I(N__29796));
    InMux I__4599 (
            .O(N__29799),
            .I(N__29793));
    Span4Mux_v I__4598 (
            .O(N__29796),
            .I(N__29790));
    LocalMux I__4597 (
            .O(N__29793),
            .I(N__29786));
    Span4Mux_v I__4596 (
            .O(N__29790),
            .I(N__29783));
    InMux I__4595 (
            .O(N__29789),
            .I(N__29780));
    Span4Mux_h I__4594 (
            .O(N__29786),
            .I(N__29777));
    Odrv4 I__4593 (
            .O(N__29783),
            .I(IAC_FLT1));
    LocalMux I__4592 (
            .O(N__29780),
            .I(IAC_FLT1));
    Odrv4 I__4591 (
            .O(N__29777),
            .I(IAC_FLT1));
    InMux I__4590 (
            .O(N__29770),
            .I(N__29767));
    LocalMux I__4589 (
            .O(N__29767),
            .I(n11982));
    CascadeMux I__4588 (
            .O(N__29764),
            .I(N__29761));
    InMux I__4587 (
            .O(N__29761),
            .I(N__29758));
    LocalMux I__4586 (
            .O(N__29758),
            .I(N__29754));
    CascadeMux I__4585 (
            .O(N__29757),
            .I(N__29751));
    Span4Mux_v I__4584 (
            .O(N__29754),
            .I(N__29747));
    InMux I__4583 (
            .O(N__29751),
            .I(N__29744));
    InMux I__4582 (
            .O(N__29750),
            .I(N__29741));
    Odrv4 I__4581 (
            .O(N__29747),
            .I(cmd_rdadctmp_18));
    LocalMux I__4580 (
            .O(N__29744),
            .I(cmd_rdadctmp_18));
    LocalMux I__4579 (
            .O(N__29741),
            .I(cmd_rdadctmp_18));
    InMux I__4578 (
            .O(N__29734),
            .I(N__29729));
    InMux I__4577 (
            .O(N__29733),
            .I(N__29726));
    InMux I__4576 (
            .O(N__29732),
            .I(N__29723));
    LocalMux I__4575 (
            .O(N__29729),
            .I(N__29720));
    LocalMux I__4574 (
            .O(N__29726),
            .I(N__29717));
    LocalMux I__4573 (
            .O(N__29723),
            .I(buf_dds1_11));
    Odrv4 I__4572 (
            .O(N__29720),
            .I(buf_dds1_11));
    Odrv4 I__4571 (
            .O(N__29717),
            .I(buf_dds1_11));
    CascadeMux I__4570 (
            .O(N__29710),
            .I(N__29707));
    CascadeBuf I__4569 (
            .O(N__29707),
            .I(N__29704));
    CascadeMux I__4568 (
            .O(N__29704),
            .I(N__29701));
    CascadeBuf I__4567 (
            .O(N__29701),
            .I(N__29698));
    CascadeMux I__4566 (
            .O(N__29698),
            .I(N__29695));
    CascadeBuf I__4565 (
            .O(N__29695),
            .I(N__29692));
    CascadeMux I__4564 (
            .O(N__29692),
            .I(N__29689));
    CascadeBuf I__4563 (
            .O(N__29689),
            .I(N__29686));
    CascadeMux I__4562 (
            .O(N__29686),
            .I(N__29683));
    CascadeBuf I__4561 (
            .O(N__29683),
            .I(N__29680));
    CascadeMux I__4560 (
            .O(N__29680),
            .I(N__29677));
    CascadeBuf I__4559 (
            .O(N__29677),
            .I(N__29674));
    CascadeMux I__4558 (
            .O(N__29674),
            .I(N__29671));
    CascadeBuf I__4557 (
            .O(N__29671),
            .I(N__29668));
    CascadeMux I__4556 (
            .O(N__29668),
            .I(N__29665));
    CascadeBuf I__4555 (
            .O(N__29665),
            .I(N__29661));
    CascadeMux I__4554 (
            .O(N__29664),
            .I(N__29658));
    CascadeMux I__4553 (
            .O(N__29661),
            .I(N__29655));
    CascadeBuf I__4552 (
            .O(N__29658),
            .I(N__29652));
    CascadeBuf I__4551 (
            .O(N__29655),
            .I(N__29649));
    CascadeMux I__4550 (
            .O(N__29652),
            .I(N__29646));
    CascadeMux I__4549 (
            .O(N__29649),
            .I(N__29643));
    InMux I__4548 (
            .O(N__29646),
            .I(N__29640));
    InMux I__4547 (
            .O(N__29643),
            .I(N__29637));
    LocalMux I__4546 (
            .O(N__29640),
            .I(N__29634));
    LocalMux I__4545 (
            .O(N__29637),
            .I(N__29631));
    Span4Mux_v I__4544 (
            .O(N__29634),
            .I(N__29627));
    Span12Mux_v I__4543 (
            .O(N__29631),
            .I(N__29624));
    InMux I__4542 (
            .O(N__29630),
            .I(N__29621));
    Span4Mux_h I__4541 (
            .O(N__29627),
            .I(N__29618));
    Span12Mux_h I__4540 (
            .O(N__29624),
            .I(N__29615));
    LocalMux I__4539 (
            .O(N__29621),
            .I(data_count_0));
    Odrv4 I__4538 (
            .O(N__29618),
            .I(data_count_0));
    Odrv12 I__4537 (
            .O(N__29615),
            .I(data_count_0));
    CascadeMux I__4536 (
            .O(N__29608),
            .I(N__29605));
    CascadeBuf I__4535 (
            .O(N__29605),
            .I(N__29602));
    CascadeMux I__4534 (
            .O(N__29602),
            .I(N__29599));
    CascadeBuf I__4533 (
            .O(N__29599),
            .I(N__29596));
    CascadeMux I__4532 (
            .O(N__29596),
            .I(N__29593));
    CascadeBuf I__4531 (
            .O(N__29593),
            .I(N__29590));
    CascadeMux I__4530 (
            .O(N__29590),
            .I(N__29587));
    CascadeBuf I__4529 (
            .O(N__29587),
            .I(N__29584));
    CascadeMux I__4528 (
            .O(N__29584),
            .I(N__29581));
    CascadeBuf I__4527 (
            .O(N__29581),
            .I(N__29578));
    CascadeMux I__4526 (
            .O(N__29578),
            .I(N__29575));
    CascadeBuf I__4525 (
            .O(N__29575),
            .I(N__29572));
    CascadeMux I__4524 (
            .O(N__29572),
            .I(N__29569));
    CascadeBuf I__4523 (
            .O(N__29569),
            .I(N__29566));
    CascadeMux I__4522 (
            .O(N__29566),
            .I(N__29563));
    CascadeBuf I__4521 (
            .O(N__29563),
            .I(N__29560));
    CascadeMux I__4520 (
            .O(N__29560),
            .I(N__29557));
    CascadeBuf I__4519 (
            .O(N__29557),
            .I(N__29553));
    CascadeMux I__4518 (
            .O(N__29556),
            .I(N__29550));
    CascadeMux I__4517 (
            .O(N__29553),
            .I(N__29547));
    CascadeBuf I__4516 (
            .O(N__29550),
            .I(N__29544));
    InMux I__4515 (
            .O(N__29547),
            .I(N__29541));
    CascadeMux I__4514 (
            .O(N__29544),
            .I(N__29538));
    LocalMux I__4513 (
            .O(N__29541),
            .I(N__29535));
    InMux I__4512 (
            .O(N__29538),
            .I(N__29532));
    Span4Mux_v I__4511 (
            .O(N__29535),
            .I(N__29529));
    LocalMux I__4510 (
            .O(N__29532),
            .I(N__29526));
    Span4Mux_h I__4509 (
            .O(N__29529),
            .I(N__29523));
    Span4Mux_v I__4508 (
            .O(N__29526),
            .I(N__29519));
    Span4Mux_h I__4507 (
            .O(N__29523),
            .I(N__29516));
    InMux I__4506 (
            .O(N__29522),
            .I(N__29513));
    Span4Mux_h I__4505 (
            .O(N__29519),
            .I(N__29510));
    Span4Mux_h I__4504 (
            .O(N__29516),
            .I(N__29507));
    LocalMux I__4503 (
            .O(N__29513),
            .I(data_count_1));
    Odrv4 I__4502 (
            .O(N__29510),
            .I(data_count_1));
    Odrv4 I__4501 (
            .O(N__29507),
            .I(data_count_1));
    InMux I__4500 (
            .O(N__29500),
            .I(n20613));
    CascadeMux I__4499 (
            .O(N__29497),
            .I(N__29494));
    CascadeBuf I__4498 (
            .O(N__29494),
            .I(N__29491));
    CascadeMux I__4497 (
            .O(N__29491),
            .I(N__29488));
    CascadeBuf I__4496 (
            .O(N__29488),
            .I(N__29485));
    CascadeMux I__4495 (
            .O(N__29485),
            .I(N__29482));
    CascadeBuf I__4494 (
            .O(N__29482),
            .I(N__29479));
    CascadeMux I__4493 (
            .O(N__29479),
            .I(N__29476));
    CascadeBuf I__4492 (
            .O(N__29476),
            .I(N__29473));
    CascadeMux I__4491 (
            .O(N__29473),
            .I(N__29470));
    CascadeBuf I__4490 (
            .O(N__29470),
            .I(N__29467));
    CascadeMux I__4489 (
            .O(N__29467),
            .I(N__29464));
    CascadeBuf I__4488 (
            .O(N__29464),
            .I(N__29461));
    CascadeMux I__4487 (
            .O(N__29461),
            .I(N__29458));
    CascadeBuf I__4486 (
            .O(N__29458),
            .I(N__29455));
    CascadeMux I__4485 (
            .O(N__29455),
            .I(N__29452));
    CascadeBuf I__4484 (
            .O(N__29452),
            .I(N__29449));
    CascadeMux I__4483 (
            .O(N__29449),
            .I(N__29445));
    CascadeMux I__4482 (
            .O(N__29448),
            .I(N__29442));
    CascadeBuf I__4481 (
            .O(N__29445),
            .I(N__29439));
    CascadeBuf I__4480 (
            .O(N__29442),
            .I(N__29436));
    CascadeMux I__4479 (
            .O(N__29439),
            .I(N__29433));
    CascadeMux I__4478 (
            .O(N__29436),
            .I(N__29430));
    InMux I__4477 (
            .O(N__29433),
            .I(N__29427));
    InMux I__4476 (
            .O(N__29430),
            .I(N__29424));
    LocalMux I__4475 (
            .O(N__29427),
            .I(N__29421));
    LocalMux I__4474 (
            .O(N__29424),
            .I(N__29418));
    Sp12to4 I__4473 (
            .O(N__29421),
            .I(N__29415));
    Span4Mux_v I__4472 (
            .O(N__29418),
            .I(N__29411));
    Span12Mux_v I__4471 (
            .O(N__29415),
            .I(N__29408));
    InMux I__4470 (
            .O(N__29414),
            .I(N__29405));
    Span4Mux_h I__4469 (
            .O(N__29411),
            .I(N__29402));
    Span12Mux_h I__4468 (
            .O(N__29408),
            .I(N__29399));
    LocalMux I__4467 (
            .O(N__29405),
            .I(data_count_2));
    Odrv4 I__4466 (
            .O(N__29402),
            .I(data_count_2));
    Odrv12 I__4465 (
            .O(N__29399),
            .I(data_count_2));
    InMux I__4464 (
            .O(N__29392),
            .I(n20614));
    CascadeMux I__4463 (
            .O(N__29389),
            .I(N__29386));
    CascadeBuf I__4462 (
            .O(N__29386),
            .I(N__29383));
    CascadeMux I__4461 (
            .O(N__29383),
            .I(N__29380));
    CascadeBuf I__4460 (
            .O(N__29380),
            .I(N__29377));
    CascadeMux I__4459 (
            .O(N__29377),
            .I(N__29374));
    CascadeBuf I__4458 (
            .O(N__29374),
            .I(N__29371));
    CascadeMux I__4457 (
            .O(N__29371),
            .I(N__29368));
    CascadeBuf I__4456 (
            .O(N__29368),
            .I(N__29365));
    CascadeMux I__4455 (
            .O(N__29365),
            .I(N__29362));
    CascadeBuf I__4454 (
            .O(N__29362),
            .I(N__29359));
    CascadeMux I__4453 (
            .O(N__29359),
            .I(N__29356));
    CascadeBuf I__4452 (
            .O(N__29356),
            .I(N__29353));
    CascadeMux I__4451 (
            .O(N__29353),
            .I(N__29350));
    CascadeBuf I__4450 (
            .O(N__29350),
            .I(N__29347));
    CascadeMux I__4449 (
            .O(N__29347),
            .I(N__29344));
    CascadeBuf I__4448 (
            .O(N__29344),
            .I(N__29340));
    CascadeMux I__4447 (
            .O(N__29343),
            .I(N__29337));
    CascadeMux I__4446 (
            .O(N__29340),
            .I(N__29334));
    CascadeBuf I__4445 (
            .O(N__29337),
            .I(N__29331));
    CascadeBuf I__4444 (
            .O(N__29334),
            .I(N__29328));
    CascadeMux I__4443 (
            .O(N__29331),
            .I(N__29325));
    CascadeMux I__4442 (
            .O(N__29328),
            .I(N__29322));
    InMux I__4441 (
            .O(N__29325),
            .I(N__29319));
    InMux I__4440 (
            .O(N__29322),
            .I(N__29316));
    LocalMux I__4439 (
            .O(N__29319),
            .I(N__29313));
    LocalMux I__4438 (
            .O(N__29316),
            .I(N__29310));
    Span4Mux_v I__4437 (
            .O(N__29313),
            .I(N__29306));
    Span12Mux_v I__4436 (
            .O(N__29310),
            .I(N__29303));
    InMux I__4435 (
            .O(N__29309),
            .I(N__29300));
    Span4Mux_h I__4434 (
            .O(N__29306),
            .I(N__29297));
    Span12Mux_h I__4433 (
            .O(N__29303),
            .I(N__29294));
    LocalMux I__4432 (
            .O(N__29300),
            .I(data_count_3));
    Odrv4 I__4431 (
            .O(N__29297),
            .I(data_count_3));
    Odrv12 I__4430 (
            .O(N__29294),
            .I(data_count_3));
    InMux I__4429 (
            .O(N__29287),
            .I(n20615));
    CascadeMux I__4428 (
            .O(N__29284),
            .I(N__29281));
    CascadeBuf I__4427 (
            .O(N__29281),
            .I(N__29278));
    CascadeMux I__4426 (
            .O(N__29278),
            .I(N__29275));
    CascadeBuf I__4425 (
            .O(N__29275),
            .I(N__29272));
    CascadeMux I__4424 (
            .O(N__29272),
            .I(N__29269));
    CascadeBuf I__4423 (
            .O(N__29269),
            .I(N__29266));
    CascadeMux I__4422 (
            .O(N__29266),
            .I(N__29263));
    CascadeBuf I__4421 (
            .O(N__29263),
            .I(N__29260));
    CascadeMux I__4420 (
            .O(N__29260),
            .I(N__29257));
    CascadeBuf I__4419 (
            .O(N__29257),
            .I(N__29254));
    CascadeMux I__4418 (
            .O(N__29254),
            .I(N__29251));
    CascadeBuf I__4417 (
            .O(N__29251),
            .I(N__29248));
    CascadeMux I__4416 (
            .O(N__29248),
            .I(N__29245));
    CascadeBuf I__4415 (
            .O(N__29245),
            .I(N__29242));
    CascadeMux I__4414 (
            .O(N__29242),
            .I(N__29239));
    CascadeBuf I__4413 (
            .O(N__29239),
            .I(N__29235));
    CascadeMux I__4412 (
            .O(N__29238),
            .I(N__29232));
    CascadeMux I__4411 (
            .O(N__29235),
            .I(N__29229));
    CascadeBuf I__4410 (
            .O(N__29232),
            .I(N__29226));
    CascadeBuf I__4409 (
            .O(N__29229),
            .I(N__29223));
    CascadeMux I__4408 (
            .O(N__29226),
            .I(N__29220));
    CascadeMux I__4407 (
            .O(N__29223),
            .I(N__29217));
    InMux I__4406 (
            .O(N__29220),
            .I(N__29214));
    InMux I__4405 (
            .O(N__29217),
            .I(N__29211));
    LocalMux I__4404 (
            .O(N__29214),
            .I(N__29208));
    LocalMux I__4403 (
            .O(N__29211),
            .I(N__29205));
    Span4Mux_h I__4402 (
            .O(N__29208),
            .I(N__29202));
    Sp12to4 I__4401 (
            .O(N__29205),
            .I(N__29199));
    Span4Mux_h I__4400 (
            .O(N__29202),
            .I(N__29195));
    Span12Mux_s8_v I__4399 (
            .O(N__29199),
            .I(N__29192));
    InMux I__4398 (
            .O(N__29198),
            .I(N__29189));
    Sp12to4 I__4397 (
            .O(N__29195),
            .I(N__29184));
    Span12Mux_h I__4396 (
            .O(N__29192),
            .I(N__29184));
    LocalMux I__4395 (
            .O(N__29189),
            .I(data_count_4));
    Odrv12 I__4394 (
            .O(N__29184),
            .I(data_count_4));
    InMux I__4393 (
            .O(N__29179),
            .I(n20616));
    CascadeMux I__4392 (
            .O(N__29176),
            .I(N__29173));
    CascadeBuf I__4391 (
            .O(N__29173),
            .I(N__29170));
    CascadeMux I__4390 (
            .O(N__29170),
            .I(N__29167));
    CascadeBuf I__4389 (
            .O(N__29167),
            .I(N__29164));
    CascadeMux I__4388 (
            .O(N__29164),
            .I(N__29161));
    CascadeBuf I__4387 (
            .O(N__29161),
            .I(N__29158));
    CascadeMux I__4386 (
            .O(N__29158),
            .I(N__29155));
    CascadeBuf I__4385 (
            .O(N__29155),
            .I(N__29152));
    CascadeMux I__4384 (
            .O(N__29152),
            .I(N__29149));
    CascadeBuf I__4383 (
            .O(N__29149),
            .I(N__29146));
    CascadeMux I__4382 (
            .O(N__29146),
            .I(N__29143));
    CascadeBuf I__4381 (
            .O(N__29143),
            .I(N__29140));
    CascadeMux I__4380 (
            .O(N__29140),
            .I(N__29137));
    CascadeBuf I__4379 (
            .O(N__29137),
            .I(N__29134));
    CascadeMux I__4378 (
            .O(N__29134),
            .I(N__29131));
    CascadeBuf I__4377 (
            .O(N__29131),
            .I(N__29127));
    CascadeMux I__4376 (
            .O(N__29130),
            .I(N__29124));
    CascadeMux I__4375 (
            .O(N__29127),
            .I(N__29121));
    CascadeBuf I__4374 (
            .O(N__29124),
            .I(N__29118));
    CascadeBuf I__4373 (
            .O(N__29121),
            .I(N__29115));
    CascadeMux I__4372 (
            .O(N__29118),
            .I(N__29112));
    CascadeMux I__4371 (
            .O(N__29115),
            .I(N__29109));
    InMux I__4370 (
            .O(N__29112),
            .I(N__29106));
    InMux I__4369 (
            .O(N__29109),
            .I(N__29103));
    LocalMux I__4368 (
            .O(N__29106),
            .I(N__29100));
    LocalMux I__4367 (
            .O(N__29103),
            .I(N__29097));
    Span4Mux_v I__4366 (
            .O(N__29100),
            .I(N__29093));
    Span12Mux_s7_v I__4365 (
            .O(N__29097),
            .I(N__29090));
    InMux I__4364 (
            .O(N__29096),
            .I(N__29087));
    Span4Mux_h I__4363 (
            .O(N__29093),
            .I(N__29084));
    Span12Mux_h I__4362 (
            .O(N__29090),
            .I(N__29081));
    LocalMux I__4361 (
            .O(N__29087),
            .I(data_count_5));
    Odrv4 I__4360 (
            .O(N__29084),
            .I(data_count_5));
    Odrv12 I__4359 (
            .O(N__29081),
            .I(data_count_5));
    InMux I__4358 (
            .O(N__29074),
            .I(n20617));
    CascadeMux I__4357 (
            .O(N__29071),
            .I(n22164_cascade_));
    InMux I__4356 (
            .O(N__29068),
            .I(N__29063));
    InMux I__4355 (
            .O(N__29067),
            .I(N__29060));
    InMux I__4354 (
            .O(N__29066),
            .I(N__29057));
    LocalMux I__4353 (
            .O(N__29063),
            .I(N__29054));
    LocalMux I__4352 (
            .O(N__29060),
            .I(buf_dds1_14));
    LocalMux I__4351 (
            .O(N__29057),
            .I(buf_dds1_14));
    Odrv4 I__4350 (
            .O(N__29054),
            .I(buf_dds1_14));
    InMux I__4349 (
            .O(N__29047),
            .I(N__29044));
    LocalMux I__4348 (
            .O(N__29044),
            .I(N__29041));
    Span4Mux_h I__4347 (
            .O(N__29041),
            .I(N__29038));
    Odrv4 I__4346 (
            .O(N__29038),
            .I(n23366));
    CascadeMux I__4345 (
            .O(N__29035),
            .I(n16_adj_1763_cascade_));
    InMux I__4344 (
            .O(N__29032),
            .I(N__29029));
    LocalMux I__4343 (
            .O(N__29029),
            .I(n23369));
    InMux I__4342 (
            .O(N__29026),
            .I(N__29023));
    LocalMux I__4341 (
            .O(N__29023),
            .I(N__29020));
    Span4Mux_v I__4340 (
            .O(N__29020),
            .I(N__29017));
    Span4Mux_h I__4339 (
            .O(N__29017),
            .I(N__29014));
    Odrv4 I__4338 (
            .O(N__29014),
            .I(n30_adj_1698));
    CascadeMux I__4337 (
            .O(N__29011),
            .I(N__29005));
    InMux I__4336 (
            .O(N__29010),
            .I(N__28998));
    InMux I__4335 (
            .O(N__29009),
            .I(N__28998));
    InMux I__4334 (
            .O(N__29008),
            .I(N__28998));
    InMux I__4333 (
            .O(N__29005),
            .I(N__28995));
    LocalMux I__4332 (
            .O(N__28998),
            .I(N__28991));
    LocalMux I__4331 (
            .O(N__28995),
            .I(N__28988));
    CascadeMux I__4330 (
            .O(N__28994),
            .I(N__28985));
    Span4Mux_h I__4329 (
            .O(N__28991),
            .I(N__28982));
    Span12Mux_h I__4328 (
            .O(N__28988),
            .I(N__28979));
    InMux I__4327 (
            .O(N__28985),
            .I(N__28976));
    Span4Mux_v I__4326 (
            .O(N__28982),
            .I(N__28973));
    Odrv12 I__4325 (
            .O(N__28979),
            .I(buf_cfgRTD_6));
    LocalMux I__4324 (
            .O(N__28976),
            .I(buf_cfgRTD_6));
    Odrv4 I__4323 (
            .O(N__28973),
            .I(buf_cfgRTD_6));
    CascadeMux I__4322 (
            .O(N__28966),
            .I(N__28962));
    CascadeMux I__4321 (
            .O(N__28965),
            .I(N__28959));
    InMux I__4320 (
            .O(N__28962),
            .I(N__28954));
    InMux I__4319 (
            .O(N__28959),
            .I(N__28954));
    LocalMux I__4318 (
            .O(N__28954),
            .I(N__28950));
    InMux I__4317 (
            .O(N__28953),
            .I(N__28947));
    Span4Mux_v I__4316 (
            .O(N__28950),
            .I(N__28942));
    LocalMux I__4315 (
            .O(N__28947),
            .I(N__28942));
    Span4Mux_h I__4314 (
            .O(N__28942),
            .I(N__28937));
    InMux I__4313 (
            .O(N__28941),
            .I(N__28934));
    InMux I__4312 (
            .O(N__28940),
            .I(N__28931));
    Odrv4 I__4311 (
            .O(N__28937),
            .I(buf_cfgRTD_2));
    LocalMux I__4310 (
            .O(N__28934),
            .I(buf_cfgRTD_2));
    LocalMux I__4309 (
            .O(N__28931),
            .I(buf_cfgRTD_2));
    CascadeMux I__4308 (
            .O(N__28924),
            .I(N__28919));
    CascadeMux I__4307 (
            .O(N__28923),
            .I(N__28916));
    InMux I__4306 (
            .O(N__28922),
            .I(N__28911));
    InMux I__4305 (
            .O(N__28919),
            .I(N__28911));
    InMux I__4304 (
            .O(N__28916),
            .I(N__28908));
    LocalMux I__4303 (
            .O(N__28911),
            .I(N__28905));
    LocalMux I__4302 (
            .O(N__28908),
            .I(N__28902));
    Span4Mux_v I__4301 (
            .O(N__28905),
            .I(N__28895));
    Span4Mux_v I__4300 (
            .O(N__28902),
            .I(N__28895));
    InMux I__4299 (
            .O(N__28901),
            .I(N__28892));
    InMux I__4298 (
            .O(N__28900),
            .I(N__28889));
    Span4Mux_h I__4297 (
            .O(N__28895),
            .I(N__28884));
    LocalMux I__4296 (
            .O(N__28892),
            .I(N__28884));
    LocalMux I__4295 (
            .O(N__28889),
            .I(buf_cfgRTD_4));
    Odrv4 I__4294 (
            .O(N__28884),
            .I(buf_cfgRTD_4));
    InMux I__4293 (
            .O(N__28879),
            .I(N__28876));
    LocalMux I__4292 (
            .O(N__28876),
            .I(N__28872));
    InMux I__4291 (
            .O(N__28875),
            .I(N__28869));
    Odrv4 I__4290 (
            .O(N__28872),
            .I(\comm_spi.n24028 ));
    LocalMux I__4289 (
            .O(N__28869),
            .I(\comm_spi.n24028 ));
    CascadeMux I__4288 (
            .O(N__28864),
            .I(\comm_spi.n24028_cascade_ ));
    InMux I__4287 (
            .O(N__28861),
            .I(N__28858));
    LocalMux I__4286 (
            .O(N__28858),
            .I(N__28855));
    Span4Mux_h I__4285 (
            .O(N__28855),
            .I(N__28852));
    Span4Mux_v I__4284 (
            .O(N__28852),
            .I(N__28848));
    CascadeMux I__4283 (
            .O(N__28851),
            .I(N__28845));
    Sp12to4 I__4282 (
            .O(N__28848),
            .I(N__28842));
    InMux I__4281 (
            .O(N__28845),
            .I(N__28839));
    Odrv12 I__4280 (
            .O(N__28842),
            .I(buf_readRTD_12));
    LocalMux I__4279 (
            .O(N__28839),
            .I(buf_readRTD_12));
    CascadeMux I__4278 (
            .O(N__28834),
            .I(N__28831));
    InMux I__4277 (
            .O(N__28831),
            .I(N__28828));
    LocalMux I__4276 (
            .O(N__28828),
            .I(n20_adj_1781));
    CascadeMux I__4275 (
            .O(N__28825),
            .I(N__28822));
    InMux I__4274 (
            .O(N__28822),
            .I(N__28818));
    CascadeMux I__4273 (
            .O(N__28821),
            .I(N__28815));
    LocalMux I__4272 (
            .O(N__28818),
            .I(N__28812));
    InMux I__4271 (
            .O(N__28815),
            .I(N__28809));
    Span4Mux_h I__4270 (
            .O(N__28812),
            .I(N__28806));
    LocalMux I__4269 (
            .O(N__28809),
            .I(N__28802));
    Span4Mux_h I__4268 (
            .O(N__28806),
            .I(N__28799));
    InMux I__4267 (
            .O(N__28805),
            .I(N__28796));
    Odrv12 I__4266 (
            .O(N__28802),
            .I(cmd_rdadctmp_19_adj_1529));
    Odrv4 I__4265 (
            .O(N__28799),
            .I(cmd_rdadctmp_19_adj_1529));
    LocalMux I__4264 (
            .O(N__28796),
            .I(cmd_rdadctmp_19_adj_1529));
    CascadeMux I__4263 (
            .O(N__28789),
            .I(N__28785));
    CascadeMux I__4262 (
            .O(N__28788),
            .I(N__28782));
    InMux I__4261 (
            .O(N__28785),
            .I(N__28779));
    InMux I__4260 (
            .O(N__28782),
            .I(N__28776));
    LocalMux I__4259 (
            .O(N__28779),
            .I(N__28773));
    LocalMux I__4258 (
            .O(N__28776),
            .I(N__28770));
    Span4Mux_v I__4257 (
            .O(N__28773),
            .I(N__28764));
    Span4Mux_h I__4256 (
            .O(N__28770),
            .I(N__28764));
    InMux I__4255 (
            .O(N__28769),
            .I(N__28761));
    Odrv4 I__4254 (
            .O(N__28764),
            .I(cmd_rdadctmp_20_adj_1528));
    LocalMux I__4253 (
            .O(N__28761),
            .I(cmd_rdadctmp_20_adj_1528));
    InMux I__4252 (
            .O(N__28756),
            .I(N__28753));
    LocalMux I__4251 (
            .O(N__28753),
            .I(n23309));
    InMux I__4250 (
            .O(N__28750),
            .I(N__28747));
    LocalMux I__4249 (
            .O(N__28747),
            .I(N__28744));
    Span4Mux_v I__4248 (
            .O(N__28744),
            .I(N__28741));
    Sp12to4 I__4247 (
            .O(N__28741),
            .I(N__28737));
    CascadeMux I__4246 (
            .O(N__28740),
            .I(N__28734));
    Span12Mux_h I__4245 (
            .O(N__28737),
            .I(N__28731));
    InMux I__4244 (
            .O(N__28734),
            .I(N__28728));
    Odrv12 I__4243 (
            .O(N__28731),
            .I(buf_readRTD_10));
    LocalMux I__4242 (
            .O(N__28728),
            .I(buf_readRTD_10));
    InMux I__4241 (
            .O(N__28723),
            .I(N__28719));
    InMux I__4240 (
            .O(N__28722),
            .I(N__28715));
    LocalMux I__4239 (
            .O(N__28719),
            .I(N__28712));
    InMux I__4238 (
            .O(N__28718),
            .I(N__28709));
    LocalMux I__4237 (
            .O(N__28715),
            .I(N__28706));
    Span4Mux_v I__4236 (
            .O(N__28712),
            .I(N__28703));
    LocalMux I__4235 (
            .O(N__28709),
            .I(buf_dds1_5));
    Odrv4 I__4234 (
            .O(N__28706),
            .I(buf_dds1_5));
    Odrv4 I__4233 (
            .O(N__28703),
            .I(buf_dds1_5));
    InMux I__4232 (
            .O(N__28696),
            .I(N__28693));
    LocalMux I__4231 (
            .O(N__28693),
            .I(N__28689));
    CascadeMux I__4230 (
            .O(N__28692),
            .I(N__28686));
    Span4Mux_v I__4229 (
            .O(N__28689),
            .I(N__28683));
    InMux I__4228 (
            .O(N__28686),
            .I(N__28680));
    Odrv4 I__4227 (
            .O(N__28683),
            .I(buf_adcdata_vdc_14));
    LocalMux I__4226 (
            .O(N__28680),
            .I(buf_adcdata_vdc_14));
    InMux I__4225 (
            .O(N__28675),
            .I(N__28672));
    LocalMux I__4224 (
            .O(N__28672),
            .I(N__28668));
    InMux I__4223 (
            .O(N__28671),
            .I(N__28665));
    Span12Mux_s10_h I__4222 (
            .O(N__28668),
            .I(N__28661));
    LocalMux I__4221 (
            .O(N__28665),
            .I(N__28658));
    InMux I__4220 (
            .O(N__28664),
            .I(N__28655));
    Span12Mux_h I__4219 (
            .O(N__28661),
            .I(N__28652));
    Span4Mux_h I__4218 (
            .O(N__28658),
            .I(N__28649));
    LocalMux I__4217 (
            .O(N__28655),
            .I(buf_adcdata_vac_14));
    Odrv12 I__4216 (
            .O(N__28652),
            .I(buf_adcdata_vac_14));
    Odrv4 I__4215 (
            .O(N__28649),
            .I(buf_adcdata_vac_14));
    CEMux I__4214 (
            .O(N__28642),
            .I(N__28639));
    LocalMux I__4213 (
            .O(N__28639),
            .I(N__28633));
    CEMux I__4212 (
            .O(N__28638),
            .I(N__28630));
    CEMux I__4211 (
            .O(N__28637),
            .I(N__28627));
    CEMux I__4210 (
            .O(N__28636),
            .I(N__28622));
    Span4Mux_v I__4209 (
            .O(N__28633),
            .I(N__28616));
    LocalMux I__4208 (
            .O(N__28630),
            .I(N__28616));
    LocalMux I__4207 (
            .O(N__28627),
            .I(N__28613));
    CEMux I__4206 (
            .O(N__28626),
            .I(N__28610));
    CEMux I__4205 (
            .O(N__28625),
            .I(N__28607));
    LocalMux I__4204 (
            .O(N__28622),
            .I(N__28604));
    CEMux I__4203 (
            .O(N__28621),
            .I(N__28601));
    Span4Mux_v I__4202 (
            .O(N__28616),
            .I(N__28598));
    Span4Mux_v I__4201 (
            .O(N__28613),
            .I(N__28593));
    LocalMux I__4200 (
            .O(N__28610),
            .I(N__28593));
    LocalMux I__4199 (
            .O(N__28607),
            .I(N__28590));
    Span4Mux_v I__4198 (
            .O(N__28604),
            .I(N__28582));
    LocalMux I__4197 (
            .O(N__28601),
            .I(N__28582));
    Span4Mux_v I__4196 (
            .O(N__28598),
            .I(N__28582));
    Span4Mux_v I__4195 (
            .O(N__28593),
            .I(N__28579));
    Span4Mux_h I__4194 (
            .O(N__28590),
            .I(N__28576));
    InMux I__4193 (
            .O(N__28589),
            .I(N__28573));
    Odrv4 I__4192 (
            .O(N__28582),
            .I(\ADC_VDC.n14120 ));
    Odrv4 I__4191 (
            .O(N__28579),
            .I(\ADC_VDC.n14120 ));
    Odrv4 I__4190 (
            .O(N__28576),
            .I(\ADC_VDC.n14120 ));
    LocalMux I__4189 (
            .O(N__28573),
            .I(\ADC_VDC.n14120 ));
    SRMux I__4188 (
            .O(N__28564),
            .I(N__28558));
    SRMux I__4187 (
            .O(N__28563),
            .I(N__28554));
    SRMux I__4186 (
            .O(N__28562),
            .I(N__28550));
    SRMux I__4185 (
            .O(N__28561),
            .I(N__28546));
    LocalMux I__4184 (
            .O(N__28558),
            .I(N__28543));
    SRMux I__4183 (
            .O(N__28557),
            .I(N__28540));
    LocalMux I__4182 (
            .O(N__28554),
            .I(N__28537));
    SRMux I__4181 (
            .O(N__28553),
            .I(N__28534));
    LocalMux I__4180 (
            .O(N__28550),
            .I(N__28531));
    SRMux I__4179 (
            .O(N__28549),
            .I(N__28528));
    LocalMux I__4178 (
            .O(N__28546),
            .I(N__28525));
    Span4Mux_h I__4177 (
            .O(N__28543),
            .I(N__28522));
    LocalMux I__4176 (
            .O(N__28540),
            .I(N__28519));
    Span4Mux_h I__4175 (
            .O(N__28537),
            .I(N__28516));
    LocalMux I__4174 (
            .O(N__28534),
            .I(N__28513));
    Span4Mux_h I__4173 (
            .O(N__28531),
            .I(N__28510));
    LocalMux I__4172 (
            .O(N__28528),
            .I(N__28507));
    Span4Mux_v I__4171 (
            .O(N__28525),
            .I(N__28504));
    Span4Mux_v I__4170 (
            .O(N__28522),
            .I(N__28497));
    Span4Mux_h I__4169 (
            .O(N__28519),
            .I(N__28497));
    Span4Mux_v I__4168 (
            .O(N__28516),
            .I(N__28497));
    Span4Mux_h I__4167 (
            .O(N__28513),
            .I(N__28492));
    Span4Mux_v I__4166 (
            .O(N__28510),
            .I(N__28492));
    Odrv12 I__4165 (
            .O(N__28507),
            .I(\ADC_VDC.n15721 ));
    Odrv4 I__4164 (
            .O(N__28504),
            .I(\ADC_VDC.n15721 ));
    Odrv4 I__4163 (
            .O(N__28497),
            .I(\ADC_VDC.n15721 ));
    Odrv4 I__4162 (
            .O(N__28492),
            .I(\ADC_VDC.n15721 ));
    InMux I__4161 (
            .O(N__28483),
            .I(N__28480));
    LocalMux I__4160 (
            .O(N__28480),
            .I(\ADC_VDC.cmd_rdadcbuf_35_N_1344_34 ));
    CascadeMux I__4159 (
            .O(N__28477),
            .I(\ADC_VDC.n4_cascade_ ));
    InMux I__4158 (
            .O(N__28474),
            .I(N__28471));
    LocalMux I__4157 (
            .O(N__28471),
            .I(N__28468));
    Span4Mux_h I__4156 (
            .O(N__28468),
            .I(N__28463));
    InMux I__4155 (
            .O(N__28467),
            .I(N__28460));
    InMux I__4154 (
            .O(N__28466),
            .I(N__28457));
    Odrv4 I__4153 (
            .O(N__28463),
            .I(cmd_rdadcbuf_34));
    LocalMux I__4152 (
            .O(N__28460),
            .I(cmd_rdadcbuf_34));
    LocalMux I__4151 (
            .O(N__28457),
            .I(cmd_rdadcbuf_34));
    CEMux I__4150 (
            .O(N__28450),
            .I(N__28447));
    LocalMux I__4149 (
            .O(N__28447),
            .I(N__28444));
    Span4Mux_h I__4148 (
            .O(N__28444),
            .I(N__28441));
    Odrv4 I__4147 (
            .O(N__28441),
            .I(\ADC_VDC.n14092 ));
    InMux I__4146 (
            .O(N__28438),
            .I(N__28434));
    InMux I__4145 (
            .O(N__28437),
            .I(N__28431));
    LocalMux I__4144 (
            .O(N__28434),
            .I(cmd_rdadcbuf_14));
    LocalMux I__4143 (
            .O(N__28431),
            .I(cmd_rdadcbuf_14));
    InMux I__4142 (
            .O(N__28426),
            .I(N__28422));
    CascadeMux I__4141 (
            .O(N__28425),
            .I(N__28418));
    LocalMux I__4140 (
            .O(N__28422),
            .I(N__28415));
    InMux I__4139 (
            .O(N__28421),
            .I(N__28412));
    InMux I__4138 (
            .O(N__28418),
            .I(N__28409));
    Odrv4 I__4137 (
            .O(N__28415),
            .I(cmd_rdadctmp_8_adj_1566));
    LocalMux I__4136 (
            .O(N__28412),
            .I(cmd_rdadctmp_8_adj_1566));
    LocalMux I__4135 (
            .O(N__28409),
            .I(cmd_rdadctmp_8_adj_1566));
    CascadeMux I__4134 (
            .O(N__28402),
            .I(N__28398));
    CascadeMux I__4133 (
            .O(N__28401),
            .I(N__28387));
    InMux I__4132 (
            .O(N__28398),
            .I(N__28382));
    CascadeMux I__4131 (
            .O(N__28397),
            .I(N__28376));
    CascadeMux I__4130 (
            .O(N__28396),
            .I(N__28373));
    CascadeMux I__4129 (
            .O(N__28395),
            .I(N__28367));
    CascadeMux I__4128 (
            .O(N__28394),
            .I(N__28364));
    CascadeMux I__4127 (
            .O(N__28393),
            .I(N__28361));
    InMux I__4126 (
            .O(N__28392),
            .I(N__28348));
    InMux I__4125 (
            .O(N__28391),
            .I(N__28348));
    InMux I__4124 (
            .O(N__28390),
            .I(N__28348));
    InMux I__4123 (
            .O(N__28387),
            .I(N__28348));
    InMux I__4122 (
            .O(N__28386),
            .I(N__28348));
    InMux I__4121 (
            .O(N__28385),
            .I(N__28348));
    LocalMux I__4120 (
            .O(N__28382),
            .I(N__28345));
    CascadeMux I__4119 (
            .O(N__28381),
            .I(N__28339));
    InMux I__4118 (
            .O(N__28380),
            .I(N__28328));
    InMux I__4117 (
            .O(N__28379),
            .I(N__28328));
    InMux I__4116 (
            .O(N__28376),
            .I(N__28328));
    InMux I__4115 (
            .O(N__28373),
            .I(N__28328));
    InMux I__4114 (
            .O(N__28372),
            .I(N__28315));
    InMux I__4113 (
            .O(N__28371),
            .I(N__28315));
    InMux I__4112 (
            .O(N__28370),
            .I(N__28315));
    InMux I__4111 (
            .O(N__28367),
            .I(N__28315));
    InMux I__4110 (
            .O(N__28364),
            .I(N__28315));
    InMux I__4109 (
            .O(N__28361),
            .I(N__28315));
    LocalMux I__4108 (
            .O(N__28348),
            .I(N__28310));
    Span4Mux_h I__4107 (
            .O(N__28345),
            .I(N__28310));
    InMux I__4106 (
            .O(N__28344),
            .I(N__28297));
    InMux I__4105 (
            .O(N__28343),
            .I(N__28297));
    InMux I__4104 (
            .O(N__28342),
            .I(N__28297));
    InMux I__4103 (
            .O(N__28339),
            .I(N__28297));
    InMux I__4102 (
            .O(N__28338),
            .I(N__28297));
    InMux I__4101 (
            .O(N__28337),
            .I(N__28297));
    LocalMux I__4100 (
            .O(N__28328),
            .I(N__28292));
    LocalMux I__4099 (
            .O(N__28315),
            .I(N__28292));
    Odrv4 I__4098 (
            .O(N__28310),
            .I(n13925));
    LocalMux I__4097 (
            .O(N__28297),
            .I(n13925));
    Odrv12 I__4096 (
            .O(N__28292),
            .I(n13925));
    InMux I__4095 (
            .O(N__28285),
            .I(N__28282));
    LocalMux I__4094 (
            .O(N__28282),
            .I(N__28278));
    CascadeMux I__4093 (
            .O(N__28281),
            .I(N__28274));
    Span4Mux_h I__4092 (
            .O(N__28278),
            .I(N__28271));
    InMux I__4091 (
            .O(N__28277),
            .I(N__28268));
    InMux I__4090 (
            .O(N__28274),
            .I(N__28265));
    Odrv4 I__4089 (
            .O(N__28271),
            .I(cmd_rdadctmp_9_adj_1565));
    LocalMux I__4088 (
            .O(N__28268),
            .I(cmd_rdadctmp_9_adj_1565));
    LocalMux I__4087 (
            .O(N__28265),
            .I(cmd_rdadctmp_9_adj_1565));
    CascadeMux I__4086 (
            .O(N__28258),
            .I(N__28255));
    InMux I__4085 (
            .O(N__28255),
            .I(N__28251));
    InMux I__4084 (
            .O(N__28254),
            .I(N__28248));
    LocalMux I__4083 (
            .O(N__28251),
            .I(cmd_rdadcbuf_22));
    LocalMux I__4082 (
            .O(N__28248),
            .I(cmd_rdadcbuf_22));
    InMux I__4081 (
            .O(N__28243),
            .I(N__28239));
    InMux I__4080 (
            .O(N__28242),
            .I(N__28236));
    LocalMux I__4079 (
            .O(N__28239),
            .I(cmd_rdadcbuf_13));
    LocalMux I__4078 (
            .O(N__28236),
            .I(cmd_rdadcbuf_13));
    CascadeMux I__4077 (
            .O(N__28231),
            .I(N__28228));
    InMux I__4076 (
            .O(N__28228),
            .I(N__28224));
    InMux I__4075 (
            .O(N__28227),
            .I(N__28221));
    LocalMux I__4074 (
            .O(N__28224),
            .I(cmd_rdadcbuf_16));
    LocalMux I__4073 (
            .O(N__28221),
            .I(cmd_rdadcbuf_16));
    InMux I__4072 (
            .O(N__28216),
            .I(N__28213));
    LocalMux I__4071 (
            .O(N__28213),
            .I(N__28210));
    Span4Mux_v I__4070 (
            .O(N__28210),
            .I(N__28207));
    Span4Mux_h I__4069 (
            .O(N__28207),
            .I(N__28203));
    InMux I__4068 (
            .O(N__28206),
            .I(N__28200));
    Odrv4 I__4067 (
            .O(N__28203),
            .I(buf_adcdata_vdc_5));
    LocalMux I__4066 (
            .O(N__28200),
            .I(buf_adcdata_vdc_5));
    InMux I__4065 (
            .O(N__28195),
            .I(N__28192));
    LocalMux I__4064 (
            .O(N__28192),
            .I(N__28188));
    InMux I__4063 (
            .O(N__28191),
            .I(N__28185));
    Odrv4 I__4062 (
            .O(N__28188),
            .I(cmd_rdadcbuf_27));
    LocalMux I__4061 (
            .O(N__28185),
            .I(cmd_rdadcbuf_27));
    InMux I__4060 (
            .O(N__28180),
            .I(N__28176));
    InMux I__4059 (
            .O(N__28179),
            .I(N__28173));
    LocalMux I__4058 (
            .O(N__28176),
            .I(\ADC_VDC.avg_cnt_10 ));
    LocalMux I__4057 (
            .O(N__28173),
            .I(\ADC_VDC.avg_cnt_10 ));
    InMux I__4056 (
            .O(N__28168),
            .I(N__28165));
    LocalMux I__4055 (
            .O(N__28165),
            .I(N__28162));
    Odrv4 I__4054 (
            .O(N__28162),
            .I(\ADC_VDC.n20 ));
    CascadeMux I__4053 (
            .O(N__28159),
            .I(\ADC_VDC.n19_cascade_ ));
    InMux I__4052 (
            .O(N__28156),
            .I(N__28153));
    LocalMux I__4051 (
            .O(N__28153),
            .I(N__28150));
    Odrv4 I__4050 (
            .O(N__28150),
            .I(\ADC_VDC.n21 ));
    InMux I__4049 (
            .O(N__28147),
            .I(N__28144));
    LocalMux I__4048 (
            .O(N__28144),
            .I(\ADC_VDC.n28 ));
    CEMux I__4047 (
            .O(N__28141),
            .I(N__28138));
    LocalMux I__4046 (
            .O(N__28138),
            .I(N__28135));
    Odrv4 I__4045 (
            .O(N__28135),
            .I(\ADC_VDC.n21871 ));
    CEMux I__4044 (
            .O(N__28132),
            .I(N__28129));
    LocalMux I__4043 (
            .O(N__28129),
            .I(\ADC_VDC.n13865 ));
    CascadeMux I__4042 (
            .O(N__28126),
            .I(\ADC_VDC.n9_cascade_ ));
    InMux I__4041 (
            .O(N__28123),
            .I(N__28118));
    InMux I__4040 (
            .O(N__28122),
            .I(N__28113));
    InMux I__4039 (
            .O(N__28121),
            .I(N__28113));
    LocalMux I__4038 (
            .O(N__28118),
            .I(\ADC_VDC.n22071 ));
    LocalMux I__4037 (
            .O(N__28113),
            .I(\ADC_VDC.n22071 ));
    SRMux I__4036 (
            .O(N__28108),
            .I(N__28105));
    LocalMux I__4035 (
            .O(N__28105),
            .I(N__28102));
    Span4Mux_h I__4034 (
            .O(N__28102),
            .I(N__28099));
    Odrv4 I__4033 (
            .O(N__28099),
            .I(\ADC_VDC.n5 ));
    CascadeMux I__4032 (
            .O(N__28096),
            .I(N__28093));
    InMux I__4031 (
            .O(N__28093),
            .I(N__28090));
    LocalMux I__4030 (
            .O(N__28090),
            .I(N__28085));
    InMux I__4029 (
            .O(N__28089),
            .I(N__28080));
    InMux I__4028 (
            .O(N__28088),
            .I(N__28080));
    Odrv4 I__4027 (
            .O(N__28085),
            .I(cmd_rdadctmp_21));
    LocalMux I__4026 (
            .O(N__28080),
            .I(cmd_rdadctmp_21));
    InMux I__4025 (
            .O(N__28075),
            .I(N__28070));
    InMux I__4024 (
            .O(N__28074),
            .I(N__28065));
    InMux I__4023 (
            .O(N__28073),
            .I(N__28065));
    LocalMux I__4022 (
            .O(N__28070),
            .I(cmd_rdadctmp_22));
    LocalMux I__4021 (
            .O(N__28065),
            .I(cmd_rdadctmp_22));
    CascadeMux I__4020 (
            .O(N__28060),
            .I(N__28056));
    InMux I__4019 (
            .O(N__28059),
            .I(N__28048));
    InMux I__4018 (
            .O(N__28056),
            .I(N__28048));
    InMux I__4017 (
            .O(N__28055),
            .I(N__28048));
    LocalMux I__4016 (
            .O(N__28048),
            .I(cmd_rdadctmp_23));
    InMux I__4015 (
            .O(N__28045),
            .I(N__28041));
    InMux I__4014 (
            .O(N__28044),
            .I(N__28038));
    LocalMux I__4013 (
            .O(N__28041),
            .I(\ADC_VDC.avg_cnt_0 ));
    LocalMux I__4012 (
            .O(N__28038),
            .I(\ADC_VDC.avg_cnt_0 ));
    InMux I__4011 (
            .O(N__28033),
            .I(N__28029));
    InMux I__4010 (
            .O(N__28032),
            .I(N__28026));
    LocalMux I__4009 (
            .O(N__28029),
            .I(\ADC_VDC.avg_cnt_5 ));
    LocalMux I__4008 (
            .O(N__28026),
            .I(\ADC_VDC.avg_cnt_5 ));
    CascadeMux I__4007 (
            .O(N__28021),
            .I(N__28018));
    InMux I__4006 (
            .O(N__28018),
            .I(N__28014));
    InMux I__4005 (
            .O(N__28017),
            .I(N__28011));
    LocalMux I__4004 (
            .O(N__28014),
            .I(N__28008));
    LocalMux I__4003 (
            .O(N__28011),
            .I(\ADC_VDC.avg_cnt_8 ));
    Odrv4 I__4002 (
            .O(N__28008),
            .I(\ADC_VDC.avg_cnt_8 ));
    InMux I__4001 (
            .O(N__28003),
            .I(N__28000));
    LocalMux I__4000 (
            .O(N__28000),
            .I(N__27997));
    Span4Mux_v I__3999 (
            .O(N__27997),
            .I(N__27994));
    Span4Mux_v I__3998 (
            .O(N__27994),
            .I(N__27989));
    InMux I__3997 (
            .O(N__27993),
            .I(N__27986));
    InMux I__3996 (
            .O(N__27992),
            .I(N__27983));
    Sp12to4 I__3995 (
            .O(N__27989),
            .I(N__27980));
    LocalMux I__3994 (
            .O(N__27986),
            .I(N__27977));
    LocalMux I__3993 (
            .O(N__27983),
            .I(buf_adcdata_iac_19));
    Odrv12 I__3992 (
            .O(N__27980),
            .I(buf_adcdata_iac_19));
    Odrv4 I__3991 (
            .O(N__27977),
            .I(buf_adcdata_iac_19));
    InMux I__3990 (
            .O(N__27970),
            .I(N__27965));
    InMux I__3989 (
            .O(N__27969),
            .I(N__27962));
    InMux I__3988 (
            .O(N__27968),
            .I(N__27959));
    LocalMux I__3987 (
            .O(N__27965),
            .I(N__27956));
    LocalMux I__3986 (
            .O(N__27962),
            .I(N__27953));
    LocalMux I__3985 (
            .O(N__27959),
            .I(buf_dds1_12));
    Odrv4 I__3984 (
            .O(N__27956),
            .I(buf_dds1_12));
    Odrv12 I__3983 (
            .O(N__27953),
            .I(buf_dds1_12));
    CascadeMux I__3982 (
            .O(N__27946),
            .I(N__27943));
    InMux I__3981 (
            .O(N__27943),
            .I(N__27940));
    LocalMux I__3980 (
            .O(N__27940),
            .I(N__27937));
    Odrv4 I__3979 (
            .O(N__27937),
            .I(n16_adj_1778));
    CascadeMux I__3978 (
            .O(N__27934),
            .I(N__27931));
    InMux I__3977 (
            .O(N__27931),
            .I(N__27928));
    LocalMux I__3976 (
            .O(N__27928),
            .I(N__27923));
    InMux I__3975 (
            .O(N__27927),
            .I(N__27918));
    InMux I__3974 (
            .O(N__27926),
            .I(N__27918));
    Odrv12 I__3973 (
            .O(N__27923),
            .I(cmd_rdadctmp_26));
    LocalMux I__3972 (
            .O(N__27918),
            .I(cmd_rdadctmp_26));
    InMux I__3971 (
            .O(N__27913),
            .I(N__27910));
    LocalMux I__3970 (
            .O(N__27910),
            .I(N__27905));
    InMux I__3969 (
            .O(N__27909),
            .I(N__27902));
    InMux I__3968 (
            .O(N__27908),
            .I(N__27899));
    Span4Mux_h I__3967 (
            .O(N__27905),
            .I(N__27896));
    LocalMux I__3966 (
            .O(N__27902),
            .I(buf_dds1_7));
    LocalMux I__3965 (
            .O(N__27899),
            .I(buf_dds1_7));
    Odrv4 I__3964 (
            .O(N__27896),
            .I(buf_dds1_7));
    IoInMux I__3963 (
            .O(N__27889),
            .I(N__27886));
    LocalMux I__3962 (
            .O(N__27886),
            .I(N__27882));
    CascadeMux I__3961 (
            .O(N__27885),
            .I(N__27879));
    Span12Mux_s9_v I__3960 (
            .O(N__27882),
            .I(N__27876));
    InMux I__3959 (
            .O(N__27879),
            .I(N__27873));
    Odrv12 I__3958 (
            .O(N__27876),
            .I(IAC_SCLK));
    LocalMux I__3957 (
            .O(N__27873),
            .I(IAC_SCLK));
    CascadeMux I__3956 (
            .O(N__27868),
            .I(N__27865));
    InMux I__3955 (
            .O(N__27865),
            .I(N__27862));
    LocalMux I__3954 (
            .O(N__27862),
            .I(N__27858));
    CascadeMux I__3953 (
            .O(N__27861),
            .I(N__27855));
    Span4Mux_v I__3952 (
            .O(N__27858),
            .I(N__27851));
    InMux I__3951 (
            .O(N__27855),
            .I(N__27846));
    InMux I__3950 (
            .O(N__27854),
            .I(N__27846));
    Odrv4 I__3949 (
            .O(N__27851),
            .I(cmd_rdadctmp_27_adj_1521));
    LocalMux I__3948 (
            .O(N__27846),
            .I(cmd_rdadctmp_27_adj_1521));
    InMux I__3947 (
            .O(N__27841),
            .I(N__27838));
    LocalMux I__3946 (
            .O(N__27838),
            .I(N__27835));
    Span4Mux_v I__3945 (
            .O(N__27835),
            .I(N__27832));
    Span4Mux_h I__3944 (
            .O(N__27832),
            .I(N__27829));
    Span4Mux_h I__3943 (
            .O(N__27829),
            .I(N__27825));
    InMux I__3942 (
            .O(N__27828),
            .I(N__27821));
    Span4Mux_h I__3941 (
            .O(N__27825),
            .I(N__27818));
    InMux I__3940 (
            .O(N__27824),
            .I(N__27815));
    LocalMux I__3939 (
            .O(N__27821),
            .I(buf_adcdata_vac_19));
    Odrv4 I__3938 (
            .O(N__27818),
            .I(buf_adcdata_vac_19));
    LocalMux I__3937 (
            .O(N__27815),
            .I(buf_adcdata_vac_19));
    CascadeMux I__3936 (
            .O(N__27808),
            .I(n23474_cascade_));
    CascadeMux I__3935 (
            .O(N__27805),
            .I(n23477_cascade_));
    InMux I__3934 (
            .O(N__27802),
            .I(N__27799));
    LocalMux I__3933 (
            .O(N__27799),
            .I(n30_adj_1784));
    InMux I__3932 (
            .O(N__27796),
            .I(N__27793));
    LocalMux I__3931 (
            .O(N__27793),
            .I(N__27790));
    Odrv4 I__3930 (
            .O(N__27790),
            .I(n112_adj_1772));
    CascadeMux I__3929 (
            .O(N__27787),
            .I(n30_adj_1768_cascade_));
    InMux I__3928 (
            .O(N__27784),
            .I(N__27781));
    LocalMux I__3927 (
            .O(N__27781),
            .I(n19_adj_1780));
    InMux I__3926 (
            .O(N__27778),
            .I(N__27775));
    LocalMux I__3925 (
            .O(N__27775),
            .I(N__27772));
    Span4Mux_h I__3924 (
            .O(N__27772),
            .I(N__27769));
    Span4Mux_h I__3923 (
            .O(N__27769),
            .I(N__27766));
    Odrv4 I__3922 (
            .O(N__27766),
            .I(n30_adj_1702));
    InMux I__3921 (
            .O(N__27763),
            .I(N__27760));
    LocalMux I__3920 (
            .O(N__27760),
            .I(n22358));
    InMux I__3919 (
            .O(N__27757),
            .I(N__27754));
    LocalMux I__3918 (
            .O(N__27754),
            .I(N__27750));
    CascadeMux I__3917 (
            .O(N__27753),
            .I(N__27747));
    Span4Mux_v I__3916 (
            .O(N__27750),
            .I(N__27744));
    InMux I__3915 (
            .O(N__27747),
            .I(N__27741));
    Odrv4 I__3914 (
            .O(N__27744),
            .I(buf_adcdata_vdc_19));
    LocalMux I__3913 (
            .O(N__27741),
            .I(buf_adcdata_vdc_19));
    InMux I__3912 (
            .O(N__27736),
            .I(N__27733));
    LocalMux I__3911 (
            .O(N__27733),
            .I(n19_adj_1789));
    InMux I__3910 (
            .O(N__27730),
            .I(N__27727));
    LocalMux I__3909 (
            .O(N__27727),
            .I(n23426));
    InMux I__3908 (
            .O(N__27724),
            .I(N__27721));
    LocalMux I__3907 (
            .O(N__27721),
            .I(n23429));
    InMux I__3906 (
            .O(N__27718),
            .I(N__27714));
    InMux I__3905 (
            .O(N__27717),
            .I(N__27711));
    LocalMux I__3904 (
            .O(N__27714),
            .I(cmd_rdadcbuf_28));
    LocalMux I__3903 (
            .O(N__27711),
            .I(cmd_rdadcbuf_28));
    InMux I__3902 (
            .O(N__27706),
            .I(\ADC_VDC.n20717 ));
    InMux I__3901 (
            .O(N__27703),
            .I(N__27699));
    InMux I__3900 (
            .O(N__27702),
            .I(N__27696));
    LocalMux I__3899 (
            .O(N__27699),
            .I(cmd_rdadcbuf_29));
    LocalMux I__3898 (
            .O(N__27696),
            .I(cmd_rdadcbuf_29));
    InMux I__3897 (
            .O(N__27691),
            .I(\ADC_VDC.n20718 ));
    InMux I__3896 (
            .O(N__27688),
            .I(N__27684));
    InMux I__3895 (
            .O(N__27687),
            .I(N__27681));
    LocalMux I__3894 (
            .O(N__27684),
            .I(cmd_rdadcbuf_30));
    LocalMux I__3893 (
            .O(N__27681),
            .I(cmd_rdadcbuf_30));
    InMux I__3892 (
            .O(N__27676),
            .I(\ADC_VDC.n20719 ));
    InMux I__3891 (
            .O(N__27673),
            .I(N__27669));
    InMux I__3890 (
            .O(N__27672),
            .I(N__27666));
    LocalMux I__3889 (
            .O(N__27669),
            .I(cmd_rdadcbuf_31));
    LocalMux I__3888 (
            .O(N__27666),
            .I(cmd_rdadcbuf_31));
    InMux I__3887 (
            .O(N__27661),
            .I(\ADC_VDC.n20720 ));
    InMux I__3886 (
            .O(N__27658),
            .I(bfn_8_10_0_));
    InMux I__3885 (
            .O(N__27655),
            .I(N__27651));
    InMux I__3884 (
            .O(N__27654),
            .I(N__27648));
    LocalMux I__3883 (
            .O(N__27651),
            .I(cmd_rdadcbuf_33));
    LocalMux I__3882 (
            .O(N__27648),
            .I(cmd_rdadcbuf_33));
    InMux I__3881 (
            .O(N__27643),
            .I(\ADC_VDC.n20722 ));
    InMux I__3880 (
            .O(N__27640),
            .I(\ADC_VDC.n20723 ));
    CascadeMux I__3879 (
            .O(N__27637),
            .I(N__27632));
    InMux I__3878 (
            .O(N__27636),
            .I(N__27627));
    InMux I__3877 (
            .O(N__27635),
            .I(N__27627));
    InMux I__3876 (
            .O(N__27632),
            .I(N__27624));
    LocalMux I__3875 (
            .O(N__27627),
            .I(cmd_rdadctmp_20_adj_1554));
    LocalMux I__3874 (
            .O(N__27624),
            .I(cmd_rdadctmp_20_adj_1554));
    InMux I__3873 (
            .O(N__27619),
            .I(N__27616));
    LocalMux I__3872 (
            .O(N__27616),
            .I(N__27612));
    InMux I__3871 (
            .O(N__27615),
            .I(N__27609));
    Odrv4 I__3870 (
            .O(N__27612),
            .I(cmd_rdadcbuf_20));
    LocalMux I__3869 (
            .O(N__27609),
            .I(cmd_rdadcbuf_20));
    InMux I__3868 (
            .O(N__27604),
            .I(\ADC_VDC.n20709 ));
    CascadeMux I__3867 (
            .O(N__27601),
            .I(N__27596));
    CascadeMux I__3866 (
            .O(N__27600),
            .I(N__27593));
    InMux I__3865 (
            .O(N__27599),
            .I(N__27590));
    InMux I__3864 (
            .O(N__27596),
            .I(N__27587));
    InMux I__3863 (
            .O(N__27593),
            .I(N__27584));
    LocalMux I__3862 (
            .O(N__27590),
            .I(cmd_rdadctmp_21_adj_1553));
    LocalMux I__3861 (
            .O(N__27587),
            .I(cmd_rdadctmp_21_adj_1553));
    LocalMux I__3860 (
            .O(N__27584),
            .I(cmd_rdadctmp_21_adj_1553));
    InMux I__3859 (
            .O(N__27577),
            .I(N__27573));
    InMux I__3858 (
            .O(N__27576),
            .I(N__27570));
    LocalMux I__3857 (
            .O(N__27573),
            .I(N__27567));
    LocalMux I__3856 (
            .O(N__27570),
            .I(N__27564));
    Odrv4 I__3855 (
            .O(N__27567),
            .I(cmd_rdadcbuf_21));
    Odrv4 I__3854 (
            .O(N__27564),
            .I(cmd_rdadcbuf_21));
    InMux I__3853 (
            .O(N__27559),
            .I(\ADC_VDC.n20710 ));
    InMux I__3852 (
            .O(N__27556),
            .I(\ADC_VDC.n20711 ));
    InMux I__3851 (
            .O(N__27553),
            .I(N__27549));
    InMux I__3850 (
            .O(N__27552),
            .I(N__27546));
    LocalMux I__3849 (
            .O(N__27549),
            .I(cmd_rdadcbuf_23));
    LocalMux I__3848 (
            .O(N__27546),
            .I(cmd_rdadcbuf_23));
    InMux I__3847 (
            .O(N__27541),
            .I(\ADC_VDC.n20712 ));
    InMux I__3846 (
            .O(N__27538),
            .I(bfn_8_9_0_));
    InMux I__3845 (
            .O(N__27535),
            .I(N__27531));
    InMux I__3844 (
            .O(N__27534),
            .I(N__27528));
    LocalMux I__3843 (
            .O(N__27531),
            .I(cmd_rdadcbuf_25));
    LocalMux I__3842 (
            .O(N__27528),
            .I(cmd_rdadcbuf_25));
    InMux I__3841 (
            .O(N__27523),
            .I(\ADC_VDC.n20714 ));
    InMux I__3840 (
            .O(N__27520),
            .I(N__27516));
    InMux I__3839 (
            .O(N__27519),
            .I(N__27513));
    LocalMux I__3838 (
            .O(N__27516),
            .I(cmd_rdadcbuf_26));
    LocalMux I__3837 (
            .O(N__27513),
            .I(cmd_rdadcbuf_26));
    InMux I__3836 (
            .O(N__27508),
            .I(\ADC_VDC.n20715 ));
    InMux I__3835 (
            .O(N__27505),
            .I(\ADC_VDC.n20716 ));
    CascadeMux I__3834 (
            .O(N__27502),
            .I(N__27497));
    CascadeMux I__3833 (
            .O(N__27501),
            .I(N__27494));
    CascadeMux I__3832 (
            .O(N__27500),
            .I(N__27491));
    InMux I__3831 (
            .O(N__27497),
            .I(N__27488));
    InMux I__3830 (
            .O(N__27494),
            .I(N__27485));
    InMux I__3829 (
            .O(N__27491),
            .I(N__27482));
    LocalMux I__3828 (
            .O(N__27488),
            .I(cmd_rdadctmp_12_adj_1562));
    LocalMux I__3827 (
            .O(N__27485),
            .I(cmd_rdadctmp_12_adj_1562));
    LocalMux I__3826 (
            .O(N__27482),
            .I(cmd_rdadctmp_12_adj_1562));
    InMux I__3825 (
            .O(N__27475),
            .I(N__27471));
    InMux I__3824 (
            .O(N__27474),
            .I(N__27468));
    LocalMux I__3823 (
            .O(N__27471),
            .I(cmd_rdadcbuf_12));
    LocalMux I__3822 (
            .O(N__27468),
            .I(cmd_rdadcbuf_12));
    InMux I__3821 (
            .O(N__27463),
            .I(\ADC_VDC.n20701 ));
    CascadeMux I__3820 (
            .O(N__27460),
            .I(N__27455));
    InMux I__3819 (
            .O(N__27459),
            .I(N__27450));
    InMux I__3818 (
            .O(N__27458),
            .I(N__27450));
    InMux I__3817 (
            .O(N__27455),
            .I(N__27447));
    LocalMux I__3816 (
            .O(N__27450),
            .I(cmd_rdadctmp_13_adj_1561));
    LocalMux I__3815 (
            .O(N__27447),
            .I(cmd_rdadctmp_13_adj_1561));
    InMux I__3814 (
            .O(N__27442),
            .I(\ADC_VDC.n20702 ));
    InMux I__3813 (
            .O(N__27439),
            .I(N__27434));
    CascadeMux I__3812 (
            .O(N__27438),
            .I(N__27431));
    InMux I__3811 (
            .O(N__27437),
            .I(N__27428));
    LocalMux I__3810 (
            .O(N__27434),
            .I(N__27425));
    InMux I__3809 (
            .O(N__27431),
            .I(N__27422));
    LocalMux I__3808 (
            .O(N__27428),
            .I(cmd_rdadctmp_14_adj_1560));
    Odrv4 I__3807 (
            .O(N__27425),
            .I(cmd_rdadctmp_14_adj_1560));
    LocalMux I__3806 (
            .O(N__27422),
            .I(cmd_rdadctmp_14_adj_1560));
    InMux I__3805 (
            .O(N__27415),
            .I(\ADC_VDC.n20703 ));
    InMux I__3804 (
            .O(N__27412),
            .I(N__27407));
    CascadeMux I__3803 (
            .O(N__27411),
            .I(N__27404));
    CascadeMux I__3802 (
            .O(N__27410),
            .I(N__27401));
    LocalMux I__3801 (
            .O(N__27407),
            .I(N__27398));
    InMux I__3800 (
            .O(N__27404),
            .I(N__27395));
    InMux I__3799 (
            .O(N__27401),
            .I(N__27392));
    Span4Mux_v I__3798 (
            .O(N__27398),
            .I(N__27389));
    LocalMux I__3797 (
            .O(N__27395),
            .I(N__27386));
    LocalMux I__3796 (
            .O(N__27392),
            .I(cmd_rdadctmp_15_adj_1559));
    Odrv4 I__3795 (
            .O(N__27389),
            .I(cmd_rdadctmp_15_adj_1559));
    Odrv4 I__3794 (
            .O(N__27386),
            .I(cmd_rdadctmp_15_adj_1559));
    InMux I__3793 (
            .O(N__27379),
            .I(N__27376));
    LocalMux I__3792 (
            .O(N__27376),
            .I(N__27372));
    InMux I__3791 (
            .O(N__27375),
            .I(N__27369));
    Odrv4 I__3790 (
            .O(N__27372),
            .I(cmd_rdadcbuf_15));
    LocalMux I__3789 (
            .O(N__27369),
            .I(cmd_rdadcbuf_15));
    InMux I__3788 (
            .O(N__27364),
            .I(\ADC_VDC.n20704 ));
    CascadeMux I__3787 (
            .O(N__27361),
            .I(N__27356));
    InMux I__3786 (
            .O(N__27360),
            .I(N__27353));
    InMux I__3785 (
            .O(N__27359),
            .I(N__27350));
    InMux I__3784 (
            .O(N__27356),
            .I(N__27347));
    LocalMux I__3783 (
            .O(N__27353),
            .I(cmd_rdadctmp_16_adj_1558));
    LocalMux I__3782 (
            .O(N__27350),
            .I(cmd_rdadctmp_16_adj_1558));
    LocalMux I__3781 (
            .O(N__27347),
            .I(cmd_rdadctmp_16_adj_1558));
    InMux I__3780 (
            .O(N__27340),
            .I(bfn_8_8_0_));
    CascadeMux I__3779 (
            .O(N__27337),
            .I(N__27333));
    CascadeMux I__3778 (
            .O(N__27336),
            .I(N__27329));
    InMux I__3777 (
            .O(N__27333),
            .I(N__27326));
    InMux I__3776 (
            .O(N__27332),
            .I(N__27323));
    InMux I__3775 (
            .O(N__27329),
            .I(N__27320));
    LocalMux I__3774 (
            .O(N__27326),
            .I(cmd_rdadctmp_17_adj_1557));
    LocalMux I__3773 (
            .O(N__27323),
            .I(cmd_rdadctmp_17_adj_1557));
    LocalMux I__3772 (
            .O(N__27320),
            .I(cmd_rdadctmp_17_adj_1557));
    InMux I__3771 (
            .O(N__27313),
            .I(N__27310));
    LocalMux I__3770 (
            .O(N__27310),
            .I(N__27306));
    InMux I__3769 (
            .O(N__27309),
            .I(N__27303));
    Odrv4 I__3768 (
            .O(N__27306),
            .I(cmd_rdadcbuf_17));
    LocalMux I__3767 (
            .O(N__27303),
            .I(cmd_rdadcbuf_17));
    InMux I__3766 (
            .O(N__27298),
            .I(\ADC_VDC.n20706 ));
    CascadeMux I__3765 (
            .O(N__27295),
            .I(N__27290));
    InMux I__3764 (
            .O(N__27294),
            .I(N__27285));
    InMux I__3763 (
            .O(N__27293),
            .I(N__27285));
    InMux I__3762 (
            .O(N__27290),
            .I(N__27282));
    LocalMux I__3761 (
            .O(N__27285),
            .I(cmd_rdadctmp_18_adj_1556));
    LocalMux I__3760 (
            .O(N__27282),
            .I(cmd_rdadctmp_18_adj_1556));
    InMux I__3759 (
            .O(N__27277),
            .I(N__27273));
    InMux I__3758 (
            .O(N__27276),
            .I(N__27270));
    LocalMux I__3757 (
            .O(N__27273),
            .I(cmd_rdadcbuf_18));
    LocalMux I__3756 (
            .O(N__27270),
            .I(cmd_rdadcbuf_18));
    InMux I__3755 (
            .O(N__27265),
            .I(\ADC_VDC.n20707 ));
    CascadeMux I__3754 (
            .O(N__27262),
            .I(N__27257));
    CascadeMux I__3753 (
            .O(N__27261),
            .I(N__27254));
    InMux I__3752 (
            .O(N__27260),
            .I(N__27251));
    InMux I__3751 (
            .O(N__27257),
            .I(N__27248));
    InMux I__3750 (
            .O(N__27254),
            .I(N__27245));
    LocalMux I__3749 (
            .O(N__27251),
            .I(cmd_rdadctmp_19_adj_1555));
    LocalMux I__3748 (
            .O(N__27248),
            .I(cmd_rdadctmp_19_adj_1555));
    LocalMux I__3747 (
            .O(N__27245),
            .I(cmd_rdadctmp_19_adj_1555));
    InMux I__3746 (
            .O(N__27238),
            .I(N__27235));
    LocalMux I__3745 (
            .O(N__27235),
            .I(N__27231));
    InMux I__3744 (
            .O(N__27234),
            .I(N__27228));
    Odrv4 I__3743 (
            .O(N__27231),
            .I(cmd_rdadcbuf_19));
    LocalMux I__3742 (
            .O(N__27228),
            .I(cmd_rdadcbuf_19));
    InMux I__3741 (
            .O(N__27223),
            .I(\ADC_VDC.n20708 ));
    CascadeMux I__3740 (
            .O(N__27220),
            .I(N__27215));
    InMux I__3739 (
            .O(N__27219),
            .I(N__27210));
    InMux I__3738 (
            .O(N__27218),
            .I(N__27210));
    InMux I__3737 (
            .O(N__27215),
            .I(N__27207));
    LocalMux I__3736 (
            .O(N__27210),
            .I(cmd_rdadctmp_4_adj_1570));
    LocalMux I__3735 (
            .O(N__27207),
            .I(cmd_rdadctmp_4_adj_1570));
    InMux I__3734 (
            .O(N__27202),
            .I(N__27199));
    LocalMux I__3733 (
            .O(N__27199),
            .I(\ADC_VDC.cmd_rdadcbuf_4 ));
    InMux I__3732 (
            .O(N__27196),
            .I(\ADC_VDC.n20693 ));
    CascadeMux I__3731 (
            .O(N__27193),
            .I(N__27189));
    CascadeMux I__3730 (
            .O(N__27192),
            .I(N__27185));
    InMux I__3729 (
            .O(N__27189),
            .I(N__27180));
    InMux I__3728 (
            .O(N__27188),
            .I(N__27180));
    InMux I__3727 (
            .O(N__27185),
            .I(N__27177));
    LocalMux I__3726 (
            .O(N__27180),
            .I(cmd_rdadctmp_5_adj_1569));
    LocalMux I__3725 (
            .O(N__27177),
            .I(cmd_rdadctmp_5_adj_1569));
    InMux I__3724 (
            .O(N__27172),
            .I(N__27169));
    LocalMux I__3723 (
            .O(N__27169),
            .I(N__27166));
    Odrv4 I__3722 (
            .O(N__27166),
            .I(\ADC_VDC.cmd_rdadcbuf_5 ));
    InMux I__3721 (
            .O(N__27163),
            .I(\ADC_VDC.n20694 ));
    CascadeMux I__3720 (
            .O(N__27160),
            .I(N__27155));
    InMux I__3719 (
            .O(N__27159),
            .I(N__27152));
    InMux I__3718 (
            .O(N__27158),
            .I(N__27149));
    InMux I__3717 (
            .O(N__27155),
            .I(N__27146));
    LocalMux I__3716 (
            .O(N__27152),
            .I(cmd_rdadctmp_6_adj_1568));
    LocalMux I__3715 (
            .O(N__27149),
            .I(cmd_rdadctmp_6_adj_1568));
    LocalMux I__3714 (
            .O(N__27146),
            .I(cmd_rdadctmp_6_adj_1568));
    InMux I__3713 (
            .O(N__27139),
            .I(N__27136));
    LocalMux I__3712 (
            .O(N__27136),
            .I(\ADC_VDC.cmd_rdadcbuf_6 ));
    InMux I__3711 (
            .O(N__27133),
            .I(\ADC_VDC.n20695 ));
    CascadeMux I__3710 (
            .O(N__27130),
            .I(N__27125));
    InMux I__3709 (
            .O(N__27129),
            .I(N__27120));
    InMux I__3708 (
            .O(N__27128),
            .I(N__27120));
    InMux I__3707 (
            .O(N__27125),
            .I(N__27117));
    LocalMux I__3706 (
            .O(N__27120),
            .I(cmd_rdadctmp_7_adj_1567));
    LocalMux I__3705 (
            .O(N__27117),
            .I(cmd_rdadctmp_7_adj_1567));
    InMux I__3704 (
            .O(N__27112),
            .I(N__27109));
    LocalMux I__3703 (
            .O(N__27109),
            .I(\ADC_VDC.cmd_rdadcbuf_7 ));
    InMux I__3702 (
            .O(N__27106),
            .I(\ADC_VDC.n20696 ));
    InMux I__3701 (
            .O(N__27103),
            .I(N__27100));
    LocalMux I__3700 (
            .O(N__27100),
            .I(\ADC_VDC.cmd_rdadcbuf_8 ));
    InMux I__3699 (
            .O(N__27097),
            .I(bfn_8_7_0_));
    InMux I__3698 (
            .O(N__27094),
            .I(N__27091));
    LocalMux I__3697 (
            .O(N__27091),
            .I(\ADC_VDC.cmd_rdadcbuf_9 ));
    InMux I__3696 (
            .O(N__27088),
            .I(\ADC_VDC.n20698 ));
    CascadeMux I__3695 (
            .O(N__27085),
            .I(N__27080));
    InMux I__3694 (
            .O(N__27084),
            .I(N__27077));
    InMux I__3693 (
            .O(N__27083),
            .I(N__27074));
    InMux I__3692 (
            .O(N__27080),
            .I(N__27071));
    LocalMux I__3691 (
            .O(N__27077),
            .I(cmd_rdadctmp_10_adj_1564));
    LocalMux I__3690 (
            .O(N__27074),
            .I(cmd_rdadctmp_10_adj_1564));
    LocalMux I__3689 (
            .O(N__27071),
            .I(cmd_rdadctmp_10_adj_1564));
    InMux I__3688 (
            .O(N__27064),
            .I(N__27061));
    LocalMux I__3687 (
            .O(N__27061),
            .I(\ADC_VDC.cmd_rdadcbuf_10 ));
    InMux I__3686 (
            .O(N__27058),
            .I(\ADC_VDC.n20699 ));
    CascadeMux I__3685 (
            .O(N__27055),
            .I(N__27050));
    InMux I__3684 (
            .O(N__27054),
            .I(N__27045));
    InMux I__3683 (
            .O(N__27053),
            .I(N__27045));
    InMux I__3682 (
            .O(N__27050),
            .I(N__27042));
    LocalMux I__3681 (
            .O(N__27045),
            .I(cmd_rdadctmp_11_adj_1563));
    LocalMux I__3680 (
            .O(N__27042),
            .I(cmd_rdadctmp_11_adj_1563));
    InMux I__3679 (
            .O(N__27037),
            .I(\ADC_VDC.n20700 ));
    CascadeMux I__3678 (
            .O(N__27034),
            .I(N__27029));
    InMux I__3677 (
            .O(N__27033),
            .I(N__27026));
    InMux I__3676 (
            .O(N__27032),
            .I(N__27023));
    InMux I__3675 (
            .O(N__27029),
            .I(N__27020));
    LocalMux I__3674 (
            .O(N__27026),
            .I(cmd_rdadctmp_0_adj_1574));
    LocalMux I__3673 (
            .O(N__27023),
            .I(cmd_rdadctmp_0_adj_1574));
    LocalMux I__3672 (
            .O(N__27020),
            .I(cmd_rdadctmp_0_adj_1574));
    InMux I__3671 (
            .O(N__27013),
            .I(N__27010));
    LocalMux I__3670 (
            .O(N__27010),
            .I(\ADC_VDC.cmd_rdadcbuf_0 ));
    CascadeMux I__3669 (
            .O(N__27007),
            .I(N__27002));
    CascadeMux I__3668 (
            .O(N__27006),
            .I(N__26999));
    CascadeMux I__3667 (
            .O(N__27005),
            .I(N__26996));
    InMux I__3666 (
            .O(N__27002),
            .I(N__26991));
    InMux I__3665 (
            .O(N__26999),
            .I(N__26991));
    InMux I__3664 (
            .O(N__26996),
            .I(N__26988));
    LocalMux I__3663 (
            .O(N__26991),
            .I(cmd_rdadctmp_1_adj_1573));
    LocalMux I__3662 (
            .O(N__26988),
            .I(cmd_rdadctmp_1_adj_1573));
    InMux I__3661 (
            .O(N__26983),
            .I(N__26980));
    LocalMux I__3660 (
            .O(N__26980),
            .I(\ADC_VDC.cmd_rdadcbuf_1 ));
    InMux I__3659 (
            .O(N__26977),
            .I(\ADC_VDC.n20690 ));
    CascadeMux I__3658 (
            .O(N__26974),
            .I(N__26971));
    InMux I__3657 (
            .O(N__26971),
            .I(N__26966));
    InMux I__3656 (
            .O(N__26970),
            .I(N__26963));
    InMux I__3655 (
            .O(N__26969),
            .I(N__26960));
    LocalMux I__3654 (
            .O(N__26966),
            .I(N__26957));
    LocalMux I__3653 (
            .O(N__26963),
            .I(cmd_rdadctmp_2_adj_1572));
    LocalMux I__3652 (
            .O(N__26960),
            .I(cmd_rdadctmp_2_adj_1572));
    Odrv4 I__3651 (
            .O(N__26957),
            .I(cmd_rdadctmp_2_adj_1572));
    InMux I__3650 (
            .O(N__26950),
            .I(N__26947));
    LocalMux I__3649 (
            .O(N__26947),
            .I(\ADC_VDC.cmd_rdadcbuf_2 ));
    InMux I__3648 (
            .O(N__26944),
            .I(\ADC_VDC.n20691 ));
    CascadeMux I__3647 (
            .O(N__26941),
            .I(N__26936));
    CascadeMux I__3646 (
            .O(N__26940),
            .I(N__26933));
    CascadeMux I__3645 (
            .O(N__26939),
            .I(N__26930));
    InMux I__3644 (
            .O(N__26936),
            .I(N__26925));
    InMux I__3643 (
            .O(N__26933),
            .I(N__26925));
    InMux I__3642 (
            .O(N__26930),
            .I(N__26922));
    LocalMux I__3641 (
            .O(N__26925),
            .I(cmd_rdadctmp_3_adj_1571));
    LocalMux I__3640 (
            .O(N__26922),
            .I(cmd_rdadctmp_3_adj_1571));
    InMux I__3639 (
            .O(N__26917),
            .I(N__26914));
    LocalMux I__3638 (
            .O(N__26914),
            .I(\ADC_VDC.cmd_rdadcbuf_3 ));
    InMux I__3637 (
            .O(N__26911),
            .I(\ADC_VDC.n20692 ));
    InMux I__3636 (
            .O(N__26908),
            .I(bfn_8_3_0_));
    InMux I__3635 (
            .O(N__26905),
            .I(N__26901));
    InMux I__3634 (
            .O(N__26904),
            .I(N__26898));
    LocalMux I__3633 (
            .O(N__26901),
            .I(\ADC_VDC.avg_cnt_9 ));
    LocalMux I__3632 (
            .O(N__26898),
            .I(\ADC_VDC.avg_cnt_9 ));
    InMux I__3631 (
            .O(N__26893),
            .I(\ADC_VDC.n20733 ));
    InMux I__3630 (
            .O(N__26890),
            .I(\ADC_VDC.n20734 ));
    InMux I__3629 (
            .O(N__26887),
            .I(\ADC_VDC.n20735 ));
    CascadeMux I__3628 (
            .O(N__26884),
            .I(N__26881));
    InMux I__3627 (
            .O(N__26881),
            .I(N__26877));
    InMux I__3626 (
            .O(N__26880),
            .I(N__26874));
    LocalMux I__3625 (
            .O(N__26877),
            .I(N__26871));
    LocalMux I__3624 (
            .O(N__26874),
            .I(\ADC_VDC.avg_cnt_11 ));
    Odrv4 I__3623 (
            .O(N__26871),
            .I(\ADC_VDC.avg_cnt_11 ));
    InMux I__3622 (
            .O(N__26866),
            .I(N__26859));
    CascadeMux I__3621 (
            .O(N__26865),
            .I(N__26849));
    InMux I__3620 (
            .O(N__26864),
            .I(N__26843));
    InMux I__3619 (
            .O(N__26863),
            .I(N__26840));
    InMux I__3618 (
            .O(N__26862),
            .I(N__26834));
    LocalMux I__3617 (
            .O(N__26859),
            .I(N__26831));
    InMux I__3616 (
            .O(N__26858),
            .I(N__26828));
    InMux I__3615 (
            .O(N__26857),
            .I(N__26823));
    InMux I__3614 (
            .O(N__26856),
            .I(N__26823));
    CascadeMux I__3613 (
            .O(N__26855),
            .I(N__26819));
    InMux I__3612 (
            .O(N__26854),
            .I(N__26814));
    InMux I__3611 (
            .O(N__26853),
            .I(N__26805));
    InMux I__3610 (
            .O(N__26852),
            .I(N__26805));
    InMux I__3609 (
            .O(N__26849),
            .I(N__26805));
    InMux I__3608 (
            .O(N__26848),
            .I(N__26805));
    InMux I__3607 (
            .O(N__26847),
            .I(N__26800));
    InMux I__3606 (
            .O(N__26846),
            .I(N__26800));
    LocalMux I__3605 (
            .O(N__26843),
            .I(N__26795));
    LocalMux I__3604 (
            .O(N__26840),
            .I(N__26792));
    CascadeMux I__3603 (
            .O(N__26839),
            .I(N__26787));
    InMux I__3602 (
            .O(N__26838),
            .I(N__26782));
    InMux I__3601 (
            .O(N__26837),
            .I(N__26779));
    LocalMux I__3600 (
            .O(N__26834),
            .I(N__26772));
    Span4Mux_v I__3599 (
            .O(N__26831),
            .I(N__26772));
    LocalMux I__3598 (
            .O(N__26828),
            .I(N__26772));
    LocalMux I__3597 (
            .O(N__26823),
            .I(N__26768));
    InMux I__3596 (
            .O(N__26822),
            .I(N__26765));
    InMux I__3595 (
            .O(N__26819),
            .I(N__26762));
    InMux I__3594 (
            .O(N__26818),
            .I(N__26759));
    InMux I__3593 (
            .O(N__26817),
            .I(N__26756));
    LocalMux I__3592 (
            .O(N__26814),
            .I(N__26749));
    LocalMux I__3591 (
            .O(N__26805),
            .I(N__26749));
    LocalMux I__3590 (
            .O(N__26800),
            .I(N__26749));
    InMux I__3589 (
            .O(N__26799),
            .I(N__26746));
    InMux I__3588 (
            .O(N__26798),
            .I(N__26743));
    Span4Mux_h I__3587 (
            .O(N__26795),
            .I(N__26738));
    Span4Mux_h I__3586 (
            .O(N__26792),
            .I(N__26738));
    InMux I__3585 (
            .O(N__26791),
            .I(N__26733));
    InMux I__3584 (
            .O(N__26790),
            .I(N__26733));
    InMux I__3583 (
            .O(N__26787),
            .I(N__26726));
    InMux I__3582 (
            .O(N__26786),
            .I(N__26726));
    InMux I__3581 (
            .O(N__26785),
            .I(N__26726));
    LocalMux I__3580 (
            .O(N__26782),
            .I(N__26721));
    LocalMux I__3579 (
            .O(N__26779),
            .I(N__26721));
    Span4Mux_h I__3578 (
            .O(N__26772),
            .I(N__26718));
    InMux I__3577 (
            .O(N__26771),
            .I(N__26715));
    Span4Mux_v I__3576 (
            .O(N__26768),
            .I(N__26710));
    LocalMux I__3575 (
            .O(N__26765),
            .I(N__26710));
    LocalMux I__3574 (
            .O(N__26762),
            .I(N__26701));
    LocalMux I__3573 (
            .O(N__26759),
            .I(N__26701));
    LocalMux I__3572 (
            .O(N__26756),
            .I(N__26701));
    Span12Mux_h I__3571 (
            .O(N__26749),
            .I(N__26701));
    LocalMux I__3570 (
            .O(N__26746),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3569 (
            .O(N__26743),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__3568 (
            .O(N__26738),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3567 (
            .O(N__26733),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3566 (
            .O(N__26726),
            .I(\RTD.adc_state_3 ));
    Odrv12 I__3565 (
            .O(N__26721),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__3564 (
            .O(N__26718),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3563 (
            .O(N__26715),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__3562 (
            .O(N__26710),
            .I(\RTD.adc_state_3 ));
    Odrv12 I__3561 (
            .O(N__26701),
            .I(\RTD.adc_state_3 ));
    InMux I__3560 (
            .O(N__26680),
            .I(N__26677));
    LocalMux I__3559 (
            .O(N__26677),
            .I(N__26664));
    InMux I__3558 (
            .O(N__26676),
            .I(N__26661));
    InMux I__3557 (
            .O(N__26675),
            .I(N__26658));
    InMux I__3556 (
            .O(N__26674),
            .I(N__26655));
    CascadeMux I__3555 (
            .O(N__26673),
            .I(N__26647));
    InMux I__3554 (
            .O(N__26672),
            .I(N__26643));
    InMux I__3553 (
            .O(N__26671),
            .I(N__26632));
    InMux I__3552 (
            .O(N__26670),
            .I(N__26632));
    InMux I__3551 (
            .O(N__26669),
            .I(N__26632));
    InMux I__3550 (
            .O(N__26668),
            .I(N__26632));
    InMux I__3549 (
            .O(N__26667),
            .I(N__26632));
    Span4Mux_v I__3548 (
            .O(N__26664),
            .I(N__26625));
    LocalMux I__3547 (
            .O(N__26661),
            .I(N__26625));
    LocalMux I__3546 (
            .O(N__26658),
            .I(N__26625));
    LocalMux I__3545 (
            .O(N__26655),
            .I(N__26622));
    InMux I__3544 (
            .O(N__26654),
            .I(N__26619));
    InMux I__3543 (
            .O(N__26653),
            .I(N__26613));
    InMux I__3542 (
            .O(N__26652),
            .I(N__26610));
    InMux I__3541 (
            .O(N__26651),
            .I(N__26599));
    InMux I__3540 (
            .O(N__26650),
            .I(N__26599));
    InMux I__3539 (
            .O(N__26647),
            .I(N__26594));
    InMux I__3538 (
            .O(N__26646),
            .I(N__26594));
    LocalMux I__3537 (
            .O(N__26643),
            .I(N__26591));
    LocalMux I__3536 (
            .O(N__26632),
            .I(N__26588));
    Span4Mux_v I__3535 (
            .O(N__26625),
            .I(N__26581));
    Span4Mux_h I__3534 (
            .O(N__26622),
            .I(N__26581));
    LocalMux I__3533 (
            .O(N__26619),
            .I(N__26581));
    InMux I__3532 (
            .O(N__26618),
            .I(N__26574));
    InMux I__3531 (
            .O(N__26617),
            .I(N__26574));
    InMux I__3530 (
            .O(N__26616),
            .I(N__26574));
    LocalMux I__3529 (
            .O(N__26613),
            .I(N__26569));
    LocalMux I__3528 (
            .O(N__26610),
            .I(N__26569));
    InMux I__3527 (
            .O(N__26609),
            .I(N__26566));
    InMux I__3526 (
            .O(N__26608),
            .I(N__26561));
    InMux I__3525 (
            .O(N__26607),
            .I(N__26561));
    InMux I__3524 (
            .O(N__26606),
            .I(N__26556));
    InMux I__3523 (
            .O(N__26605),
            .I(N__26556));
    InMux I__3522 (
            .O(N__26604),
            .I(N__26553));
    LocalMux I__3521 (
            .O(N__26599),
            .I(N__26550));
    LocalMux I__3520 (
            .O(N__26594),
            .I(N__26547));
    Span4Mux_v I__3519 (
            .O(N__26591),
            .I(N__26536));
    Span4Mux_h I__3518 (
            .O(N__26588),
            .I(N__26536));
    Span4Mux_h I__3517 (
            .O(N__26581),
            .I(N__26536));
    LocalMux I__3516 (
            .O(N__26574),
            .I(N__26536));
    Span4Mux_h I__3515 (
            .O(N__26569),
            .I(N__26536));
    LocalMux I__3514 (
            .O(N__26566),
            .I(\RTD.adc_state_1 ));
    LocalMux I__3513 (
            .O(N__26561),
            .I(\RTD.adc_state_1 ));
    LocalMux I__3512 (
            .O(N__26556),
            .I(\RTD.adc_state_1 ));
    LocalMux I__3511 (
            .O(N__26553),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__3510 (
            .O(N__26550),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__3509 (
            .O(N__26547),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__3508 (
            .O(N__26536),
            .I(\RTD.adc_state_1 ));
    CascadeMux I__3507 (
            .O(N__26521),
            .I(N__26511));
    CascadeMux I__3506 (
            .O(N__26520),
            .I(N__26507));
    CascadeMux I__3505 (
            .O(N__26519),
            .I(N__26504));
    CascadeMux I__3504 (
            .O(N__26518),
            .I(N__26487));
    CascadeMux I__3503 (
            .O(N__26517),
            .I(N__26483));
    InMux I__3502 (
            .O(N__26516),
            .I(N__26476));
    InMux I__3501 (
            .O(N__26515),
            .I(N__26476));
    InMux I__3500 (
            .O(N__26514),
            .I(N__26476));
    InMux I__3499 (
            .O(N__26511),
            .I(N__26469));
    InMux I__3498 (
            .O(N__26510),
            .I(N__26466));
    InMux I__3497 (
            .O(N__26507),
            .I(N__26463));
    InMux I__3496 (
            .O(N__26504),
            .I(N__26460));
    CascadeMux I__3495 (
            .O(N__26503),
            .I(N__26456));
    InMux I__3494 (
            .O(N__26502),
            .I(N__26441));
    InMux I__3493 (
            .O(N__26501),
            .I(N__26441));
    InMux I__3492 (
            .O(N__26500),
            .I(N__26441));
    InMux I__3491 (
            .O(N__26499),
            .I(N__26441));
    InMux I__3490 (
            .O(N__26498),
            .I(N__26441));
    InMux I__3489 (
            .O(N__26497),
            .I(N__26441));
    InMux I__3488 (
            .O(N__26496),
            .I(N__26441));
    InMux I__3487 (
            .O(N__26495),
            .I(N__26438));
    InMux I__3486 (
            .O(N__26494),
            .I(N__26425));
    InMux I__3485 (
            .O(N__26493),
            .I(N__26425));
    InMux I__3484 (
            .O(N__26492),
            .I(N__26418));
    InMux I__3483 (
            .O(N__26491),
            .I(N__26418));
    InMux I__3482 (
            .O(N__26490),
            .I(N__26418));
    InMux I__3481 (
            .O(N__26487),
            .I(N__26415));
    InMux I__3480 (
            .O(N__26486),
            .I(N__26412));
    InMux I__3479 (
            .O(N__26483),
            .I(N__26409));
    LocalMux I__3478 (
            .O(N__26476),
            .I(N__26406));
    InMux I__3477 (
            .O(N__26475),
            .I(N__26399));
    InMux I__3476 (
            .O(N__26474),
            .I(N__26399));
    InMux I__3475 (
            .O(N__26473),
            .I(N__26399));
    CascadeMux I__3474 (
            .O(N__26472),
            .I(N__26395));
    LocalMux I__3473 (
            .O(N__26469),
            .I(N__26389));
    LocalMux I__3472 (
            .O(N__26466),
            .I(N__26382));
    LocalMux I__3471 (
            .O(N__26463),
            .I(N__26382));
    LocalMux I__3470 (
            .O(N__26460),
            .I(N__26382));
    CascadeMux I__3469 (
            .O(N__26459),
            .I(N__26379));
    InMux I__3468 (
            .O(N__26456),
            .I(N__26376));
    LocalMux I__3467 (
            .O(N__26441),
            .I(N__26367));
    LocalMux I__3466 (
            .O(N__26438),
            .I(N__26367));
    InMux I__3465 (
            .O(N__26437),
            .I(N__26356));
    InMux I__3464 (
            .O(N__26436),
            .I(N__26356));
    InMux I__3463 (
            .O(N__26435),
            .I(N__26356));
    InMux I__3462 (
            .O(N__26434),
            .I(N__26356));
    InMux I__3461 (
            .O(N__26433),
            .I(N__26356));
    InMux I__3460 (
            .O(N__26432),
            .I(N__26349));
    InMux I__3459 (
            .O(N__26431),
            .I(N__26349));
    InMux I__3458 (
            .O(N__26430),
            .I(N__26349));
    LocalMux I__3457 (
            .O(N__26425),
            .I(N__26340));
    LocalMux I__3456 (
            .O(N__26418),
            .I(N__26340));
    LocalMux I__3455 (
            .O(N__26415),
            .I(N__26340));
    LocalMux I__3454 (
            .O(N__26412),
            .I(N__26340));
    LocalMux I__3453 (
            .O(N__26409),
            .I(N__26337));
    Span4Mux_v I__3452 (
            .O(N__26406),
            .I(N__26332));
    LocalMux I__3451 (
            .O(N__26399),
            .I(N__26332));
    CascadeMux I__3450 (
            .O(N__26398),
            .I(N__26329));
    InMux I__3449 (
            .O(N__26395),
            .I(N__26326));
    InMux I__3448 (
            .O(N__26394),
            .I(N__26323));
    InMux I__3447 (
            .O(N__26393),
            .I(N__26318));
    InMux I__3446 (
            .O(N__26392),
            .I(N__26318));
    Span4Mux_v I__3445 (
            .O(N__26389),
            .I(N__26313));
    Span4Mux_v I__3444 (
            .O(N__26382),
            .I(N__26313));
    InMux I__3443 (
            .O(N__26379),
            .I(N__26310));
    LocalMux I__3442 (
            .O(N__26376),
            .I(N__26307));
    InMux I__3441 (
            .O(N__26375),
            .I(N__26298));
    InMux I__3440 (
            .O(N__26374),
            .I(N__26298));
    InMux I__3439 (
            .O(N__26373),
            .I(N__26298));
    InMux I__3438 (
            .O(N__26372),
            .I(N__26298));
    Span12Mux_h I__3437 (
            .O(N__26367),
            .I(N__26291));
    LocalMux I__3436 (
            .O(N__26356),
            .I(N__26291));
    LocalMux I__3435 (
            .O(N__26349),
            .I(N__26291));
    Span4Mux_v I__3434 (
            .O(N__26340),
            .I(N__26284));
    Span4Mux_v I__3433 (
            .O(N__26337),
            .I(N__26284));
    Span4Mux_v I__3432 (
            .O(N__26332),
            .I(N__26284));
    InMux I__3431 (
            .O(N__26329),
            .I(N__26281));
    LocalMux I__3430 (
            .O(N__26326),
            .I(N__26278));
    LocalMux I__3429 (
            .O(N__26323),
            .I(adc_state_2));
    LocalMux I__3428 (
            .O(N__26318),
            .I(adc_state_2));
    Odrv4 I__3427 (
            .O(N__26313),
            .I(adc_state_2));
    LocalMux I__3426 (
            .O(N__26310),
            .I(adc_state_2));
    Odrv12 I__3425 (
            .O(N__26307),
            .I(adc_state_2));
    LocalMux I__3424 (
            .O(N__26298),
            .I(adc_state_2));
    Odrv12 I__3423 (
            .O(N__26291),
            .I(adc_state_2));
    Odrv4 I__3422 (
            .O(N__26284),
            .I(adc_state_2));
    LocalMux I__3421 (
            .O(N__26281),
            .I(adc_state_2));
    Odrv4 I__3420 (
            .O(N__26278),
            .I(adc_state_2));
    CascadeMux I__3419 (
            .O(N__26257),
            .I(N__26254));
    InMux I__3418 (
            .O(N__26254),
            .I(N__26239));
    InMux I__3417 (
            .O(N__26253),
            .I(N__26239));
    InMux I__3416 (
            .O(N__26252),
            .I(N__26239));
    InMux I__3415 (
            .O(N__26251),
            .I(N__26239));
    InMux I__3414 (
            .O(N__26250),
            .I(N__26236));
    InMux I__3413 (
            .O(N__26249),
            .I(N__26230));
    CascadeMux I__3412 (
            .O(N__26248),
            .I(N__26226));
    LocalMux I__3411 (
            .O(N__26239),
            .I(N__26217));
    LocalMux I__3410 (
            .O(N__26236),
            .I(N__26217));
    InMux I__3409 (
            .O(N__26235),
            .I(N__26214));
    InMux I__3408 (
            .O(N__26234),
            .I(N__26210));
    InMux I__3407 (
            .O(N__26233),
            .I(N__26207));
    LocalMux I__3406 (
            .O(N__26230),
            .I(N__26203));
    InMux I__3405 (
            .O(N__26229),
            .I(N__26200));
    InMux I__3404 (
            .O(N__26226),
            .I(N__26197));
    InMux I__3403 (
            .O(N__26225),
            .I(N__26194));
    CascadeMux I__3402 (
            .O(N__26224),
            .I(N__26182));
    InMux I__3401 (
            .O(N__26223),
            .I(N__26178));
    InMux I__3400 (
            .O(N__26222),
            .I(N__26175));
    Span4Mux_h I__3399 (
            .O(N__26217),
            .I(N__26169));
    LocalMux I__3398 (
            .O(N__26214),
            .I(N__26169));
    InMux I__3397 (
            .O(N__26213),
            .I(N__26166));
    LocalMux I__3396 (
            .O(N__26210),
            .I(N__26160));
    LocalMux I__3395 (
            .O(N__26207),
            .I(N__26160));
    InMux I__3394 (
            .O(N__26206),
            .I(N__26157));
    Span4Mux_v I__3393 (
            .O(N__26203),
            .I(N__26152));
    LocalMux I__3392 (
            .O(N__26200),
            .I(N__26152));
    LocalMux I__3391 (
            .O(N__26197),
            .I(N__26147));
    LocalMux I__3390 (
            .O(N__26194),
            .I(N__26147));
    InMux I__3389 (
            .O(N__26193),
            .I(N__26127));
    InMux I__3388 (
            .O(N__26192),
            .I(N__26127));
    InMux I__3387 (
            .O(N__26191),
            .I(N__26127));
    InMux I__3386 (
            .O(N__26190),
            .I(N__26127));
    InMux I__3385 (
            .O(N__26189),
            .I(N__26127));
    InMux I__3384 (
            .O(N__26188),
            .I(N__26127));
    InMux I__3383 (
            .O(N__26187),
            .I(N__26127));
    InMux I__3382 (
            .O(N__26186),
            .I(N__26127));
    InMux I__3381 (
            .O(N__26185),
            .I(N__26124));
    InMux I__3380 (
            .O(N__26182),
            .I(N__26121));
    InMux I__3379 (
            .O(N__26181),
            .I(N__26118));
    LocalMux I__3378 (
            .O(N__26178),
            .I(N__26114));
    LocalMux I__3377 (
            .O(N__26175),
            .I(N__26111));
    InMux I__3376 (
            .O(N__26174),
            .I(N__26108));
    Span4Mux_v I__3375 (
            .O(N__26169),
            .I(N__26103));
    LocalMux I__3374 (
            .O(N__26166),
            .I(N__26103));
    InMux I__3373 (
            .O(N__26165),
            .I(N__26100));
    Span4Mux_h I__3372 (
            .O(N__26160),
            .I(N__26097));
    LocalMux I__3371 (
            .O(N__26157),
            .I(N__26092));
    Span4Mux_h I__3370 (
            .O(N__26152),
            .I(N__26092));
    Span4Mux_v I__3369 (
            .O(N__26147),
            .I(N__26089));
    InMux I__3368 (
            .O(N__26146),
            .I(N__26082));
    InMux I__3367 (
            .O(N__26145),
            .I(N__26082));
    InMux I__3366 (
            .O(N__26144),
            .I(N__26082));
    LocalMux I__3365 (
            .O(N__26127),
            .I(N__26077));
    LocalMux I__3364 (
            .O(N__26124),
            .I(N__26077));
    LocalMux I__3363 (
            .O(N__26121),
            .I(N__26072));
    LocalMux I__3362 (
            .O(N__26118),
            .I(N__26072));
    InMux I__3361 (
            .O(N__26117),
            .I(N__26069));
    Span4Mux_h I__3360 (
            .O(N__26114),
            .I(N__26060));
    Span4Mux_v I__3359 (
            .O(N__26111),
            .I(N__26060));
    LocalMux I__3358 (
            .O(N__26108),
            .I(N__26060));
    Span4Mux_h I__3357 (
            .O(N__26103),
            .I(N__26060));
    LocalMux I__3356 (
            .O(N__26100),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3355 (
            .O(N__26097),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3354 (
            .O(N__26092),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3353 (
            .O(N__26089),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3352 (
            .O(N__26082),
            .I(\RTD.adc_state_0 ));
    Odrv12 I__3351 (
            .O(N__26077),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3350 (
            .O(N__26072),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3349 (
            .O(N__26069),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3348 (
            .O(N__26060),
            .I(\RTD.adc_state_0 ));
    CascadeMux I__3347 (
            .O(N__26041),
            .I(\ADC_VDC.n22071_cascade_ ));
    InMux I__3346 (
            .O(N__26038),
            .I(N__26035));
    LocalMux I__3345 (
            .O(N__26035),
            .I(N__26032));
    Span12Mux_h I__3344 (
            .O(N__26032),
            .I(N__26029));
    Odrv12 I__3343 (
            .O(N__26029),
            .I(EIS_SYNCCLK));
    IoInMux I__3342 (
            .O(N__26026),
            .I(N__26022));
    IoInMux I__3341 (
            .O(N__26025),
            .I(N__26019));
    LocalMux I__3340 (
            .O(N__26022),
            .I(N__26016));
    LocalMux I__3339 (
            .O(N__26019),
            .I(N__26013));
    Span4Mux_s3_h I__3338 (
            .O(N__26016),
            .I(N__26010));
    Span4Mux_s3_v I__3337 (
            .O(N__26013),
            .I(N__26007));
    Span4Mux_h I__3336 (
            .O(N__26010),
            .I(N__26004));
    Span4Mux_h I__3335 (
            .O(N__26007),
            .I(N__26001));
    Span4Mux_h I__3334 (
            .O(N__26004),
            .I(N__25998));
    Sp12to4 I__3333 (
            .O(N__26001),
            .I(N__25993));
    Sp12to4 I__3332 (
            .O(N__25998),
            .I(N__25993));
    Span12Mux_v I__3331 (
            .O(N__25993),
            .I(N__25990));
    Odrv12 I__3330 (
            .O(N__25990),
            .I(IAC_CLK));
    InMux I__3329 (
            .O(N__25987),
            .I(bfn_8_2_0_));
    InMux I__3328 (
            .O(N__25984),
            .I(N__25980));
    InMux I__3327 (
            .O(N__25983),
            .I(N__25977));
    LocalMux I__3326 (
            .O(N__25980),
            .I(\ADC_VDC.avg_cnt_1 ));
    LocalMux I__3325 (
            .O(N__25977),
            .I(\ADC_VDC.avg_cnt_1 ));
    InMux I__3324 (
            .O(N__25972),
            .I(\ADC_VDC.n20725 ));
    CascadeMux I__3323 (
            .O(N__25969),
            .I(N__25965));
    InMux I__3322 (
            .O(N__25968),
            .I(N__25962));
    InMux I__3321 (
            .O(N__25965),
            .I(N__25959));
    LocalMux I__3320 (
            .O(N__25962),
            .I(\ADC_VDC.avg_cnt_2 ));
    LocalMux I__3319 (
            .O(N__25959),
            .I(\ADC_VDC.avg_cnt_2 ));
    InMux I__3318 (
            .O(N__25954),
            .I(\ADC_VDC.n20726 ));
    InMux I__3317 (
            .O(N__25951),
            .I(N__25947));
    InMux I__3316 (
            .O(N__25950),
            .I(N__25944));
    LocalMux I__3315 (
            .O(N__25947),
            .I(\ADC_VDC.avg_cnt_3 ));
    LocalMux I__3314 (
            .O(N__25944),
            .I(\ADC_VDC.avg_cnt_3 ));
    InMux I__3313 (
            .O(N__25939),
            .I(\ADC_VDC.n20727 ));
    InMux I__3312 (
            .O(N__25936),
            .I(N__25932));
    InMux I__3311 (
            .O(N__25935),
            .I(N__25929));
    LocalMux I__3310 (
            .O(N__25932),
            .I(\ADC_VDC.avg_cnt_4 ));
    LocalMux I__3309 (
            .O(N__25929),
            .I(\ADC_VDC.avg_cnt_4 ));
    InMux I__3308 (
            .O(N__25924),
            .I(\ADC_VDC.n20728 ));
    InMux I__3307 (
            .O(N__25921),
            .I(\ADC_VDC.n20729 ));
    InMux I__3306 (
            .O(N__25918),
            .I(N__25914));
    InMux I__3305 (
            .O(N__25917),
            .I(N__25911));
    LocalMux I__3304 (
            .O(N__25914),
            .I(\ADC_VDC.avg_cnt_6 ));
    LocalMux I__3303 (
            .O(N__25911),
            .I(\ADC_VDC.avg_cnt_6 ));
    InMux I__3302 (
            .O(N__25906),
            .I(\ADC_VDC.n20730 ));
    InMux I__3301 (
            .O(N__25903),
            .I(N__25899));
    InMux I__3300 (
            .O(N__25902),
            .I(N__25896));
    LocalMux I__3299 (
            .O(N__25899),
            .I(\ADC_VDC.avg_cnt_7 ));
    LocalMux I__3298 (
            .O(N__25896),
            .I(\ADC_VDC.avg_cnt_7 ));
    InMux I__3297 (
            .O(N__25891),
            .I(\ADC_VDC.n20731 ));
    CascadeMux I__3296 (
            .O(N__25888),
            .I(\ADC_IAC.n22384_cascade_ ));
    CEMux I__3295 (
            .O(N__25885),
            .I(N__25882));
    LocalMux I__3294 (
            .O(N__25882),
            .I(N__25879));
    Odrv4 I__3293 (
            .O(N__25879),
            .I(\ADC_IAC.n22032 ));
    InMux I__3292 (
            .O(N__25876),
            .I(N__25870));
    InMux I__3291 (
            .O(N__25875),
            .I(N__25870));
    LocalMux I__3290 (
            .O(N__25870),
            .I(N__25864));
    InMux I__3289 (
            .O(N__25869),
            .I(N__25859));
    InMux I__3288 (
            .O(N__25868),
            .I(N__25859));
    InMux I__3287 (
            .O(N__25867),
            .I(N__25856));
    Span4Mux_h I__3286 (
            .O(N__25864),
            .I(N__25853));
    LocalMux I__3285 (
            .O(N__25859),
            .I(N__25850));
    LocalMux I__3284 (
            .O(N__25856),
            .I(acadc_trig));
    Odrv4 I__3283 (
            .O(N__25853),
            .I(acadc_trig));
    Odrv4 I__3282 (
            .O(N__25850),
            .I(acadc_trig));
    CascadeMux I__3281 (
            .O(N__25843),
            .I(\ADC_IAC.n17_cascade_ ));
    CEMux I__3280 (
            .O(N__25840),
            .I(N__25837));
    LocalMux I__3279 (
            .O(N__25837),
            .I(N__25834));
    Odrv4 I__3278 (
            .O(N__25834),
            .I(\ADC_IAC.n12 ));
    InMux I__3277 (
            .O(N__25831),
            .I(N__25828));
    LocalMux I__3276 (
            .O(N__25828),
            .I(n21892));
    InMux I__3275 (
            .O(N__25825),
            .I(N__25822));
    LocalMux I__3274 (
            .O(N__25822),
            .I(n14_adj_1578));
    CascadeMux I__3273 (
            .O(N__25819),
            .I(N__25813));
    InMux I__3272 (
            .O(N__25818),
            .I(N__25807));
    InMux I__3271 (
            .O(N__25817),
            .I(N__25807));
    InMux I__3270 (
            .O(N__25816),
            .I(N__25802));
    InMux I__3269 (
            .O(N__25813),
            .I(N__25802));
    InMux I__3268 (
            .O(N__25812),
            .I(N__25799));
    LocalMux I__3267 (
            .O(N__25807),
            .I(N__25796));
    LocalMux I__3266 (
            .O(N__25802),
            .I(N__25793));
    LocalMux I__3265 (
            .O(N__25799),
            .I(N__25790));
    Span4Mux_v I__3264 (
            .O(N__25796),
            .I(N__25787));
    Span4Mux_v I__3263 (
            .O(N__25793),
            .I(N__25782));
    Span4Mux_v I__3262 (
            .O(N__25790),
            .I(N__25782));
    Sp12to4 I__3261 (
            .O(N__25787),
            .I(N__25777));
    Sp12to4 I__3260 (
            .O(N__25782),
            .I(N__25777));
    Span12Mux_h I__3259 (
            .O(N__25777),
            .I(N__25774));
    Odrv12 I__3258 (
            .O(N__25774),
            .I(IAC_DRDY));
    IoInMux I__3257 (
            .O(N__25771),
            .I(N__25768));
    LocalMux I__3256 (
            .O(N__25768),
            .I(N__25765));
    Span12Mux_s8_v I__3255 (
            .O(N__25765),
            .I(N__25761));
    InMux I__3254 (
            .O(N__25764),
            .I(N__25758));
    Odrv12 I__3253 (
            .O(N__25761),
            .I(IAC_CS));
    LocalMux I__3252 (
            .O(N__25758),
            .I(IAC_CS));
    InMux I__3251 (
            .O(N__25753),
            .I(N__25747));
    InMux I__3250 (
            .O(N__25752),
            .I(N__25747));
    LocalMux I__3249 (
            .O(N__25747),
            .I(cmd_rdadctmp_2));
    InMux I__3248 (
            .O(N__25744),
            .I(N__25738));
    InMux I__3247 (
            .O(N__25743),
            .I(N__25738));
    LocalMux I__3246 (
            .O(N__25738),
            .I(cmd_rdadctmp_3));
    CascadeMux I__3245 (
            .O(N__25735),
            .I(N__25731));
    InMux I__3244 (
            .O(N__25734),
            .I(N__25726));
    InMux I__3243 (
            .O(N__25731),
            .I(N__25726));
    LocalMux I__3242 (
            .O(N__25726),
            .I(cmd_rdadctmp_4));
    CascadeMux I__3241 (
            .O(N__25723),
            .I(N__25720));
    InMux I__3240 (
            .O(N__25720),
            .I(N__25716));
    InMux I__3239 (
            .O(N__25719),
            .I(N__25713));
    LocalMux I__3238 (
            .O(N__25716),
            .I(cmd_rdadctmp_0));
    LocalMux I__3237 (
            .O(N__25713),
            .I(cmd_rdadctmp_0));
    CascadeMux I__3236 (
            .O(N__25708),
            .I(N__25705));
    InMux I__3235 (
            .O(N__25705),
            .I(N__25699));
    InMux I__3234 (
            .O(N__25704),
            .I(N__25699));
    LocalMux I__3233 (
            .O(N__25699),
            .I(cmd_rdadctmp_1));
    InMux I__3232 (
            .O(N__25696),
            .I(\ADC_IAC.n20680 ));
    InMux I__3231 (
            .O(N__25693),
            .I(\ADC_IAC.n20681 ));
    InMux I__3230 (
            .O(N__25690),
            .I(\ADC_IAC.n20682 ));
    CEMux I__3229 (
            .O(N__25687),
            .I(N__25684));
    LocalMux I__3228 (
            .O(N__25684),
            .I(N__25681));
    Span4Mux_v I__3227 (
            .O(N__25681),
            .I(N__25678));
    Span4Mux_h I__3226 (
            .O(N__25678),
            .I(N__25674));
    InMux I__3225 (
            .O(N__25677),
            .I(N__25671));
    Odrv4 I__3224 (
            .O(N__25674),
            .I(\ADC_IAC.n13667 ));
    LocalMux I__3223 (
            .O(N__25671),
            .I(\ADC_IAC.n13667 ));
    SRMux I__3222 (
            .O(N__25666),
            .I(N__25663));
    LocalMux I__3221 (
            .O(N__25663),
            .I(N__25660));
    Span4Mux_v I__3220 (
            .O(N__25660),
            .I(N__25657));
    Odrv4 I__3219 (
            .O(N__25657),
            .I(\ADC_IAC.n15622 ));
    InMux I__3218 (
            .O(N__25654),
            .I(N__25651));
    LocalMux I__3217 (
            .O(N__25651),
            .I(\ADC_IAC.n22031 ));
    InMux I__3216 (
            .O(N__25648),
            .I(N__25644));
    InMux I__3215 (
            .O(N__25647),
            .I(N__25641));
    LocalMux I__3214 (
            .O(N__25644),
            .I(\ADC_IAC.bit_cnt_4 ));
    LocalMux I__3213 (
            .O(N__25641),
            .I(\ADC_IAC.bit_cnt_4 ));
    InMux I__3212 (
            .O(N__25636),
            .I(N__25632));
    InMux I__3211 (
            .O(N__25635),
            .I(N__25629));
    LocalMux I__3210 (
            .O(N__25632),
            .I(\ADC_IAC.bit_cnt_3 ));
    LocalMux I__3209 (
            .O(N__25629),
            .I(\ADC_IAC.bit_cnt_3 ));
    CascadeMux I__3208 (
            .O(N__25624),
            .I(N__25620));
    InMux I__3207 (
            .O(N__25623),
            .I(N__25617));
    InMux I__3206 (
            .O(N__25620),
            .I(N__25614));
    LocalMux I__3205 (
            .O(N__25617),
            .I(\ADC_IAC.bit_cnt_1 ));
    LocalMux I__3204 (
            .O(N__25614),
            .I(\ADC_IAC.bit_cnt_1 ));
    InMux I__3203 (
            .O(N__25609),
            .I(N__25605));
    InMux I__3202 (
            .O(N__25608),
            .I(N__25602));
    LocalMux I__3201 (
            .O(N__25605),
            .I(\ADC_IAC.bit_cnt_2 ));
    LocalMux I__3200 (
            .O(N__25602),
            .I(\ADC_IAC.bit_cnt_2 ));
    InMux I__3199 (
            .O(N__25597),
            .I(N__25593));
    InMux I__3198 (
            .O(N__25596),
            .I(N__25590));
    LocalMux I__3197 (
            .O(N__25593),
            .I(\ADC_IAC.bit_cnt_6 ));
    LocalMux I__3196 (
            .O(N__25590),
            .I(\ADC_IAC.bit_cnt_6 ));
    InMux I__3195 (
            .O(N__25585),
            .I(N__25581));
    InMux I__3194 (
            .O(N__25584),
            .I(N__25578));
    LocalMux I__3193 (
            .O(N__25581),
            .I(\ADC_IAC.bit_cnt_0 ));
    LocalMux I__3192 (
            .O(N__25578),
            .I(\ADC_IAC.bit_cnt_0 ));
    CascadeMux I__3191 (
            .O(N__25573),
            .I(\ADC_IAC.n22113_cascade_ ));
    InMux I__3190 (
            .O(N__25570),
            .I(N__25566));
    InMux I__3189 (
            .O(N__25569),
            .I(N__25563));
    LocalMux I__3188 (
            .O(N__25566),
            .I(\ADC_IAC.bit_cnt_7 ));
    LocalMux I__3187 (
            .O(N__25563),
            .I(\ADC_IAC.bit_cnt_7 ));
    InMux I__3186 (
            .O(N__25558),
            .I(N__25554));
    InMux I__3185 (
            .O(N__25557),
            .I(N__25551));
    LocalMux I__3184 (
            .O(N__25554),
            .I(\ADC_IAC.bit_cnt_5 ));
    LocalMux I__3183 (
            .O(N__25551),
            .I(\ADC_IAC.bit_cnt_5 ));
    CascadeMux I__3182 (
            .O(N__25546),
            .I(\ADC_IAC.n22128_cascade_ ));
    InMux I__3181 (
            .O(N__25543),
            .I(N__25540));
    LocalMux I__3180 (
            .O(N__25540),
            .I(N__25537));
    Odrv4 I__3179 (
            .O(N__25537),
            .I(n19));
    CascadeMux I__3178 (
            .O(N__25534),
            .I(N__25531));
    InMux I__3177 (
            .O(N__25531),
            .I(N__25528));
    LocalMux I__3176 (
            .O(N__25528),
            .I(N__25525));
    Span4Mux_v I__3175 (
            .O(N__25525),
            .I(N__25521));
    CascadeMux I__3174 (
            .O(N__25524),
            .I(N__25518));
    Span4Mux_v I__3173 (
            .O(N__25521),
            .I(N__25515));
    InMux I__3172 (
            .O(N__25518),
            .I(N__25512));
    Odrv4 I__3171 (
            .O(N__25515),
            .I(buf_readRTD_0));
    LocalMux I__3170 (
            .O(N__25512),
            .I(buf_readRTD_0));
    CascadeMux I__3169 (
            .O(N__25507),
            .I(n22041_cascade_));
    InMux I__3168 (
            .O(N__25504),
            .I(bfn_7_16_0_));
    InMux I__3167 (
            .O(N__25501),
            .I(\ADC_IAC.n20676 ));
    InMux I__3166 (
            .O(N__25498),
            .I(\ADC_IAC.n20677 ));
    InMux I__3165 (
            .O(N__25495),
            .I(\ADC_IAC.n20678 ));
    InMux I__3164 (
            .O(N__25492),
            .I(\ADC_IAC.n20679 ));
    CascadeMux I__3163 (
            .O(N__25489),
            .I(N__25486));
    InMux I__3162 (
            .O(N__25486),
            .I(N__25483));
    LocalMux I__3161 (
            .O(N__25483),
            .I(n20_adj_1790));
    CascadeMux I__3160 (
            .O(N__25480),
            .I(n23498_cascade_));
    InMux I__3159 (
            .O(N__25477),
            .I(N__25473));
    CascadeMux I__3158 (
            .O(N__25476),
            .I(N__25470));
    LocalMux I__3157 (
            .O(N__25473),
            .I(N__25467));
    InMux I__3156 (
            .O(N__25470),
            .I(N__25464));
    Odrv4 I__3155 (
            .O(N__25467),
            .I(buf_adcdata_vdc_20));
    LocalMux I__3154 (
            .O(N__25464),
            .I(buf_adcdata_vdc_20));
    InMux I__3153 (
            .O(N__25459),
            .I(N__25456));
    LocalMux I__3152 (
            .O(N__25456),
            .I(N__25453));
    Span4Mux_v I__3151 (
            .O(N__25453),
            .I(N__25450));
    Sp12to4 I__3150 (
            .O(N__25450),
            .I(N__25447));
    Span12Mux_h I__3149 (
            .O(N__25447),
            .I(N__25442));
    InMux I__3148 (
            .O(N__25446),
            .I(N__25439));
    InMux I__3147 (
            .O(N__25445),
            .I(N__25436));
    Span12Mux_v I__3146 (
            .O(N__25442),
            .I(N__25433));
    LocalMux I__3145 (
            .O(N__25439),
            .I(N__25428));
    LocalMux I__3144 (
            .O(N__25436),
            .I(N__25428));
    Odrv12 I__3143 (
            .O(N__25433),
            .I(buf_adcdata_vac_20));
    Odrv4 I__3142 (
            .O(N__25428),
            .I(buf_adcdata_vac_20));
    InMux I__3141 (
            .O(N__25423),
            .I(N__25420));
    LocalMux I__3140 (
            .O(N__25420),
            .I(n16_adj_1787));
    InMux I__3139 (
            .O(N__25417),
            .I(N__25414));
    LocalMux I__3138 (
            .O(N__25414),
            .I(n17_adj_1788));
    InMux I__3137 (
            .O(N__25411),
            .I(N__25408));
    LocalMux I__3136 (
            .O(N__25408),
            .I(N__25405));
    Odrv4 I__3135 (
            .O(N__25405),
            .I(n23540));
    InMux I__3134 (
            .O(N__25402),
            .I(N__25399));
    LocalMux I__3133 (
            .O(N__25399),
            .I(N__25396));
    Span12Mux_s9_h I__3132 (
            .O(N__25396),
            .I(N__25393));
    Span12Mux_h I__3131 (
            .O(N__25393),
            .I(N__25389));
    CascadeMux I__3130 (
            .O(N__25392),
            .I(N__25385));
    Span12Mux_v I__3129 (
            .O(N__25389),
            .I(N__25382));
    InMux I__3128 (
            .O(N__25388),
            .I(N__25377));
    InMux I__3127 (
            .O(N__25385),
            .I(N__25377));
    Odrv12 I__3126 (
            .O(N__25382),
            .I(buf_adcdata_iac_23));
    LocalMux I__3125 (
            .O(N__25377),
            .I(buf_adcdata_iac_23));
    CascadeMux I__3124 (
            .O(N__25372),
            .I(N__25368));
    CascadeMux I__3123 (
            .O(N__25371),
            .I(N__25365));
    InMux I__3122 (
            .O(N__25368),
            .I(N__25360));
    InMux I__3121 (
            .O(N__25365),
            .I(N__25360));
    LocalMux I__3120 (
            .O(N__25360),
            .I(cmd_rdadctmp_31));
    InMux I__3119 (
            .O(N__25357),
            .I(N__25351));
    InMux I__3118 (
            .O(N__25356),
            .I(N__25351));
    LocalMux I__3117 (
            .O(N__25351),
            .I(comm_test_buf_24_22));
    InMux I__3116 (
            .O(N__25348),
            .I(N__25344));
    CascadeMux I__3115 (
            .O(N__25347),
            .I(N__25341));
    LocalMux I__3114 (
            .O(N__25344),
            .I(N__25337));
    InMux I__3113 (
            .O(N__25341),
            .I(N__25334));
    InMux I__3112 (
            .O(N__25340),
            .I(N__25331));
    Span4Mux_h I__3111 (
            .O(N__25337),
            .I(N__25328));
    LocalMux I__3110 (
            .O(N__25334),
            .I(buf_dds1_15));
    LocalMux I__3109 (
            .O(N__25331),
            .I(buf_dds1_15));
    Odrv4 I__3108 (
            .O(N__25328),
            .I(buf_dds1_15));
    InMux I__3107 (
            .O(N__25321),
            .I(N__25318));
    LocalMux I__3106 (
            .O(N__25318),
            .I(n111_adj_1771));
    InMux I__3105 (
            .O(N__25315),
            .I(N__25312));
    LocalMux I__3104 (
            .O(N__25312),
            .I(N__25308));
    InMux I__3103 (
            .O(N__25311),
            .I(N__25305));
    Odrv4 I__3102 (
            .O(N__25308),
            .I(buf_adcdata_vdc_8));
    LocalMux I__3101 (
            .O(N__25305),
            .I(buf_adcdata_vdc_8));
    InMux I__3100 (
            .O(N__25300),
            .I(N__25297));
    LocalMux I__3099 (
            .O(N__25297),
            .I(N__25294));
    Span4Mux_v I__3098 (
            .O(N__25294),
            .I(N__25291));
    Sp12to4 I__3097 (
            .O(N__25291),
            .I(N__25287));
    InMux I__3096 (
            .O(N__25290),
            .I(N__25284));
    Span12Mux_h I__3095 (
            .O(N__25287),
            .I(N__25280));
    LocalMux I__3094 (
            .O(N__25284),
            .I(N__25277));
    InMux I__3093 (
            .O(N__25283),
            .I(N__25274));
    Span12Mux_h I__3092 (
            .O(N__25280),
            .I(N__25271));
    Span4Mux_v I__3091 (
            .O(N__25277),
            .I(N__25268));
    LocalMux I__3090 (
            .O(N__25274),
            .I(buf_adcdata_vac_8));
    Odrv12 I__3089 (
            .O(N__25271),
            .I(buf_adcdata_vac_8));
    Odrv4 I__3088 (
            .O(N__25268),
            .I(buf_adcdata_vac_8));
    InMux I__3087 (
            .O(N__25261),
            .I(N__25258));
    LocalMux I__3086 (
            .O(N__25258),
            .I(N__25255));
    Span4Mux_h I__3085 (
            .O(N__25255),
            .I(N__25252));
    Odrv4 I__3084 (
            .O(N__25252),
            .I(n30_adj_1695));
    InMux I__3083 (
            .O(N__25249),
            .I(N__25246));
    LocalMux I__3082 (
            .O(N__25246),
            .I(N__25243));
    Span4Mux_v I__3081 (
            .O(N__25243),
            .I(N__25239));
    CascadeMux I__3080 (
            .O(N__25242),
            .I(N__25236));
    Span4Mux_h I__3079 (
            .O(N__25239),
            .I(N__25233));
    InMux I__3078 (
            .O(N__25236),
            .I(N__25230));
    Odrv4 I__3077 (
            .O(N__25233),
            .I(buf_readRTD_11));
    LocalMux I__3076 (
            .O(N__25230),
            .I(buf_readRTD_11));
    CascadeMux I__3075 (
            .O(N__25225),
            .I(N__25221));
    CascadeMux I__3074 (
            .O(N__25224),
            .I(N__25218));
    InMux I__3073 (
            .O(N__25221),
            .I(N__25212));
    InMux I__3072 (
            .O(N__25218),
            .I(N__25212));
    CascadeMux I__3071 (
            .O(N__25217),
            .I(N__25209));
    LocalMux I__3070 (
            .O(N__25212),
            .I(N__25206));
    InMux I__3069 (
            .O(N__25209),
            .I(N__25203));
    Span4Mux_v I__3068 (
            .O(N__25206),
            .I(N__25198));
    LocalMux I__3067 (
            .O(N__25203),
            .I(N__25198));
    Span4Mux_v I__3066 (
            .O(N__25198),
            .I(N__25193));
    InMux I__3065 (
            .O(N__25197),
            .I(N__25188));
    InMux I__3064 (
            .O(N__25196),
            .I(N__25188));
    Odrv4 I__3063 (
            .O(N__25193),
            .I(buf_cfgRTD_3));
    LocalMux I__3062 (
            .O(N__25188),
            .I(buf_cfgRTD_3));
    InMux I__3061 (
            .O(N__25183),
            .I(N__25180));
    LocalMux I__3060 (
            .O(N__25180),
            .I(N__25176));
    CascadeMux I__3059 (
            .O(N__25179),
            .I(N__25173));
    Span4Mux_h I__3058 (
            .O(N__25176),
            .I(N__25170));
    InMux I__3057 (
            .O(N__25173),
            .I(N__25167));
    Odrv4 I__3056 (
            .O(N__25170),
            .I(buf_adcdata_vdc_6));
    LocalMux I__3055 (
            .O(N__25167),
            .I(buf_adcdata_vdc_6));
    InMux I__3054 (
            .O(N__25162),
            .I(N__25159));
    LocalMux I__3053 (
            .O(N__25159),
            .I(N__25155));
    CascadeMux I__3052 (
            .O(N__25158),
            .I(N__25152));
    Span12Mux_s10_h I__3051 (
            .O(N__25155),
            .I(N__25149));
    InMux I__3050 (
            .O(N__25152),
            .I(N__25146));
    Odrv12 I__3049 (
            .O(N__25149),
            .I(buf_adcdata_vdc_22));
    LocalMux I__3048 (
            .O(N__25146),
            .I(buf_adcdata_vdc_22));
    CascadeMux I__3047 (
            .O(N__25141),
            .I(N__25138));
    InMux I__3046 (
            .O(N__25138),
            .I(N__25134));
    CascadeMux I__3045 (
            .O(N__25137),
            .I(N__25131));
    LocalMux I__3044 (
            .O(N__25134),
            .I(N__25128));
    InMux I__3043 (
            .O(N__25131),
            .I(N__25125));
    Span4Mux_h I__3042 (
            .O(N__25128),
            .I(N__25121));
    LocalMux I__3041 (
            .O(N__25125),
            .I(N__25118));
    InMux I__3040 (
            .O(N__25124),
            .I(N__25115));
    Odrv4 I__3039 (
            .O(N__25121),
            .I(cmd_rdadctmp_26_adj_1522));
    Odrv4 I__3038 (
            .O(N__25118),
            .I(cmd_rdadctmp_26_adj_1522));
    LocalMux I__3037 (
            .O(N__25115),
            .I(cmd_rdadctmp_26_adj_1522));
    CascadeMux I__3036 (
            .O(N__25108),
            .I(n112_adj_1786_cascade_));
    InMux I__3035 (
            .O(N__25105),
            .I(N__25101));
    CascadeMux I__3034 (
            .O(N__25104),
            .I(N__25098));
    LocalMux I__3033 (
            .O(N__25101),
            .I(N__25095));
    InMux I__3032 (
            .O(N__25098),
            .I(N__25092));
    Odrv4 I__3031 (
            .O(N__25095),
            .I(buf_adcdata_vdc_10));
    LocalMux I__3030 (
            .O(N__25092),
            .I(buf_adcdata_vdc_10));
    InMux I__3029 (
            .O(N__25087),
            .I(N__25084));
    LocalMux I__3028 (
            .O(N__25084),
            .I(N__25081));
    Span4Mux_h I__3027 (
            .O(N__25081),
            .I(N__25078));
    Span4Mux_v I__3026 (
            .O(N__25078),
            .I(N__25073));
    InMux I__3025 (
            .O(N__25077),
            .I(N__25070));
    InMux I__3024 (
            .O(N__25076),
            .I(N__25067));
    Sp12to4 I__3023 (
            .O(N__25073),
            .I(N__25064));
    LocalMux I__3022 (
            .O(N__25070),
            .I(N__25059));
    LocalMux I__3021 (
            .O(N__25067),
            .I(N__25059));
    Span12Mux_h I__3020 (
            .O(N__25064),
            .I(N__25056));
    Odrv4 I__3019 (
            .O(N__25059),
            .I(buf_adcdata_vac_10));
    Odrv12 I__3018 (
            .O(N__25056),
            .I(buf_adcdata_vac_10));
    InMux I__3017 (
            .O(N__25051),
            .I(N__25048));
    LocalMux I__3016 (
            .O(N__25048),
            .I(n19_adj_1747));
    InMux I__3015 (
            .O(N__25045),
            .I(N__25041));
    CascadeMux I__3014 (
            .O(N__25044),
            .I(N__25038));
    LocalMux I__3013 (
            .O(N__25041),
            .I(N__25035));
    InMux I__3012 (
            .O(N__25038),
            .I(N__25032));
    Odrv4 I__3011 (
            .O(N__25035),
            .I(buf_adcdata_vdc_15));
    LocalMux I__3010 (
            .O(N__25032),
            .I(buf_adcdata_vdc_15));
    InMux I__3009 (
            .O(N__25027),
            .I(N__25023));
    CascadeMux I__3008 (
            .O(N__25026),
            .I(N__25020));
    LocalMux I__3007 (
            .O(N__25023),
            .I(N__25017));
    InMux I__3006 (
            .O(N__25020),
            .I(N__25014));
    Odrv12 I__3005 (
            .O(N__25017),
            .I(buf_adcdata_vdc_7));
    LocalMux I__3004 (
            .O(N__25014),
            .I(buf_adcdata_vdc_7));
    CascadeMux I__3003 (
            .O(N__25009),
            .I(N__25006));
    InMux I__3002 (
            .O(N__25006),
            .I(N__25003));
    LocalMux I__3001 (
            .O(N__25003),
            .I(N__24999));
    CascadeMux I__3000 (
            .O(N__25002),
            .I(N__24996));
    Span12Mux_v I__2999 (
            .O(N__24999),
            .I(N__24993));
    InMux I__2998 (
            .O(N__24996),
            .I(N__24990));
    Odrv12 I__2997 (
            .O(N__24993),
            .I(buf_adcdata_vdc_23));
    LocalMux I__2996 (
            .O(N__24990),
            .I(buf_adcdata_vdc_23));
    InMux I__2995 (
            .O(N__24985),
            .I(N__24982));
    LocalMux I__2994 (
            .O(N__24982),
            .I(N__24979));
    Span4Mux_v I__2993 (
            .O(N__24979),
            .I(N__24975));
    CascadeMux I__2992 (
            .O(N__24978),
            .I(N__24972));
    Span4Mux_h I__2991 (
            .O(N__24975),
            .I(N__24969));
    InMux I__2990 (
            .O(N__24972),
            .I(N__24966));
    Odrv4 I__2989 (
            .O(N__24969),
            .I(buf_adcdata_vdc_4));
    LocalMux I__2988 (
            .O(N__24966),
            .I(buf_adcdata_vdc_4));
    InMux I__2987 (
            .O(N__24961),
            .I(N__24958));
    LocalMux I__2986 (
            .O(N__24958),
            .I(N__24954));
    InMux I__2985 (
            .O(N__24957),
            .I(N__24951));
    Odrv4 I__2984 (
            .O(N__24954),
            .I(buf_adcdata_vdc_9));
    LocalMux I__2983 (
            .O(N__24951),
            .I(buf_adcdata_vdc_9));
    InMux I__2982 (
            .O(N__24946),
            .I(N__24943));
    LocalMux I__2981 (
            .O(N__24943),
            .I(\RTD.n17 ));
    CascadeMux I__2980 (
            .O(N__24940),
            .I(N__24937));
    InMux I__2979 (
            .O(N__24937),
            .I(N__24934));
    LocalMux I__2978 (
            .O(N__24934),
            .I(N__24930));
    CascadeMux I__2977 (
            .O(N__24933),
            .I(N__24925));
    Span4Mux_h I__2976 (
            .O(N__24930),
            .I(N__24919));
    InMux I__2975 (
            .O(N__24929),
            .I(N__24914));
    InMux I__2974 (
            .O(N__24928),
            .I(N__24914));
    InMux I__2973 (
            .O(N__24925),
            .I(N__24905));
    InMux I__2972 (
            .O(N__24924),
            .I(N__24905));
    InMux I__2971 (
            .O(N__24923),
            .I(N__24905));
    InMux I__2970 (
            .O(N__24922),
            .I(N__24905));
    Span4Mux_v I__2969 (
            .O(N__24919),
            .I(N__24902));
    LocalMux I__2968 (
            .O(N__24914),
            .I(\RTD.n79 ));
    LocalMux I__2967 (
            .O(N__24905),
            .I(\RTD.n79 ));
    Odrv4 I__2966 (
            .O(N__24902),
            .I(\RTD.n79 ));
    CascadeMux I__2965 (
            .O(N__24895),
            .I(N__24892));
    InMux I__2964 (
            .O(N__24892),
            .I(N__24889));
    LocalMux I__2963 (
            .O(N__24889),
            .I(n12356));
    InMux I__2962 (
            .O(N__24886),
            .I(N__24883));
    LocalMux I__2961 (
            .O(N__24883),
            .I(N__24880));
    Odrv4 I__2960 (
            .O(N__24880),
            .I(n22388));
    IoInMux I__2959 (
            .O(N__24877),
            .I(N__24874));
    LocalMux I__2958 (
            .O(N__24874),
            .I(N__24871));
    Span4Mux_s1_h I__2957 (
            .O(N__24871),
            .I(N__24868));
    Span4Mux_h I__2956 (
            .O(N__24868),
            .I(N__24865));
    Span4Mux_h I__2955 (
            .O(N__24865),
            .I(N__24861));
    InMux I__2954 (
            .O(N__24864),
            .I(N__24858));
    Odrv4 I__2953 (
            .O(N__24861),
            .I(VDC_SCLK));
    LocalMux I__2952 (
            .O(N__24858),
            .I(VDC_SCLK));
    CascadeMux I__2951 (
            .O(N__24853),
            .I(n21892_cascade_));
    CascadeMux I__2950 (
            .O(N__24850),
            .I(N__24847));
    InMux I__2949 (
            .O(N__24847),
            .I(N__24844));
    LocalMux I__2948 (
            .O(N__24844),
            .I(N__24841));
    Span4Mux_v I__2947 (
            .O(N__24841),
            .I(N__24838));
    Span4Mux_v I__2946 (
            .O(N__24838),
            .I(N__24835));
    IoSpan4Mux I__2945 (
            .O(N__24835),
            .I(N__24832));
    Odrv4 I__2944 (
            .O(N__24832),
            .I(IAC_MISO));
    IoInMux I__2943 (
            .O(N__24829),
            .I(N__24826));
    LocalMux I__2942 (
            .O(N__24826),
            .I(N__24823));
    Span12Mux_s6_v I__2941 (
            .O(N__24823),
            .I(N__24820));
    Odrv12 I__2940 (
            .O(N__24820),
            .I(GB_BUFFER_DDS_MCLK1_THRU_CO));
    CascadeMux I__2939 (
            .O(N__24817),
            .I(N__24814));
    InMux I__2938 (
            .O(N__24814),
            .I(N__24811));
    LocalMux I__2937 (
            .O(N__24811),
            .I(\CLK_DDS.tmp_buf_0 ));
    CascadeMux I__2936 (
            .O(N__24808),
            .I(N__24805));
    InMux I__2935 (
            .O(N__24805),
            .I(N__24802));
    LocalMux I__2934 (
            .O(N__24802),
            .I(\CLK_DDS.tmp_buf_1 ));
    CascadeMux I__2933 (
            .O(N__24799),
            .I(N__24796));
    InMux I__2932 (
            .O(N__24796),
            .I(N__24793));
    LocalMux I__2931 (
            .O(N__24793),
            .I(\CLK_DDS.tmp_buf_2 ));
    CascadeMux I__2930 (
            .O(N__24790),
            .I(N__24787));
    InMux I__2929 (
            .O(N__24787),
            .I(N__24784));
    LocalMux I__2928 (
            .O(N__24784),
            .I(\CLK_DDS.tmp_buf_3 ));
    CascadeMux I__2927 (
            .O(N__24781),
            .I(N__24778));
    InMux I__2926 (
            .O(N__24778),
            .I(N__24775));
    LocalMux I__2925 (
            .O(N__24775),
            .I(\CLK_DDS.tmp_buf_4 ));
    CascadeMux I__2924 (
            .O(N__24772),
            .I(N__24769));
    InMux I__2923 (
            .O(N__24769),
            .I(N__24766));
    LocalMux I__2922 (
            .O(N__24766),
            .I(\CLK_DDS.tmp_buf_5 ));
    InMux I__2921 (
            .O(N__24763),
            .I(N__24731));
    InMux I__2920 (
            .O(N__24762),
            .I(N__24731));
    InMux I__2919 (
            .O(N__24761),
            .I(N__24731));
    InMux I__2918 (
            .O(N__24760),
            .I(N__24731));
    InMux I__2917 (
            .O(N__24759),
            .I(N__24731));
    InMux I__2916 (
            .O(N__24758),
            .I(N__24731));
    InMux I__2915 (
            .O(N__24757),
            .I(N__24731));
    InMux I__2914 (
            .O(N__24756),
            .I(N__24731));
    InMux I__2913 (
            .O(N__24755),
            .I(N__24714));
    InMux I__2912 (
            .O(N__24754),
            .I(N__24714));
    InMux I__2911 (
            .O(N__24753),
            .I(N__24714));
    InMux I__2910 (
            .O(N__24752),
            .I(N__24714));
    InMux I__2909 (
            .O(N__24751),
            .I(N__24714));
    InMux I__2908 (
            .O(N__24750),
            .I(N__24714));
    InMux I__2907 (
            .O(N__24749),
            .I(N__24714));
    InMux I__2906 (
            .O(N__24748),
            .I(N__24714));
    LocalMux I__2905 (
            .O(N__24731),
            .I(N__24711));
    LocalMux I__2904 (
            .O(N__24714),
            .I(N__24708));
    Span4Mux_v I__2903 (
            .O(N__24711),
            .I(N__24698));
    Span4Mux_v I__2902 (
            .O(N__24708),
            .I(N__24698));
    InMux I__2901 (
            .O(N__24707),
            .I(N__24695));
    InMux I__2900 (
            .O(N__24706),
            .I(N__24692));
    CascadeMux I__2899 (
            .O(N__24705),
            .I(N__24685));
    InMux I__2898 (
            .O(N__24704),
            .I(N__24679));
    InMux I__2897 (
            .O(N__24703),
            .I(N__24679));
    Span4Mux_h I__2896 (
            .O(N__24698),
            .I(N__24672));
    LocalMux I__2895 (
            .O(N__24695),
            .I(N__24672));
    LocalMux I__2894 (
            .O(N__24692),
            .I(N__24672));
    InMux I__2893 (
            .O(N__24691),
            .I(N__24669));
    InMux I__2892 (
            .O(N__24690),
            .I(N__24666));
    InMux I__2891 (
            .O(N__24689),
            .I(N__24663));
    InMux I__2890 (
            .O(N__24688),
            .I(N__24656));
    InMux I__2889 (
            .O(N__24685),
            .I(N__24656));
    InMux I__2888 (
            .O(N__24684),
            .I(N__24656));
    LocalMux I__2887 (
            .O(N__24679),
            .I(N__24647));
    Span4Mux_v I__2886 (
            .O(N__24672),
            .I(N__24647));
    LocalMux I__2885 (
            .O(N__24669),
            .I(N__24647));
    LocalMux I__2884 (
            .O(N__24666),
            .I(N__24647));
    LocalMux I__2883 (
            .O(N__24663),
            .I(dds_state_2_adj_1508));
    LocalMux I__2882 (
            .O(N__24656),
            .I(dds_state_2_adj_1508));
    Odrv4 I__2881 (
            .O(N__24647),
            .I(dds_state_2_adj_1508));
    CEMux I__2880 (
            .O(N__24640),
            .I(N__24636));
    CascadeMux I__2879 (
            .O(N__24639),
            .I(N__24615));
    LocalMux I__2878 (
            .O(N__24636),
            .I(N__24606));
    SRMux I__2877 (
            .O(N__24635),
            .I(N__24603));
    InMux I__2876 (
            .O(N__24634),
            .I(N__24588));
    InMux I__2875 (
            .O(N__24633),
            .I(N__24588));
    InMux I__2874 (
            .O(N__24632),
            .I(N__24588));
    InMux I__2873 (
            .O(N__24631),
            .I(N__24588));
    InMux I__2872 (
            .O(N__24630),
            .I(N__24588));
    InMux I__2871 (
            .O(N__24629),
            .I(N__24588));
    InMux I__2870 (
            .O(N__24628),
            .I(N__24588));
    InMux I__2869 (
            .O(N__24627),
            .I(N__24585));
    InMux I__2868 (
            .O(N__24626),
            .I(N__24568));
    InMux I__2867 (
            .O(N__24625),
            .I(N__24568));
    InMux I__2866 (
            .O(N__24624),
            .I(N__24568));
    InMux I__2865 (
            .O(N__24623),
            .I(N__24568));
    InMux I__2864 (
            .O(N__24622),
            .I(N__24568));
    InMux I__2863 (
            .O(N__24621),
            .I(N__24568));
    InMux I__2862 (
            .O(N__24620),
            .I(N__24568));
    InMux I__2861 (
            .O(N__24619),
            .I(N__24568));
    InMux I__2860 (
            .O(N__24618),
            .I(N__24565));
    InMux I__2859 (
            .O(N__24615),
            .I(N__24560));
    InMux I__2858 (
            .O(N__24614),
            .I(N__24560));
    InMux I__2857 (
            .O(N__24613),
            .I(N__24557));
    InMux I__2856 (
            .O(N__24612),
            .I(N__24550));
    InMux I__2855 (
            .O(N__24611),
            .I(N__24550));
    InMux I__2854 (
            .O(N__24610),
            .I(N__24550));
    CascadeMux I__2853 (
            .O(N__24609),
            .I(N__24547));
    Span4Mux_v I__2852 (
            .O(N__24606),
            .I(N__24543));
    LocalMux I__2851 (
            .O(N__24603),
            .I(N__24540));
    LocalMux I__2850 (
            .O(N__24588),
            .I(N__24537));
    LocalMux I__2849 (
            .O(N__24585),
            .I(N__24530));
    LocalMux I__2848 (
            .O(N__24568),
            .I(N__24530));
    LocalMux I__2847 (
            .O(N__24565),
            .I(N__24530));
    LocalMux I__2846 (
            .O(N__24560),
            .I(N__24523));
    LocalMux I__2845 (
            .O(N__24557),
            .I(N__24523));
    LocalMux I__2844 (
            .O(N__24550),
            .I(N__24523));
    InMux I__2843 (
            .O(N__24547),
            .I(N__24519));
    InMux I__2842 (
            .O(N__24546),
            .I(N__24516));
    Span4Mux_h I__2841 (
            .O(N__24543),
            .I(N__24507));
    Span4Mux_v I__2840 (
            .O(N__24540),
            .I(N__24507));
    Span4Mux_v I__2839 (
            .O(N__24537),
            .I(N__24507));
    Span4Mux_v I__2838 (
            .O(N__24530),
            .I(N__24507));
    Span4Mux_v I__2837 (
            .O(N__24523),
            .I(N__24504));
    InMux I__2836 (
            .O(N__24522),
            .I(N__24501));
    LocalMux I__2835 (
            .O(N__24519),
            .I(N__24496));
    LocalMux I__2834 (
            .O(N__24516),
            .I(N__24496));
    Odrv4 I__2833 (
            .O(N__24507),
            .I(dds_state_1_adj_1509));
    Odrv4 I__2832 (
            .O(N__24504),
            .I(dds_state_1_adj_1509));
    LocalMux I__2831 (
            .O(N__24501),
            .I(dds_state_1_adj_1509));
    Odrv4 I__2830 (
            .O(N__24496),
            .I(dds_state_1_adj_1509));
    CascadeMux I__2829 (
            .O(N__24487),
            .I(N__24484));
    InMux I__2828 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__2827 (
            .O(N__24481),
            .I(\CLK_DDS.tmp_buf_6 ));
    CascadeMux I__2826 (
            .O(N__24478),
            .I(N__24475));
    InMux I__2825 (
            .O(N__24475),
            .I(N__24472));
    LocalMux I__2824 (
            .O(N__24472),
            .I(\CLK_DDS.tmp_buf_7 ));
    CEMux I__2823 (
            .O(N__24469),
            .I(N__24466));
    LocalMux I__2822 (
            .O(N__24466),
            .I(N__24462));
    CEMux I__2821 (
            .O(N__24465),
            .I(N__24459));
    Span4Mux_v I__2820 (
            .O(N__24462),
            .I(N__24456));
    LocalMux I__2819 (
            .O(N__24459),
            .I(N__24453));
    Span4Mux_v I__2818 (
            .O(N__24456),
            .I(N__24450));
    Span4Mux_h I__2817 (
            .O(N__24453),
            .I(N__24447));
    Span4Mux_h I__2816 (
            .O(N__24450),
            .I(N__24442));
    Span4Mux_v I__2815 (
            .O(N__24447),
            .I(N__24442));
    Span4Mux_v I__2814 (
            .O(N__24442),
            .I(N__24439));
    Odrv4 I__2813 (
            .O(N__24439),
            .I(\CLK_DDS.n13376 ));
    InMux I__2812 (
            .O(N__24436),
            .I(N__24433));
    LocalMux I__2811 (
            .O(N__24433),
            .I(n19_adj_1765));
    CascadeMux I__2810 (
            .O(N__24430),
            .I(N__24427));
    InMux I__2809 (
            .O(N__24427),
            .I(N__24424));
    LocalMux I__2808 (
            .O(N__24424),
            .I(N__24421));
    Span12Mux_v I__2807 (
            .O(N__24421),
            .I(N__24418));
    Odrv12 I__2806 (
            .O(N__24418),
            .I(n20_adj_1766));
    CascadeMux I__2805 (
            .O(N__24415),
            .I(N__24412));
    InMux I__2804 (
            .O(N__24412),
            .I(N__24409));
    LocalMux I__2803 (
            .O(N__24409),
            .I(\CLK_DDS.tmp_buf_10 ));
    CascadeMux I__2802 (
            .O(N__24406),
            .I(N__24403));
    InMux I__2801 (
            .O(N__24403),
            .I(N__24400));
    LocalMux I__2800 (
            .O(N__24400),
            .I(\CLK_DDS.tmp_buf_11 ));
    CascadeMux I__2799 (
            .O(N__24397),
            .I(N__24394));
    InMux I__2798 (
            .O(N__24394),
            .I(N__24391));
    LocalMux I__2797 (
            .O(N__24391),
            .I(\CLK_DDS.tmp_buf_12 ));
    CascadeMux I__2796 (
            .O(N__24388),
            .I(N__24385));
    InMux I__2795 (
            .O(N__24385),
            .I(N__24382));
    LocalMux I__2794 (
            .O(N__24382),
            .I(\CLK_DDS.tmp_buf_13 ));
    InMux I__2793 (
            .O(N__24379),
            .I(N__24376));
    LocalMux I__2792 (
            .O(N__24376),
            .I(\CLK_DDS.tmp_buf_14 ));
    CascadeMux I__2791 (
            .O(N__24373),
            .I(N__24370));
    InMux I__2790 (
            .O(N__24370),
            .I(N__24367));
    LocalMux I__2789 (
            .O(N__24367),
            .I(\CLK_DDS.tmp_buf_9 ));
    CascadeMux I__2788 (
            .O(N__24364),
            .I(N__24361));
    InMux I__2787 (
            .O(N__24361),
            .I(N__24358));
    LocalMux I__2786 (
            .O(N__24358),
            .I(\CLK_DDS.tmp_buf_8 ));
    InMux I__2785 (
            .O(N__24355),
            .I(N__24351));
    InMux I__2784 (
            .O(N__24354),
            .I(N__24348));
    LocalMux I__2783 (
            .O(N__24351),
            .I(tmp_buf_15_adj_1511));
    LocalMux I__2782 (
            .O(N__24348),
            .I(tmp_buf_15_adj_1511));
    InMux I__2781 (
            .O(N__24343),
            .I(N__24340));
    LocalMux I__2780 (
            .O(N__24340),
            .I(N__24336));
    CascadeMux I__2779 (
            .O(N__24339),
            .I(N__24333));
    Span4Mux_v I__2778 (
            .O(N__24336),
            .I(N__24330));
    InMux I__2777 (
            .O(N__24333),
            .I(N__24327));
    Odrv4 I__2776 (
            .O(N__24330),
            .I(buf_readRTD_2));
    LocalMux I__2775 (
            .O(N__24327),
            .I(buf_readRTD_2));
    CascadeMux I__2774 (
            .O(N__24322),
            .I(N__24318));
    CascadeMux I__2773 (
            .O(N__24321),
            .I(N__24315));
    InMux I__2772 (
            .O(N__24318),
            .I(N__24312));
    InMux I__2771 (
            .O(N__24315),
            .I(N__24309));
    LocalMux I__2770 (
            .O(N__24312),
            .I(N__24306));
    LocalMux I__2769 (
            .O(N__24309),
            .I(N__24302));
    Span12Mux_s9_h I__2768 (
            .O(N__24306),
            .I(N__24299));
    InMux I__2767 (
            .O(N__24305),
            .I(N__24296));
    Odrv12 I__2766 (
            .O(N__24302),
            .I(cmd_rdadctmp_12_adj_1536));
    Odrv12 I__2765 (
            .O(N__24299),
            .I(cmd_rdadctmp_12_adj_1536));
    LocalMux I__2764 (
            .O(N__24296),
            .I(cmd_rdadctmp_12_adj_1536));
    IoInMux I__2763 (
            .O(N__24289),
            .I(N__24286));
    LocalMux I__2762 (
            .O(N__24286),
            .I(N__24283));
    Span4Mux_s3_v I__2761 (
            .O(N__24283),
            .I(N__24280));
    Span4Mux_v I__2760 (
            .O(N__24280),
            .I(N__24277));
    Span4Mux_v I__2759 (
            .O(N__24277),
            .I(N__24274));
    Span4Mux_v I__2758 (
            .O(N__24274),
            .I(N__24270));
    InMux I__2757 (
            .O(N__24273),
            .I(N__24267));
    Odrv4 I__2756 (
            .O(N__24270),
            .I(DDS_MOSI1));
    LocalMux I__2755 (
            .O(N__24267),
            .I(DDS_MOSI1));
    CascadeMux I__2754 (
            .O(N__24262),
            .I(N__24259));
    InMux I__2753 (
            .O(N__24259),
            .I(N__24255));
    CascadeMux I__2752 (
            .O(N__24258),
            .I(N__24252));
    LocalMux I__2751 (
            .O(N__24255),
            .I(N__24249));
    InMux I__2750 (
            .O(N__24252),
            .I(N__24245));
    Span4Mux_h I__2749 (
            .O(N__24249),
            .I(N__24242));
    InMux I__2748 (
            .O(N__24248),
            .I(N__24239));
    LocalMux I__2747 (
            .O(N__24245),
            .I(cmd_rdadctmp_22_adj_1526));
    Odrv4 I__2746 (
            .O(N__24242),
            .I(cmd_rdadctmp_22_adj_1526));
    LocalMux I__2745 (
            .O(N__24239),
            .I(cmd_rdadctmp_22_adj_1526));
    InMux I__2744 (
            .O(N__24232),
            .I(N__24229));
    LocalMux I__2743 (
            .O(N__24229),
            .I(N__24225));
    CascadeMux I__2742 (
            .O(N__24228),
            .I(N__24222));
    Span4Mux_v I__2741 (
            .O(N__24225),
            .I(N__24219));
    InMux I__2740 (
            .O(N__24222),
            .I(N__24215));
    Sp12to4 I__2739 (
            .O(N__24219),
            .I(N__24212));
    InMux I__2738 (
            .O(N__24218),
            .I(N__24209));
    LocalMux I__2737 (
            .O(N__24215),
            .I(N__24204));
    Span12Mux_h I__2736 (
            .O(N__24212),
            .I(N__24204));
    LocalMux I__2735 (
            .O(N__24209),
            .I(buf_adcdata_vac_15));
    Odrv12 I__2734 (
            .O(N__24204),
            .I(buf_adcdata_vac_15));
    CascadeMux I__2733 (
            .O(N__24199),
            .I(n19_adj_1714_cascade_));
    InMux I__2732 (
            .O(N__24196),
            .I(N__24193));
    LocalMux I__2731 (
            .O(N__24193),
            .I(N__24189));
    InMux I__2730 (
            .O(N__24192),
            .I(N__24186));
    Odrv4 I__2729 (
            .O(N__24189),
            .I(buf_readRTD_7));
    LocalMux I__2728 (
            .O(N__24186),
            .I(buf_readRTD_7));
    CascadeMux I__2727 (
            .O(N__24181),
            .I(N__24177));
    InMux I__2726 (
            .O(N__24180),
            .I(N__24172));
    InMux I__2725 (
            .O(N__24177),
            .I(N__24172));
    LocalMux I__2724 (
            .O(N__24172),
            .I(\RTD.adress_2 ));
    CascadeMux I__2723 (
            .O(N__24169),
            .I(N__24166));
    InMux I__2722 (
            .O(N__24166),
            .I(N__24163));
    LocalMux I__2721 (
            .O(N__24163),
            .I(\RTD.adress_0 ));
    CEMux I__2720 (
            .O(N__24160),
            .I(N__24151));
    InMux I__2719 (
            .O(N__24159),
            .I(N__24138));
    InMux I__2718 (
            .O(N__24158),
            .I(N__24138));
    InMux I__2717 (
            .O(N__24157),
            .I(N__24138));
    InMux I__2716 (
            .O(N__24156),
            .I(N__24138));
    InMux I__2715 (
            .O(N__24155),
            .I(N__24138));
    InMux I__2714 (
            .O(N__24154),
            .I(N__24138));
    LocalMux I__2713 (
            .O(N__24151),
            .I(\RTD.n13441 ));
    LocalMux I__2712 (
            .O(N__24138),
            .I(\RTD.n13441 ));
    CascadeMux I__2711 (
            .O(N__24133),
            .I(N__24129));
    InMux I__2710 (
            .O(N__24132),
            .I(N__24126));
    InMux I__2709 (
            .O(N__24129),
            .I(N__24123));
    LocalMux I__2708 (
            .O(N__24126),
            .I(\RTD.adress_1 ));
    LocalMux I__2707 (
            .O(N__24123),
            .I(\RTD.adress_1 ));
    InMux I__2706 (
            .O(N__24118),
            .I(N__24115));
    LocalMux I__2705 (
            .O(N__24115),
            .I(N__24111));
    CascadeMux I__2704 (
            .O(N__24114),
            .I(N__24108));
    Span4Mux_v I__2703 (
            .O(N__24111),
            .I(N__24104));
    InMux I__2702 (
            .O(N__24108),
            .I(N__24101));
    InMux I__2701 (
            .O(N__24107),
            .I(N__24098));
    Odrv4 I__2700 (
            .O(N__24104),
            .I(read_buf_6));
    LocalMux I__2699 (
            .O(N__24101),
            .I(read_buf_6));
    LocalMux I__2698 (
            .O(N__24098),
            .I(read_buf_6));
    CascadeMux I__2697 (
            .O(N__24091),
            .I(N__24084));
    CascadeMux I__2696 (
            .O(N__24090),
            .I(N__24080));
    InMux I__2695 (
            .O(N__24089),
            .I(N__24073));
    InMux I__2694 (
            .O(N__24088),
            .I(N__24068));
    InMux I__2693 (
            .O(N__24087),
            .I(N__24068));
    InMux I__2692 (
            .O(N__24084),
            .I(N__24062));
    InMux I__2691 (
            .O(N__24083),
            .I(N__24062));
    InMux I__2690 (
            .O(N__24080),
            .I(N__24055));
    InMux I__2689 (
            .O(N__24079),
            .I(N__24055));
    InMux I__2688 (
            .O(N__24078),
            .I(N__24055));
    InMux I__2687 (
            .O(N__24077),
            .I(N__24049));
    InMux I__2686 (
            .O(N__24076),
            .I(N__24046));
    LocalMux I__2685 (
            .O(N__24073),
            .I(N__24041));
    LocalMux I__2684 (
            .O(N__24068),
            .I(N__24041));
    CascadeMux I__2683 (
            .O(N__24067),
            .I(N__24038));
    LocalMux I__2682 (
            .O(N__24062),
            .I(N__24032));
    LocalMux I__2681 (
            .O(N__24055),
            .I(N__24032));
    InMux I__2680 (
            .O(N__24054),
            .I(N__24027));
    InMux I__2679 (
            .O(N__24053),
            .I(N__24027));
    InMux I__2678 (
            .O(N__24052),
            .I(N__24024));
    LocalMux I__2677 (
            .O(N__24049),
            .I(N__24019));
    LocalMux I__2676 (
            .O(N__24046),
            .I(N__24019));
    Span4Mux_v I__2675 (
            .O(N__24041),
            .I(N__24016));
    InMux I__2674 (
            .O(N__24038),
            .I(N__24013));
    InMux I__2673 (
            .O(N__24037),
            .I(N__24010));
    Span4Mux_h I__2672 (
            .O(N__24032),
            .I(N__24007));
    LocalMux I__2671 (
            .O(N__24027),
            .I(N__24004));
    LocalMux I__2670 (
            .O(N__24024),
            .I(N__23999));
    Span4Mux_v I__2669 (
            .O(N__24019),
            .I(N__23999));
    Odrv4 I__2668 (
            .O(N__24016),
            .I(n21989));
    LocalMux I__2667 (
            .O(N__24013),
            .I(n21989));
    LocalMux I__2666 (
            .O(N__24010),
            .I(n21989));
    Odrv4 I__2665 (
            .O(N__24007),
            .I(n21989));
    Odrv12 I__2664 (
            .O(N__24004),
            .I(n21989));
    Odrv4 I__2663 (
            .O(N__23999),
            .I(n21989));
    InMux I__2662 (
            .O(N__23986),
            .I(N__23967));
    InMux I__2661 (
            .O(N__23985),
            .I(N__23967));
    InMux I__2660 (
            .O(N__23984),
            .I(N__23967));
    InMux I__2659 (
            .O(N__23983),
            .I(N__23960));
    InMux I__2658 (
            .O(N__23982),
            .I(N__23960));
    InMux I__2657 (
            .O(N__23981),
            .I(N__23960));
    InMux I__2656 (
            .O(N__23980),
            .I(N__23955));
    InMux I__2655 (
            .O(N__23979),
            .I(N__23955));
    InMux I__2654 (
            .O(N__23978),
            .I(N__23950));
    InMux I__2653 (
            .O(N__23977),
            .I(N__23950));
    InMux I__2652 (
            .O(N__23976),
            .I(N__23945));
    InMux I__2651 (
            .O(N__23975),
            .I(N__23945));
    InMux I__2650 (
            .O(N__23974),
            .I(N__23942));
    LocalMux I__2649 (
            .O(N__23967),
            .I(N__23934));
    LocalMux I__2648 (
            .O(N__23960),
            .I(N__23934));
    LocalMux I__2647 (
            .O(N__23955),
            .I(N__23931));
    LocalMux I__2646 (
            .O(N__23950),
            .I(N__23928));
    LocalMux I__2645 (
            .O(N__23945),
            .I(N__23925));
    LocalMux I__2644 (
            .O(N__23942),
            .I(N__23922));
    InMux I__2643 (
            .O(N__23941),
            .I(N__23915));
    InMux I__2642 (
            .O(N__23940),
            .I(N__23915));
    InMux I__2641 (
            .O(N__23939),
            .I(N__23915));
    Span4Mux_v I__2640 (
            .O(N__23934),
            .I(N__23912));
    Span4Mux_h I__2639 (
            .O(N__23931),
            .I(N__23907));
    Span4Mux_v I__2638 (
            .O(N__23928),
            .I(N__23907));
    Span4Mux_v I__2637 (
            .O(N__23925),
            .I(N__23902));
    Span4Mux_v I__2636 (
            .O(N__23922),
            .I(N__23902));
    LocalMux I__2635 (
            .O(N__23915),
            .I(n13584));
    Odrv4 I__2634 (
            .O(N__23912),
            .I(n13584));
    Odrv4 I__2633 (
            .O(N__23907),
            .I(n13584));
    Odrv4 I__2632 (
            .O(N__23902),
            .I(n13584));
    CascadeMux I__2631 (
            .O(N__23893),
            .I(N__23888));
    InMux I__2630 (
            .O(N__23892),
            .I(N__23881));
    InMux I__2629 (
            .O(N__23891),
            .I(N__23881));
    InMux I__2628 (
            .O(N__23888),
            .I(N__23881));
    LocalMux I__2627 (
            .O(N__23881),
            .I(read_buf_7));
    InMux I__2626 (
            .O(N__23878),
            .I(N__23875));
    LocalMux I__2625 (
            .O(N__23875),
            .I(N__23872));
    Span4Mux_h I__2624 (
            .O(N__23872),
            .I(N__23869));
    Span4Mux_v I__2623 (
            .O(N__23869),
            .I(N__23865));
    CascadeMux I__2622 (
            .O(N__23868),
            .I(N__23862));
    Span4Mux_v I__2621 (
            .O(N__23865),
            .I(N__23858));
    InMux I__2620 (
            .O(N__23862),
            .I(N__23855));
    InMux I__2619 (
            .O(N__23861),
            .I(N__23852));
    Sp12to4 I__2618 (
            .O(N__23858),
            .I(N__23849));
    LocalMux I__2617 (
            .O(N__23855),
            .I(buf_adcdata_vac_9));
    LocalMux I__2616 (
            .O(N__23852),
            .I(buf_adcdata_vac_9));
    Odrv12 I__2615 (
            .O(N__23849),
            .I(buf_adcdata_vac_9));
    InMux I__2614 (
            .O(N__23842),
            .I(N__23839));
    LocalMux I__2613 (
            .O(N__23839),
            .I(n19_adj_1752));
    CascadeMux I__2612 (
            .O(N__23836),
            .I(N__23831));
    InMux I__2611 (
            .O(N__23835),
            .I(N__23828));
    InMux I__2610 (
            .O(N__23834),
            .I(N__23823));
    InMux I__2609 (
            .O(N__23831),
            .I(N__23823));
    LocalMux I__2608 (
            .O(N__23828),
            .I(read_buf_8));
    LocalMux I__2607 (
            .O(N__23823),
            .I(read_buf_8));
    InMux I__2606 (
            .O(N__23818),
            .I(N__23807));
    InMux I__2605 (
            .O(N__23817),
            .I(N__23804));
    InMux I__2604 (
            .O(N__23816),
            .I(N__23799));
    InMux I__2603 (
            .O(N__23815),
            .I(N__23799));
    InMux I__2602 (
            .O(N__23814),
            .I(N__23796));
    CascadeMux I__2601 (
            .O(N__23813),
            .I(N__23793));
    CascadeMux I__2600 (
            .O(N__23812),
            .I(N__23789));
    InMux I__2599 (
            .O(N__23811),
            .I(N__23784));
    InMux I__2598 (
            .O(N__23810),
            .I(N__23784));
    LocalMux I__2597 (
            .O(N__23807),
            .I(N__23772));
    LocalMux I__2596 (
            .O(N__23804),
            .I(N__23772));
    LocalMux I__2595 (
            .O(N__23799),
            .I(N__23772));
    LocalMux I__2594 (
            .O(N__23796),
            .I(N__23769));
    InMux I__2593 (
            .O(N__23793),
            .I(N__23764));
    InMux I__2592 (
            .O(N__23792),
            .I(N__23764));
    InMux I__2591 (
            .O(N__23789),
            .I(N__23761));
    LocalMux I__2590 (
            .O(N__23784),
            .I(N__23758));
    InMux I__2589 (
            .O(N__23783),
            .I(N__23749));
    InMux I__2588 (
            .O(N__23782),
            .I(N__23749));
    InMux I__2587 (
            .O(N__23781),
            .I(N__23749));
    InMux I__2586 (
            .O(N__23780),
            .I(N__23749));
    InMux I__2585 (
            .O(N__23779),
            .I(N__23746));
    Span4Mux_v I__2584 (
            .O(N__23772),
            .I(N__23741));
    Span4Mux_v I__2583 (
            .O(N__23769),
            .I(N__23741));
    LocalMux I__2582 (
            .O(N__23764),
            .I(N__23736));
    LocalMux I__2581 (
            .O(N__23761),
            .I(N__23736));
    Span4Mux_h I__2580 (
            .O(N__23758),
            .I(N__23733));
    LocalMux I__2579 (
            .O(N__23749),
            .I(n13603));
    LocalMux I__2578 (
            .O(N__23746),
            .I(n13603));
    Odrv4 I__2577 (
            .O(N__23741),
            .I(n13603));
    Odrv12 I__2576 (
            .O(N__23736),
            .I(n13603));
    Odrv4 I__2575 (
            .O(N__23733),
            .I(n13603));
    CascadeMux I__2574 (
            .O(N__23722),
            .I(N__23719));
    InMux I__2573 (
            .O(N__23719),
            .I(N__23716));
    LocalMux I__2572 (
            .O(N__23716),
            .I(N__23711));
    CascadeMux I__2571 (
            .O(N__23715),
            .I(N__23708));
    CascadeMux I__2570 (
            .O(N__23714),
            .I(N__23705));
    Span4Mux_h I__2569 (
            .O(N__23711),
            .I(N__23702));
    InMux I__2568 (
            .O(N__23708),
            .I(N__23699));
    InMux I__2567 (
            .O(N__23705),
            .I(N__23696));
    Odrv4 I__2566 (
            .O(N__23702),
            .I(read_buf_9));
    LocalMux I__2565 (
            .O(N__23699),
            .I(read_buf_9));
    LocalMux I__2564 (
            .O(N__23696),
            .I(read_buf_9));
    InMux I__2563 (
            .O(N__23689),
            .I(N__23682));
    InMux I__2562 (
            .O(N__23688),
            .I(N__23679));
    InMux I__2561 (
            .O(N__23687),
            .I(N__23675));
    InMux I__2560 (
            .O(N__23686),
            .I(N__23670));
    InMux I__2559 (
            .O(N__23685),
            .I(N__23670));
    LocalMux I__2558 (
            .O(N__23682),
            .I(N__23667));
    LocalMux I__2557 (
            .O(N__23679),
            .I(N__23664));
    InMux I__2556 (
            .O(N__23678),
            .I(N__23661));
    LocalMux I__2555 (
            .O(N__23675),
            .I(\RTD.adress_7_N_1009_7 ));
    LocalMux I__2554 (
            .O(N__23670),
            .I(\RTD.adress_7_N_1009_7 ));
    Odrv12 I__2553 (
            .O(N__23667),
            .I(\RTD.adress_7_N_1009_7 ));
    Odrv4 I__2552 (
            .O(N__23664),
            .I(\RTD.adress_7_N_1009_7 ));
    LocalMux I__2551 (
            .O(N__23661),
            .I(\RTD.adress_7_N_1009_7 ));
    InMux I__2550 (
            .O(N__23650),
            .I(N__23645));
    InMux I__2549 (
            .O(N__23649),
            .I(N__23640));
    InMux I__2548 (
            .O(N__23648),
            .I(N__23640));
    LocalMux I__2547 (
            .O(N__23645),
            .I(\RTD.n11 ));
    LocalMux I__2546 (
            .O(N__23640),
            .I(\RTD.n11 ));
    CascadeMux I__2545 (
            .O(N__23635),
            .I(\RTD.n11_cascade_ ));
    CEMux I__2544 (
            .O(N__23632),
            .I(N__23629));
    LocalMux I__2543 (
            .O(N__23629),
            .I(N__23626));
    Span4Mux_v I__2542 (
            .O(N__23626),
            .I(N__23623));
    Odrv4 I__2541 (
            .O(N__23623),
            .I(\RTD.n13488 ));
    CascadeMux I__2540 (
            .O(N__23620),
            .I(\RTD.n13488_cascade_ ));
    SRMux I__2539 (
            .O(N__23617),
            .I(N__23614));
    LocalMux I__2538 (
            .O(N__23614),
            .I(N__23611));
    Span4Mux_h I__2537 (
            .O(N__23611),
            .I(N__23608));
    Odrv4 I__2536 (
            .O(N__23608),
            .I(\RTD.n15585 ));
    InMux I__2535 (
            .O(N__23605),
            .I(N__23602));
    LocalMux I__2534 (
            .O(N__23602),
            .I(\RTD.n22081 ));
    CascadeMux I__2533 (
            .O(N__23599),
            .I(N__23595));
    InMux I__2532 (
            .O(N__23598),
            .I(N__23592));
    InMux I__2531 (
            .O(N__23595),
            .I(N__23589));
    LocalMux I__2530 (
            .O(N__23592),
            .I(\RTD.adress_6 ));
    LocalMux I__2529 (
            .O(N__23589),
            .I(\RTD.adress_6 ));
    InMux I__2528 (
            .O(N__23584),
            .I(N__23578));
    InMux I__2527 (
            .O(N__23583),
            .I(N__23578));
    LocalMux I__2526 (
            .O(N__23578),
            .I(\RTD.adress_5 ));
    CascadeMux I__2525 (
            .O(N__23575),
            .I(N__23571));
    InMux I__2524 (
            .O(N__23574),
            .I(N__23566));
    InMux I__2523 (
            .O(N__23571),
            .I(N__23566));
    LocalMux I__2522 (
            .O(N__23566),
            .I(\RTD.adress_4 ));
    InMux I__2521 (
            .O(N__23563),
            .I(N__23557));
    InMux I__2520 (
            .O(N__23562),
            .I(N__23557));
    LocalMux I__2519 (
            .O(N__23557),
            .I(\RTD.adress_3 ));
    InMux I__2518 (
            .O(N__23554),
            .I(N__23548));
    InMux I__2517 (
            .O(N__23553),
            .I(N__23548));
    LocalMux I__2516 (
            .O(N__23548),
            .I(\RTD.cfg_buf_6 ));
    InMux I__2515 (
            .O(N__23545),
            .I(N__23539));
    InMux I__2514 (
            .O(N__23544),
            .I(N__23539));
    LocalMux I__2513 (
            .O(N__23539),
            .I(\RTD.cfg_buf_5 ));
    InMux I__2512 (
            .O(N__23536),
            .I(N__23533));
    LocalMux I__2511 (
            .O(N__23533),
            .I(\RTD.n12 ));
    CascadeMux I__2510 (
            .O(N__23530),
            .I(N__23527));
    InMux I__2509 (
            .O(N__23527),
            .I(N__23523));
    InMux I__2508 (
            .O(N__23526),
            .I(N__23520));
    LocalMux I__2507 (
            .O(N__23523),
            .I(\RTD.cfg_buf_1 ));
    LocalMux I__2506 (
            .O(N__23520),
            .I(\RTD.cfg_buf_1 ));
    InMux I__2505 (
            .O(N__23515),
            .I(N__23512));
    LocalMux I__2504 (
            .O(N__23512),
            .I(\RTD.n20093 ));
    InMux I__2503 (
            .O(N__23509),
            .I(N__23499));
    InMux I__2502 (
            .O(N__23508),
            .I(N__23492));
    InMux I__2501 (
            .O(N__23507),
            .I(N__23492));
    InMux I__2500 (
            .O(N__23506),
            .I(N__23492));
    InMux I__2499 (
            .O(N__23505),
            .I(N__23483));
    InMux I__2498 (
            .O(N__23504),
            .I(N__23483));
    InMux I__2497 (
            .O(N__23503),
            .I(N__23483));
    InMux I__2496 (
            .O(N__23502),
            .I(N__23483));
    LocalMux I__2495 (
            .O(N__23499),
            .I(\RTD.n13482 ));
    LocalMux I__2494 (
            .O(N__23492),
            .I(\RTD.n13482 ));
    LocalMux I__2493 (
            .O(N__23483),
            .I(\RTD.n13482 ));
    CascadeMux I__2492 (
            .O(N__23476),
            .I(N__23471));
    CascadeMux I__2491 (
            .O(N__23475),
            .I(N__23468));
    CascadeMux I__2490 (
            .O(N__23474),
            .I(N__23465));
    InMux I__2489 (
            .O(N__23471),
            .I(N__23455));
    InMux I__2488 (
            .O(N__23468),
            .I(N__23446));
    InMux I__2487 (
            .O(N__23465),
            .I(N__23446));
    InMux I__2486 (
            .O(N__23464),
            .I(N__23446));
    InMux I__2485 (
            .O(N__23463),
            .I(N__23446));
    InMux I__2484 (
            .O(N__23462),
            .I(N__23443));
    InMux I__2483 (
            .O(N__23461),
            .I(N__23436));
    InMux I__2482 (
            .O(N__23460),
            .I(N__23436));
    InMux I__2481 (
            .O(N__23459),
            .I(N__23436));
    InMux I__2480 (
            .O(N__23458),
            .I(N__23433));
    LocalMux I__2479 (
            .O(N__23455),
            .I(N__23428));
    LocalMux I__2478 (
            .O(N__23446),
            .I(N__23428));
    LocalMux I__2477 (
            .O(N__23443),
            .I(N__23425));
    LocalMux I__2476 (
            .O(N__23436),
            .I(\RTD.n68 ));
    LocalMux I__2475 (
            .O(N__23433),
            .I(\RTD.n68 ));
    Odrv4 I__2474 (
            .O(N__23428),
            .I(\RTD.n68 ));
    Odrv4 I__2473 (
            .O(N__23425),
            .I(\RTD.n68 ));
    InMux I__2472 (
            .O(N__23416),
            .I(N__23412));
    InMux I__2471 (
            .O(N__23415),
            .I(N__23409));
    LocalMux I__2470 (
            .O(N__23412),
            .I(\RTD.cfg_buf_7 ));
    LocalMux I__2469 (
            .O(N__23409),
            .I(\RTD.cfg_buf_7 ));
    InMux I__2468 (
            .O(N__23404),
            .I(N__23400));
    CascadeMux I__2467 (
            .O(N__23403),
            .I(N__23397));
    LocalMux I__2466 (
            .O(N__23400),
            .I(N__23394));
    InMux I__2465 (
            .O(N__23397),
            .I(N__23391));
    Odrv4 I__2464 (
            .O(N__23394),
            .I(buf_readRTD_14));
    LocalMux I__2463 (
            .O(N__23391),
            .I(buf_readRTD_14));
    InMux I__2462 (
            .O(N__23386),
            .I(N__23383));
    LocalMux I__2461 (
            .O(N__23383),
            .I(N__23380));
    Odrv4 I__2460 (
            .O(N__23380),
            .I(\RTD.n68_adj_1498 ));
    CEMux I__2459 (
            .O(N__23377),
            .I(N__23374));
    LocalMux I__2458 (
            .O(N__23374),
            .I(N__23371));
    Span4Mux_v I__2457 (
            .O(N__23371),
            .I(N__23368));
    Odrv4 I__2456 (
            .O(N__23368),
            .I(\RTD.n21954 ));
    InMux I__2455 (
            .O(N__23365),
            .I(N__23360));
    InMux I__2454 (
            .O(N__23364),
            .I(N__23357));
    CascadeMux I__2453 (
            .O(N__23363),
            .I(N__23354));
    LocalMux I__2452 (
            .O(N__23360),
            .I(N__23349));
    LocalMux I__2451 (
            .O(N__23357),
            .I(N__23349));
    InMux I__2450 (
            .O(N__23354),
            .I(N__23346));
    Span4Mux_v I__2449 (
            .O(N__23349),
            .I(N__23342));
    LocalMux I__2448 (
            .O(N__23346),
            .I(N__23339));
    InMux I__2447 (
            .O(N__23345),
            .I(N__23336));
    Span4Mux_v I__2446 (
            .O(N__23342),
            .I(N__23333));
    Span4Mux_v I__2445 (
            .O(N__23339),
            .I(N__23328));
    LocalMux I__2444 (
            .O(N__23336),
            .I(N__23328));
    Span4Mux_h I__2443 (
            .O(N__23333),
            .I(N__23325));
    Span4Mux_v I__2442 (
            .O(N__23328),
            .I(N__23322));
    Sp12to4 I__2441 (
            .O(N__23325),
            .I(N__23317));
    Sp12to4 I__2440 (
            .O(N__23322),
            .I(N__23317));
    Odrv12 I__2439 (
            .O(N__23317),
            .I(RTD_DRDY));
    CascadeMux I__2438 (
            .O(N__23314),
            .I(\RTD.n21954_cascade_ ));
    InMux I__2437 (
            .O(N__23311),
            .I(N__23308));
    LocalMux I__2436 (
            .O(N__23308),
            .I(\RTD.n21955 ));
    InMux I__2435 (
            .O(N__23305),
            .I(N__23302));
    LocalMux I__2434 (
            .O(N__23302),
            .I(\RTD.n21988 ));
    CascadeMux I__2433 (
            .O(N__23299),
            .I(\RTD.n7_adj_1497_cascade_ ));
    CascadeMux I__2432 (
            .O(N__23296),
            .I(n13603_cascade_));
    InMux I__2431 (
            .O(N__23293),
            .I(N__23288));
    InMux I__2430 (
            .O(N__23292),
            .I(N__23283));
    InMux I__2429 (
            .O(N__23291),
            .I(N__23283));
    LocalMux I__2428 (
            .O(N__23288),
            .I(read_buf_5));
    LocalMux I__2427 (
            .O(N__23283),
            .I(read_buf_5));
    InMux I__2426 (
            .O(N__23278),
            .I(N__23275));
    LocalMux I__2425 (
            .O(N__23275),
            .I(\RTD.n62 ));
    CEMux I__2424 (
            .O(N__23272),
            .I(N__23268));
    CEMux I__2423 (
            .O(N__23271),
            .I(N__23265));
    LocalMux I__2422 (
            .O(N__23268),
            .I(\RTD.n12274 ));
    LocalMux I__2421 (
            .O(N__23265),
            .I(\RTD.n12274 ));
    InMux I__2420 (
            .O(N__23260),
            .I(N__23257));
    LocalMux I__2419 (
            .O(N__23257),
            .I(\RTD.n11_adj_1500 ));
    InMux I__2418 (
            .O(N__23254),
            .I(N__23251));
    LocalMux I__2417 (
            .O(N__23251),
            .I(N__23247));
    InMux I__2416 (
            .O(N__23250),
            .I(N__23244));
    Span12Mux_s11_h I__2415 (
            .O(N__23247),
            .I(N__23241));
    LocalMux I__2414 (
            .O(N__23244),
            .I(N__23238));
    Span12Mux_v I__2413 (
            .O(N__23241),
            .I(N__23234));
    Span4Mux_v I__2412 (
            .O(N__23238),
            .I(N__23231));
    InMux I__2411 (
            .O(N__23237),
            .I(N__23228));
    Span12Mux_h I__2410 (
            .O(N__23234),
            .I(N__23225));
    Span4Mux_v I__2409 (
            .O(N__23231),
            .I(N__23222));
    LocalMux I__2408 (
            .O(N__23228),
            .I(buf_adcdata_vac_23));
    Odrv12 I__2407 (
            .O(N__23225),
            .I(buf_adcdata_vac_23));
    Odrv4 I__2406 (
            .O(N__23222),
            .I(buf_adcdata_vac_23));
    InMux I__2405 (
            .O(N__23215),
            .I(N__23212));
    LocalMux I__2404 (
            .O(N__23212),
            .I(N__23209));
    Span12Mux_v I__2403 (
            .O(N__23209),
            .I(N__23206));
    Odrv12 I__2402 (
            .O(N__23206),
            .I(n23435));
    InMux I__2401 (
            .O(N__23203),
            .I(N__23197));
    InMux I__2400 (
            .O(N__23202),
            .I(N__23194));
    CascadeMux I__2399 (
            .O(N__23201),
            .I(N__23191));
    InMux I__2398 (
            .O(N__23200),
            .I(N__23188));
    LocalMux I__2397 (
            .O(N__23197),
            .I(N__23185));
    LocalMux I__2396 (
            .O(N__23194),
            .I(N__23182));
    InMux I__2395 (
            .O(N__23191),
            .I(N__23179));
    LocalMux I__2394 (
            .O(N__23188),
            .I(N__23176));
    Span4Mux_h I__2393 (
            .O(N__23185),
            .I(N__23173));
    Span4Mux_v I__2392 (
            .O(N__23182),
            .I(N__23170));
    LocalMux I__2391 (
            .O(N__23179),
            .I(\RTD.mode ));
    Odrv4 I__2390 (
            .O(N__23176),
            .I(\RTD.mode ));
    Odrv4 I__2389 (
            .O(N__23173),
            .I(\RTD.mode ));
    Odrv4 I__2388 (
            .O(N__23170),
            .I(\RTD.mode ));
    InMux I__2387 (
            .O(N__23161),
            .I(N__23155));
    InMux I__2386 (
            .O(N__23160),
            .I(N__23155));
    LocalMux I__2385 (
            .O(N__23155),
            .I(cmd_rdadctmp_31_adj_1517));
    InMux I__2384 (
            .O(N__23152),
            .I(N__23149));
    LocalMux I__2383 (
            .O(N__23149),
            .I(N__23146));
    Span4Mux_v I__2382 (
            .O(N__23146),
            .I(N__23142));
    CascadeMux I__2381 (
            .O(N__23145),
            .I(N__23139));
    Span4Mux_v I__2380 (
            .O(N__23142),
            .I(N__23135));
    InMux I__2379 (
            .O(N__23139),
            .I(N__23130));
    InMux I__2378 (
            .O(N__23138),
            .I(N__23130));
    Odrv4 I__2377 (
            .O(N__23135),
            .I(cmd_rdadctmp_29_adj_1519));
    LocalMux I__2376 (
            .O(N__23130),
            .I(cmd_rdadctmp_29_adj_1519));
    CascadeMux I__2375 (
            .O(N__23125),
            .I(N__23120));
    CascadeMux I__2374 (
            .O(N__23124),
            .I(N__23117));
    InMux I__2373 (
            .O(N__23123),
            .I(N__23110));
    InMux I__2372 (
            .O(N__23120),
            .I(N__23110));
    InMux I__2371 (
            .O(N__23117),
            .I(N__23110));
    LocalMux I__2370 (
            .O(N__23110),
            .I(cmd_rdadctmp_30_adj_1518));
    CascadeMux I__2369 (
            .O(N__23107),
            .I(n21948_cascade_));
    InMux I__2368 (
            .O(N__23104),
            .I(N__23101));
    LocalMux I__2367 (
            .O(N__23101),
            .I(N__23098));
    Span4Mux_h I__2366 (
            .O(N__23098),
            .I(N__23095));
    Sp12to4 I__2365 (
            .O(N__23095),
            .I(N__23092));
    Span12Mux_v I__2364 (
            .O(N__23092),
            .I(N__23088));
    InMux I__2363 (
            .O(N__23091),
            .I(N__23084));
    Span12Mux_h I__2362 (
            .O(N__23088),
            .I(N__23081));
    InMux I__2361 (
            .O(N__23087),
            .I(N__23078));
    LocalMux I__2360 (
            .O(N__23084),
            .I(buf_adcdata_vac_22));
    Odrv12 I__2359 (
            .O(N__23081),
            .I(buf_adcdata_vac_22));
    LocalMux I__2358 (
            .O(N__23078),
            .I(buf_adcdata_vac_22));
    IoInMux I__2357 (
            .O(N__23071),
            .I(N__23068));
    LocalMux I__2356 (
            .O(N__23068),
            .I(N__23065));
    IoSpan4Mux I__2355 (
            .O(N__23065),
            .I(N__23062));
    Span4Mux_s3_v I__2354 (
            .O(N__23062),
            .I(N__23059));
    Span4Mux_v I__2353 (
            .O(N__23059),
            .I(N__23056));
    Odrv4 I__2352 (
            .O(N__23056),
            .I(AC_ADC_SYNC));
    CascadeMux I__2351 (
            .O(N__23053),
            .I(N__23049));
    InMux I__2350 (
            .O(N__23052),
            .I(N__23044));
    InMux I__2349 (
            .O(N__23049),
            .I(N__23044));
    LocalMux I__2348 (
            .O(N__23044),
            .I(N__23041));
    Span4Mux_h I__2347 (
            .O(N__23041),
            .I(N__23037));
    InMux I__2346 (
            .O(N__23040),
            .I(N__23034));
    Odrv4 I__2345 (
            .O(N__23037),
            .I(cmd_rdadctmp_23_adj_1525));
    LocalMux I__2344 (
            .O(N__23034),
            .I(cmd_rdadctmp_23_adj_1525));
    CascadeMux I__2343 (
            .O(N__23029),
            .I(N__23026));
    InMux I__2342 (
            .O(N__23026),
            .I(N__23023));
    LocalMux I__2341 (
            .O(N__23023),
            .I(N__23018));
    InMux I__2340 (
            .O(N__23022),
            .I(N__23013));
    InMux I__2339 (
            .O(N__23021),
            .I(N__23013));
    Odrv4 I__2338 (
            .O(N__23018),
            .I(cmd_rdadctmp_24_adj_1524));
    LocalMux I__2337 (
            .O(N__23013),
            .I(cmd_rdadctmp_24_adj_1524));
    CascadeMux I__2336 (
            .O(N__23008),
            .I(N__23005));
    InMux I__2335 (
            .O(N__23005),
            .I(N__23001));
    CascadeMux I__2334 (
            .O(N__23004),
            .I(N__22998));
    LocalMux I__2333 (
            .O(N__23001),
            .I(N__22995));
    InMux I__2332 (
            .O(N__22998),
            .I(N__22991));
    Span4Mux_h I__2331 (
            .O(N__22995),
            .I(N__22988));
    InMux I__2330 (
            .O(N__22994),
            .I(N__22985));
    LocalMux I__2329 (
            .O(N__22991),
            .I(cmd_rdadctmp_28_adj_1520));
    Odrv4 I__2328 (
            .O(N__22988),
            .I(cmd_rdadctmp_28_adj_1520));
    LocalMux I__2327 (
            .O(N__22985),
            .I(cmd_rdadctmp_28_adj_1520));
    CascadeMux I__2326 (
            .O(N__22978),
            .I(N__22975));
    InMux I__2325 (
            .O(N__22975),
            .I(N__22972));
    LocalMux I__2324 (
            .O(N__22972),
            .I(N__22969));
    Span4Mux_h I__2323 (
            .O(N__22969),
            .I(N__22964));
    InMux I__2322 (
            .O(N__22968),
            .I(N__22959));
    InMux I__2321 (
            .O(N__22967),
            .I(N__22959));
    Odrv4 I__2320 (
            .O(N__22964),
            .I(cmd_rdadctmp_15));
    LocalMux I__2319 (
            .O(N__22959),
            .I(cmd_rdadctmp_15));
    CascadeMux I__2318 (
            .O(N__22954),
            .I(N__22951));
    InMux I__2317 (
            .O(N__22951),
            .I(N__22947));
    CascadeMux I__2316 (
            .O(N__22950),
            .I(N__22944));
    LocalMux I__2315 (
            .O(N__22947),
            .I(N__22940));
    InMux I__2314 (
            .O(N__22944),
            .I(N__22935));
    InMux I__2313 (
            .O(N__22943),
            .I(N__22935));
    Odrv12 I__2312 (
            .O(N__22940),
            .I(cmd_rdadctmp_13_adj_1535));
    LocalMux I__2311 (
            .O(N__22935),
            .I(cmd_rdadctmp_13_adj_1535));
    InMux I__2310 (
            .O(N__22930),
            .I(N__22927));
    LocalMux I__2309 (
            .O(N__22927),
            .I(N__22922));
    InMux I__2308 (
            .O(N__22926),
            .I(N__22919));
    InMux I__2307 (
            .O(N__22925),
            .I(N__22916));
    Span12Mux_v I__2306 (
            .O(N__22922),
            .I(N__22913));
    LocalMux I__2305 (
            .O(N__22919),
            .I(N__22910));
    LocalMux I__2304 (
            .O(N__22916),
            .I(buf_adcdata_vac_5));
    Odrv12 I__2303 (
            .O(N__22913),
            .I(buf_adcdata_vac_5));
    Odrv4 I__2302 (
            .O(N__22910),
            .I(buf_adcdata_vac_5));
    CascadeMux I__2301 (
            .O(N__22903),
            .I(N__22900));
    InMux I__2300 (
            .O(N__22900),
            .I(N__22897));
    LocalMux I__2299 (
            .O(N__22897),
            .I(N__22892));
    InMux I__2298 (
            .O(N__22896),
            .I(N__22887));
    InMux I__2297 (
            .O(N__22895),
            .I(N__22887));
    Odrv4 I__2296 (
            .O(N__22892),
            .I(cmd_rdadctmp_17_adj_1531));
    LocalMux I__2295 (
            .O(N__22887),
            .I(cmd_rdadctmp_17_adj_1531));
    CascadeMux I__2294 (
            .O(N__22882),
            .I(N__22878));
    CascadeMux I__2293 (
            .O(N__22881),
            .I(N__22875));
    InMux I__2292 (
            .O(N__22878),
            .I(N__22870));
    InMux I__2291 (
            .O(N__22875),
            .I(N__22870));
    LocalMux I__2290 (
            .O(N__22870),
            .I(N__22866));
    InMux I__2289 (
            .O(N__22869),
            .I(N__22863));
    Odrv12 I__2288 (
            .O(N__22866),
            .I(cmd_rdadctmp_18_adj_1530));
    LocalMux I__2287 (
            .O(N__22863),
            .I(cmd_rdadctmp_18_adj_1530));
    CascadeMux I__2286 (
            .O(N__22858),
            .I(n23543_cascade_));
    InMux I__2285 (
            .O(N__22855),
            .I(N__22852));
    LocalMux I__2284 (
            .O(N__22852),
            .I(N__22849));
    Odrv4 I__2283 (
            .O(N__22849),
            .I(n19_adj_1696));
    InMux I__2282 (
            .O(N__22846),
            .I(N__22843));
    LocalMux I__2281 (
            .O(N__22843),
            .I(N__22840));
    Span4Mux_v I__2280 (
            .O(N__22840),
            .I(N__22837));
    Odrv4 I__2279 (
            .O(N__22837),
            .I(buf_data_iac_7));
    InMux I__2278 (
            .O(N__22834),
            .I(N__22831));
    LocalMux I__2277 (
            .O(N__22831),
            .I(N__22828));
    Span4Mux_v I__2276 (
            .O(N__22828),
            .I(N__22825));
    Odrv4 I__2275 (
            .O(N__22825),
            .I(n22_adj_1691));
    CascadeMux I__2274 (
            .O(N__22822),
            .I(N__22819));
    InMux I__2273 (
            .O(N__22819),
            .I(N__22815));
    CascadeMux I__2272 (
            .O(N__22818),
            .I(N__22812));
    LocalMux I__2271 (
            .O(N__22815),
            .I(N__22809));
    InMux I__2270 (
            .O(N__22812),
            .I(N__22805));
    Span4Mux_h I__2269 (
            .O(N__22809),
            .I(N__22802));
    InMux I__2268 (
            .O(N__22808),
            .I(N__22799));
    LocalMux I__2267 (
            .O(N__22805),
            .I(cmd_rdadctmp_16_adj_1532));
    Odrv4 I__2266 (
            .O(N__22802),
            .I(cmd_rdadctmp_16_adj_1532));
    LocalMux I__2265 (
            .O(N__22799),
            .I(cmd_rdadctmp_16_adj_1532));
    InMux I__2264 (
            .O(N__22792),
            .I(N__22789));
    LocalMux I__2263 (
            .O(N__22789),
            .I(\RTD.cfg_tmp_3 ));
    InMux I__2262 (
            .O(N__22786),
            .I(N__22783));
    LocalMux I__2261 (
            .O(N__22783),
            .I(\RTD.cfg_tmp_4 ));
    InMux I__2260 (
            .O(N__22780),
            .I(N__22777));
    LocalMux I__2259 (
            .O(N__22777),
            .I(\RTD.cfg_tmp_5 ));
    InMux I__2258 (
            .O(N__22774),
            .I(N__22771));
    LocalMux I__2257 (
            .O(N__22771),
            .I(\RTD.cfg_tmp_6 ));
    CascadeMux I__2256 (
            .O(N__22768),
            .I(N__22765));
    InMux I__2255 (
            .O(N__22765),
            .I(N__22762));
    LocalMux I__2254 (
            .O(N__22762),
            .I(N__22759));
    Span4Mux_v I__2253 (
            .O(N__22759),
            .I(N__22755));
    InMux I__2252 (
            .O(N__22758),
            .I(N__22752));
    Odrv4 I__2251 (
            .O(N__22755),
            .I(\RTD.cfg_tmp_7 ));
    LocalMux I__2250 (
            .O(N__22752),
            .I(\RTD.cfg_tmp_7 ));
    InMux I__2249 (
            .O(N__22747),
            .I(N__22744));
    LocalMux I__2248 (
            .O(N__22744),
            .I(N__22741));
    Span4Mux_v I__2247 (
            .O(N__22741),
            .I(N__22738));
    Odrv4 I__2246 (
            .O(N__22738),
            .I(buf_data_iac_6));
    InMux I__2245 (
            .O(N__22735),
            .I(N__22732));
    LocalMux I__2244 (
            .O(N__22732),
            .I(N__22729));
    Odrv4 I__2243 (
            .O(N__22729),
            .I(n22_adj_1694));
    InMux I__2242 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__2241 (
            .O(N__22723),
            .I(N__22719));
    CascadeMux I__2240 (
            .O(N__22722),
            .I(N__22716));
    Span4Mux_v I__2239 (
            .O(N__22719),
            .I(N__22713));
    InMux I__2238 (
            .O(N__22716),
            .I(N__22710));
    Odrv4 I__2237 (
            .O(N__22713),
            .I(buf_readRTD_1));
    LocalMux I__2236 (
            .O(N__22710),
            .I(buf_readRTD_1));
    InMux I__2235 (
            .O(N__22705),
            .I(N__22702));
    LocalMux I__2234 (
            .O(N__22702),
            .I(N__22699));
    Span4Mux_h I__2233 (
            .O(N__22699),
            .I(N__22695));
    InMux I__2232 (
            .O(N__22698),
            .I(N__22692));
    Odrv4 I__2231 (
            .O(N__22695),
            .I(cmd_rdadctmp_2_adj_1546));
    LocalMux I__2230 (
            .O(N__22692),
            .I(cmd_rdadctmp_2_adj_1546));
    CascadeMux I__2229 (
            .O(N__22687),
            .I(N__22683));
    CascadeMux I__2228 (
            .O(N__22686),
            .I(N__22680));
    InMux I__2227 (
            .O(N__22683),
            .I(N__22677));
    InMux I__2226 (
            .O(N__22680),
            .I(N__22674));
    LocalMux I__2225 (
            .O(N__22677),
            .I(N__22671));
    LocalMux I__2224 (
            .O(N__22674),
            .I(N__22665));
    Span4Mux_v I__2223 (
            .O(N__22671),
            .I(N__22665));
    InMux I__2222 (
            .O(N__22670),
            .I(N__22662));
    Odrv4 I__2221 (
            .O(N__22665),
            .I(cmd_rdadctmp_12));
    LocalMux I__2220 (
            .O(N__22662),
            .I(cmd_rdadctmp_12));
    InMux I__2219 (
            .O(N__22657),
            .I(N__22654));
    LocalMux I__2218 (
            .O(N__22654),
            .I(N__22650));
    CascadeMux I__2217 (
            .O(N__22653),
            .I(N__22647));
    Span4Mux_v I__2216 (
            .O(N__22650),
            .I(N__22644));
    InMux I__2215 (
            .O(N__22647),
            .I(N__22641));
    Span4Mux_h I__2214 (
            .O(N__22644),
            .I(N__22638));
    LocalMux I__2213 (
            .O(N__22641),
            .I(\RTD.adress_7 ));
    Odrv4 I__2212 (
            .O(N__22638),
            .I(\RTD.adress_7 ));
    CascadeMux I__2211 (
            .O(N__22633),
            .I(\RTD.n19_cascade_ ));
    SRMux I__2210 (
            .O(N__22630),
            .I(N__22627));
    LocalMux I__2209 (
            .O(N__22627),
            .I(\RTD.n15396 ));
    InMux I__2208 (
            .O(N__22624),
            .I(N__22621));
    LocalMux I__2207 (
            .O(N__22621),
            .I(\RTD.n1 ));
    CascadeMux I__2206 (
            .O(N__22618),
            .I(\RTD.n1_cascade_ ));
    InMux I__2205 (
            .O(N__22615),
            .I(N__22612));
    LocalMux I__2204 (
            .O(N__22612),
            .I(\RTD.cfg_tmp_0 ));
    CascadeMux I__2203 (
            .O(N__22609),
            .I(N__22606));
    InMux I__2202 (
            .O(N__22606),
            .I(N__22603));
    LocalMux I__2201 (
            .O(N__22603),
            .I(\RTD.cfg_tmp_1 ));
    InMux I__2200 (
            .O(N__22600),
            .I(N__22597));
    LocalMux I__2199 (
            .O(N__22597),
            .I(\RTD.cfg_tmp_2 ));
    CascadeMux I__2198 (
            .O(N__22594),
            .I(\RTD.n68_cascade_ ));
    InMux I__2197 (
            .O(N__22591),
            .I(N__22585));
    InMux I__2196 (
            .O(N__22590),
            .I(N__22585));
    LocalMux I__2195 (
            .O(N__22585),
            .I(\RTD.cfg_buf_4 ));
    InMux I__2194 (
            .O(N__22582),
            .I(N__22576));
    InMux I__2193 (
            .O(N__22581),
            .I(N__22576));
    LocalMux I__2192 (
            .O(N__22576),
            .I(\RTD.cfg_buf_2 ));
    InMux I__2191 (
            .O(N__22573),
            .I(N__22567));
    InMux I__2190 (
            .O(N__22572),
            .I(N__22567));
    LocalMux I__2189 (
            .O(N__22567),
            .I(\RTD.cfg_buf_0 ));
    InMux I__2188 (
            .O(N__22564),
            .I(N__22561));
    LocalMux I__2187 (
            .O(N__22561),
            .I(\RTD.n10 ));
    CascadeMux I__2186 (
            .O(N__22558),
            .I(\RTD.n9_cascade_ ));
    InMux I__2185 (
            .O(N__22555),
            .I(N__22549));
    InMux I__2184 (
            .O(N__22554),
            .I(N__22549));
    LocalMux I__2183 (
            .O(N__22549),
            .I(\RTD.cfg_buf_3 ));
    InMux I__2182 (
            .O(N__22546),
            .I(N__22540));
    InMux I__2181 (
            .O(N__22545),
            .I(N__22540));
    LocalMux I__2180 (
            .O(N__22540),
            .I(\RTD.n20051 ));
    InMux I__2179 (
            .O(N__22537),
            .I(N__22534));
    LocalMux I__2178 (
            .O(N__22534),
            .I(N__22531));
    Span4Mux_h I__2177 (
            .O(N__22531),
            .I(N__22526));
    InMux I__2176 (
            .O(N__22530),
            .I(N__22521));
    InMux I__2175 (
            .O(N__22529),
            .I(N__22521));
    Odrv4 I__2174 (
            .O(N__22526),
            .I(read_buf_0));
    LocalMux I__2173 (
            .O(N__22521),
            .I(read_buf_0));
    InMux I__2172 (
            .O(N__22516),
            .I(N__22512));
    InMux I__2171 (
            .O(N__22515),
            .I(N__22509));
    LocalMux I__2170 (
            .O(N__22512),
            .I(N__22503));
    LocalMux I__2169 (
            .O(N__22509),
            .I(N__22503));
    InMux I__2168 (
            .O(N__22508),
            .I(N__22500));
    Odrv12 I__2167 (
            .O(N__22503),
            .I(\RTD.read_buf_4 ));
    LocalMux I__2166 (
            .O(N__22500),
            .I(\RTD.read_buf_4 ));
    CascadeMux I__2165 (
            .O(N__22495),
            .I(n21989_cascade_));
    InMux I__2164 (
            .O(N__22492),
            .I(N__22486));
    InMux I__2163 (
            .O(N__22491),
            .I(N__22486));
    LocalMux I__2162 (
            .O(N__22486),
            .I(N__22483));
    Span4Mux_h I__2161 (
            .O(N__22483),
            .I(N__22479));
    InMux I__2160 (
            .O(N__22482),
            .I(N__22476));
    Odrv4 I__2159 (
            .O(N__22479),
            .I(read_buf_1));
    LocalMux I__2158 (
            .O(N__22476),
            .I(read_buf_1));
    InMux I__2157 (
            .O(N__22471),
            .I(N__22468));
    LocalMux I__2156 (
            .O(N__22468),
            .I(N__22464));
    CascadeMux I__2155 (
            .O(N__22467),
            .I(N__22460));
    Span4Mux_v I__2154 (
            .O(N__22464),
            .I(N__22457));
    InMux I__2153 (
            .O(N__22463),
            .I(N__22452));
    InMux I__2152 (
            .O(N__22460),
            .I(N__22452));
    Odrv4 I__2151 (
            .O(N__22457),
            .I(read_buf_2));
    LocalMux I__2150 (
            .O(N__22452),
            .I(read_buf_2));
    CascadeMux I__2149 (
            .O(N__22447),
            .I(\RTD.n20051_cascade_ ));
    InMux I__2148 (
            .O(N__22444),
            .I(N__22441));
    LocalMux I__2147 (
            .O(N__22441),
            .I(N__22438));
    Span4Mux_h I__2146 (
            .O(N__22438),
            .I(N__22435));
    Odrv4 I__2145 (
            .O(N__22435),
            .I(\RTD.n22079 ));
    CascadeMux I__2144 (
            .O(N__22432),
            .I(\RTD.n22599_cascade_ ));
    InMux I__2143 (
            .O(N__22429),
            .I(N__22425));
    InMux I__2142 (
            .O(N__22428),
            .I(N__22422));
    LocalMux I__2141 (
            .O(N__22425),
            .I(N__22419));
    LocalMux I__2140 (
            .O(N__22422),
            .I(\RTD.n23689 ));
    Odrv4 I__2139 (
            .O(N__22419),
            .I(\RTD.n23689 ));
    CascadeMux I__2138 (
            .O(N__22414),
            .I(\RTD.n56_cascade_ ));
    InMux I__2137 (
            .O(N__22411),
            .I(N__22408));
    LocalMux I__2136 (
            .O(N__22408),
            .I(N__22405));
    Odrv4 I__2135 (
            .O(N__22405),
            .I(\RTD.n5 ));
    InMux I__2134 (
            .O(N__22402),
            .I(N__22399));
    LocalMux I__2133 (
            .O(N__22399),
            .I(\RTD.n71 ));
    CascadeMux I__2132 (
            .O(N__22396),
            .I(\RTD.n71_cascade_ ));
    InMux I__2131 (
            .O(N__22393),
            .I(N__22390));
    LocalMux I__2130 (
            .O(N__22390),
            .I(\RTD.n22623 ));
    InMux I__2129 (
            .O(N__22387),
            .I(N__22383));
    InMux I__2128 (
            .O(N__22386),
            .I(N__22380));
    LocalMux I__2127 (
            .O(N__22383),
            .I(\ADC_VAC.bit_cnt_6 ));
    LocalMux I__2126 (
            .O(N__22380),
            .I(\ADC_VAC.bit_cnt_6 ));
    InMux I__2125 (
            .O(N__22375),
            .I(N__22371));
    InMux I__2124 (
            .O(N__22374),
            .I(N__22368));
    LocalMux I__2123 (
            .O(N__22371),
            .I(\ADC_VAC.bit_cnt_0 ));
    LocalMux I__2122 (
            .O(N__22368),
            .I(\ADC_VAC.bit_cnt_0 ));
    CascadeMux I__2121 (
            .O(N__22363),
            .I(\ADC_VAC.n22109_cascade_ ));
    InMux I__2120 (
            .O(N__22360),
            .I(N__22356));
    InMux I__2119 (
            .O(N__22359),
            .I(N__22353));
    LocalMux I__2118 (
            .O(N__22356),
            .I(\ADC_VAC.bit_cnt_7 ));
    LocalMux I__2117 (
            .O(N__22353),
            .I(\ADC_VAC.bit_cnt_7 ));
    CascadeMux I__2116 (
            .O(N__22348),
            .I(\ADC_VAC.n22126_cascade_ ));
    InMux I__2115 (
            .O(N__22345),
            .I(N__22341));
    InMux I__2114 (
            .O(N__22344),
            .I(N__22338));
    LocalMux I__2113 (
            .O(N__22341),
            .I(\ADC_VAC.bit_cnt_5 ));
    LocalMux I__2112 (
            .O(N__22338),
            .I(\ADC_VAC.bit_cnt_5 ));
    CascadeMux I__2111 (
            .O(N__22333),
            .I(\ADC_VAC.n22389_cascade_ ));
    CEMux I__2110 (
            .O(N__22330),
            .I(N__22327));
    LocalMux I__2109 (
            .O(N__22327),
            .I(N__22324));
    Odrv4 I__2108 (
            .O(N__22324),
            .I(\ADC_VAC.n22030 ));
    InMux I__2107 (
            .O(N__22321),
            .I(N__22318));
    LocalMux I__2106 (
            .O(N__22318),
            .I(\ADC_VAC.n17 ));
    CascadeMux I__2105 (
            .O(N__22315),
            .I(N__22312));
    InMux I__2104 (
            .O(N__22312),
            .I(N__22307));
    InMux I__2103 (
            .O(N__22311),
            .I(N__22304));
    InMux I__2102 (
            .O(N__22310),
            .I(N__22301));
    LocalMux I__2101 (
            .O(N__22307),
            .I(N__22296));
    LocalMux I__2100 (
            .O(N__22304),
            .I(N__22296));
    LocalMux I__2099 (
            .O(N__22301),
            .I(N__22291));
    Span4Mux_v I__2098 (
            .O(N__22296),
            .I(N__22288));
    InMux I__2097 (
            .O(N__22295),
            .I(N__22283));
    InMux I__2096 (
            .O(N__22294),
            .I(N__22283));
    Span4Mux_v I__2095 (
            .O(N__22291),
            .I(N__22280));
    Sp12to4 I__2094 (
            .O(N__22288),
            .I(N__22275));
    LocalMux I__2093 (
            .O(N__22283),
            .I(N__22275));
    Span4Mux_h I__2092 (
            .O(N__22280),
            .I(N__22272));
    Odrv12 I__2091 (
            .O(N__22275),
            .I(VAC_DRDY));
    Odrv4 I__2090 (
            .O(N__22272),
            .I(VAC_DRDY));
    CEMux I__2089 (
            .O(N__22267),
            .I(N__22263));
    CEMux I__2088 (
            .O(N__22266),
            .I(N__22260));
    LocalMux I__2087 (
            .O(N__22263),
            .I(N__22257));
    LocalMux I__2086 (
            .O(N__22260),
            .I(N__22254));
    Span4Mux_h I__2085 (
            .O(N__22257),
            .I(N__22251));
    Span4Mux_v I__2084 (
            .O(N__22254),
            .I(N__22248));
    Odrv4 I__2083 (
            .O(N__22251),
            .I(\ADC_VAC.n12 ));
    Odrv4 I__2082 (
            .O(N__22248),
            .I(\ADC_VAC.n12 ));
    IoInMux I__2081 (
            .O(N__22243),
            .I(N__22240));
    LocalMux I__2080 (
            .O(N__22240),
            .I(N__22237));
    Span12Mux_s8_h I__2079 (
            .O(N__22237),
            .I(N__22234));
    Odrv12 I__2078 (
            .O(N__22234),
            .I(RTD_CS));
    InMux I__2077 (
            .O(N__22231),
            .I(N__22228));
    LocalMux I__2076 (
            .O(N__22228),
            .I(\RTD.n22382 ));
    InMux I__2075 (
            .O(N__22225),
            .I(N__22222));
    LocalMux I__2074 (
            .O(N__22222),
            .I(n22_adj_1697));
    CascadeMux I__2073 (
            .O(N__22219),
            .I(N__22216));
    InMux I__2072 (
            .O(N__22216),
            .I(N__22213));
    LocalMux I__2071 (
            .O(N__22213),
            .I(N__22209));
    CascadeMux I__2070 (
            .O(N__22212),
            .I(N__22206));
    Span4Mux_h I__2069 (
            .O(N__22209),
            .I(N__22202));
    InMux I__2068 (
            .O(N__22206),
            .I(N__22199));
    InMux I__2067 (
            .O(N__22205),
            .I(N__22196));
    Odrv4 I__2066 (
            .O(N__22202),
            .I(cmd_rdadctmp_15_adj_1533));
    LocalMux I__2065 (
            .O(N__22199),
            .I(cmd_rdadctmp_15_adj_1533));
    LocalMux I__2064 (
            .O(N__22196),
            .I(cmd_rdadctmp_15_adj_1533));
    CascadeMux I__2063 (
            .O(N__22189),
            .I(N__22186));
    InMux I__2062 (
            .O(N__22186),
            .I(N__22182));
    CascadeMux I__2061 (
            .O(N__22185),
            .I(N__22179));
    LocalMux I__2060 (
            .O(N__22182),
            .I(N__22175));
    InMux I__2059 (
            .O(N__22179),
            .I(N__22170));
    InMux I__2058 (
            .O(N__22178),
            .I(N__22170));
    Odrv4 I__2057 (
            .O(N__22175),
            .I(cmd_rdadctmp_13));
    LocalMux I__2056 (
            .O(N__22170),
            .I(cmd_rdadctmp_13));
    InMux I__2055 (
            .O(N__22165),
            .I(N__22162));
    LocalMux I__2054 (
            .O(N__22162),
            .I(N__22158));
    InMux I__2053 (
            .O(N__22161),
            .I(N__22154));
    Span4Mux_v I__2052 (
            .O(N__22158),
            .I(N__22151));
    InMux I__2051 (
            .O(N__22157),
            .I(N__22148));
    LocalMux I__2050 (
            .O(N__22154),
            .I(buf_adcdata_iac_5));
    Odrv4 I__2049 (
            .O(N__22151),
            .I(buf_adcdata_iac_5));
    LocalMux I__2048 (
            .O(N__22148),
            .I(buf_adcdata_iac_5));
    CascadeMux I__2047 (
            .O(N__22141),
            .I(\ADC_VAC.n13747_cascade_ ));
    InMux I__2046 (
            .O(N__22138),
            .I(N__22135));
    LocalMux I__2045 (
            .O(N__22135),
            .I(\ADC_VAC.n13842 ));
    InMux I__2044 (
            .O(N__22132),
            .I(N__22128));
    InMux I__2043 (
            .O(N__22131),
            .I(N__22125));
    LocalMux I__2042 (
            .O(N__22128),
            .I(\ADC_VAC.bit_cnt_2 ));
    LocalMux I__2041 (
            .O(N__22125),
            .I(\ADC_VAC.bit_cnt_2 ));
    InMux I__2040 (
            .O(N__22120),
            .I(N__22116));
    InMux I__2039 (
            .O(N__22119),
            .I(N__22113));
    LocalMux I__2038 (
            .O(N__22116),
            .I(\ADC_VAC.bit_cnt_1 ));
    LocalMux I__2037 (
            .O(N__22113),
            .I(\ADC_VAC.bit_cnt_1 ));
    CascadeMux I__2036 (
            .O(N__22108),
            .I(N__22104));
    InMux I__2035 (
            .O(N__22107),
            .I(N__22101));
    InMux I__2034 (
            .O(N__22104),
            .I(N__22098));
    LocalMux I__2033 (
            .O(N__22101),
            .I(\ADC_VAC.bit_cnt_3 ));
    LocalMux I__2032 (
            .O(N__22098),
            .I(\ADC_VAC.bit_cnt_3 ));
    InMux I__2031 (
            .O(N__22093),
            .I(N__22089));
    InMux I__2030 (
            .O(N__22092),
            .I(N__22086));
    LocalMux I__2029 (
            .O(N__22089),
            .I(\ADC_VAC.bit_cnt_4 ));
    LocalMux I__2028 (
            .O(N__22086),
            .I(\ADC_VAC.bit_cnt_4 ));
    InMux I__2027 (
            .O(N__22081),
            .I(N__22078));
    LocalMux I__2026 (
            .O(N__22078),
            .I(N__22075));
    Span4Mux_h I__2025 (
            .O(N__22075),
            .I(N__22072));
    Odrv4 I__2024 (
            .O(N__22072),
            .I(buf_data_iac_5));
    InMux I__2023 (
            .O(N__22069),
            .I(N__22066));
    LocalMux I__2022 (
            .O(N__22066),
            .I(N__22063));
    Span4Mux_h I__2021 (
            .O(N__22063),
            .I(N__22058));
    InMux I__2020 (
            .O(N__22062),
            .I(N__22053));
    InMux I__2019 (
            .O(N__22061),
            .I(N__22053));
    Odrv4 I__2018 (
            .O(N__22058),
            .I(buf_adcdata_iac_6));
    LocalMux I__2017 (
            .O(N__22053),
            .I(buf_adcdata_iac_6));
    InMux I__2016 (
            .O(N__22048),
            .I(N__22045));
    LocalMux I__2015 (
            .O(N__22045),
            .I(N__22041));
    InMux I__2014 (
            .O(N__22044),
            .I(N__22037));
    Span4Mux_v I__2013 (
            .O(N__22041),
            .I(N__22034));
    InMux I__2012 (
            .O(N__22040),
            .I(N__22031));
    LocalMux I__2011 (
            .O(N__22037),
            .I(buf_adcdata_iac_7));
    Odrv4 I__2010 (
            .O(N__22034),
            .I(buf_adcdata_iac_7));
    LocalMux I__2009 (
            .O(N__22031),
            .I(buf_adcdata_iac_7));
    CascadeMux I__2008 (
            .O(N__22024),
            .I(N__22021));
    InMux I__2007 (
            .O(N__22021),
            .I(N__22012));
    InMux I__2006 (
            .O(N__22020),
            .I(N__22012));
    InMux I__2005 (
            .O(N__22019),
            .I(N__22012));
    LocalMux I__2004 (
            .O(N__22012),
            .I(cmd_rdadctmp_14));
    InMux I__2003 (
            .O(N__22009),
            .I(N__22006));
    LocalMux I__2002 (
            .O(N__22006),
            .I(n19_adj_1700));
    InMux I__2001 (
            .O(N__22003),
            .I(N__22000));
    LocalMux I__2000 (
            .O(N__22000),
            .I(N__21997));
    Span4Mux_h I__1999 (
            .O(N__21997),
            .I(N__21994));
    Odrv4 I__1998 (
            .O(N__21994),
            .I(buf_data_iac_4));
    CascadeMux I__1997 (
            .O(N__21991),
            .I(n22_adj_1701_cascade_));
    InMux I__1996 (
            .O(N__21988),
            .I(N__21985));
    LocalMux I__1995 (
            .O(N__21985),
            .I(N__21980));
    InMux I__1994 (
            .O(N__21984),
            .I(N__21977));
    InMux I__1993 (
            .O(N__21983),
            .I(N__21974));
    Span4Mux_v I__1992 (
            .O(N__21980),
            .I(N__21971));
    LocalMux I__1991 (
            .O(N__21977),
            .I(N__21968));
    LocalMux I__1990 (
            .O(N__21974),
            .I(buf_adcdata_vac_7));
    Odrv4 I__1989 (
            .O(N__21971),
            .I(buf_adcdata_vac_7));
    Odrv4 I__1988 (
            .O(N__21968),
            .I(buf_adcdata_vac_7));
    InMux I__1987 (
            .O(N__21961),
            .I(N__21958));
    LocalMux I__1986 (
            .O(N__21958),
            .I(N__21953));
    InMux I__1985 (
            .O(N__21957),
            .I(N__21948));
    InMux I__1984 (
            .O(N__21956),
            .I(N__21948));
    Odrv4 I__1983 (
            .O(N__21953),
            .I(buf_adcdata_iac_4));
    LocalMux I__1982 (
            .O(N__21948),
            .I(buf_adcdata_iac_4));
    InMux I__1981 (
            .O(N__21943),
            .I(N__21938));
    InMux I__1980 (
            .O(N__21942),
            .I(N__21935));
    CascadeMux I__1979 (
            .O(N__21941),
            .I(N__21932));
    LocalMux I__1978 (
            .O(N__21938),
            .I(N__21929));
    LocalMux I__1977 (
            .O(N__21935),
            .I(N__21926));
    InMux I__1976 (
            .O(N__21932),
            .I(N__21923));
    Odrv4 I__1975 (
            .O(N__21929),
            .I(read_buf_14));
    Odrv4 I__1974 (
            .O(N__21926),
            .I(read_buf_14));
    LocalMux I__1973 (
            .O(N__21923),
            .I(read_buf_14));
    CascadeMux I__1972 (
            .O(N__21916),
            .I(N__21911));
    CascadeMux I__1971 (
            .O(N__21915),
            .I(N__21908));
    InMux I__1970 (
            .O(N__21914),
            .I(N__21905));
    InMux I__1969 (
            .O(N__21911),
            .I(N__21902));
    InMux I__1968 (
            .O(N__21908),
            .I(N__21899));
    LocalMux I__1967 (
            .O(N__21905),
            .I(N__21896));
    LocalMux I__1966 (
            .O(N__21902),
            .I(N__21893));
    LocalMux I__1965 (
            .O(N__21899),
            .I(read_buf_3));
    Odrv4 I__1964 (
            .O(N__21896),
            .I(read_buf_3));
    Odrv4 I__1963 (
            .O(N__21893),
            .I(read_buf_3));
    CascadeMux I__1962 (
            .O(N__21886),
            .I(N__21881));
    InMux I__1961 (
            .O(N__21885),
            .I(N__21878));
    InMux I__1960 (
            .O(N__21884),
            .I(N__21873));
    InMux I__1959 (
            .O(N__21881),
            .I(N__21873));
    LocalMux I__1958 (
            .O(N__21878),
            .I(read_buf_13));
    LocalMux I__1957 (
            .O(N__21873),
            .I(read_buf_13));
    CascadeMux I__1956 (
            .O(N__21868),
            .I(n19_adj_1690_cascade_));
    InMux I__1955 (
            .O(N__21865),
            .I(N__21862));
    LocalMux I__1954 (
            .O(N__21862),
            .I(N__21858));
    InMux I__1953 (
            .O(N__21861),
            .I(N__21854));
    Span4Mux_h I__1952 (
            .O(N__21858),
            .I(N__21851));
    InMux I__1951 (
            .O(N__21857),
            .I(N__21848));
    LocalMux I__1950 (
            .O(N__21854),
            .I(buf_adcdata_vac_6));
    Odrv4 I__1949 (
            .O(N__21851),
            .I(buf_adcdata_vac_6));
    LocalMux I__1948 (
            .O(N__21848),
            .I(buf_adcdata_vac_6));
    CascadeMux I__1947 (
            .O(N__21841),
            .I(n19_adj_1693_cascade_));
    InMux I__1946 (
            .O(N__21838),
            .I(N__21833));
    InMux I__1945 (
            .O(N__21837),
            .I(N__21828));
    InMux I__1944 (
            .O(N__21836),
            .I(N__21828));
    LocalMux I__1943 (
            .O(N__21833),
            .I(read_buf_10));
    LocalMux I__1942 (
            .O(N__21828),
            .I(read_buf_10));
    CascadeMux I__1941 (
            .O(N__21823),
            .I(N__21819));
    InMux I__1940 (
            .O(N__21822),
            .I(N__21815));
    InMux I__1939 (
            .O(N__21819),
            .I(N__21810));
    InMux I__1938 (
            .O(N__21818),
            .I(N__21810));
    LocalMux I__1937 (
            .O(N__21815),
            .I(N__21807));
    LocalMux I__1936 (
            .O(N__21810),
            .I(bit_cnt_2));
    Odrv4 I__1935 (
            .O(N__21807),
            .I(bit_cnt_2));
    CascadeMux I__1934 (
            .O(N__21802),
            .I(N__21799));
    InMux I__1933 (
            .O(N__21799),
            .I(N__21793));
    InMux I__1932 (
            .O(N__21798),
            .I(N__21786));
    InMux I__1931 (
            .O(N__21797),
            .I(N__21786));
    InMux I__1930 (
            .O(N__21796),
            .I(N__21786));
    LocalMux I__1929 (
            .O(N__21793),
            .I(N__21783));
    LocalMux I__1928 (
            .O(N__21786),
            .I(bit_cnt_1));
    Odrv4 I__1927 (
            .O(N__21783),
            .I(bit_cnt_1));
    InMux I__1926 (
            .O(N__21778),
            .I(N__21769));
    InMux I__1925 (
            .O(N__21777),
            .I(N__21769));
    InMux I__1924 (
            .O(N__21776),
            .I(N__21764));
    InMux I__1923 (
            .O(N__21775),
            .I(N__21758));
    InMux I__1922 (
            .O(N__21774),
            .I(N__21758));
    LocalMux I__1921 (
            .O(N__21769),
            .I(N__21755));
    InMux I__1920 (
            .O(N__21768),
            .I(N__21751));
    InMux I__1919 (
            .O(N__21767),
            .I(N__21748));
    LocalMux I__1918 (
            .O(N__21764),
            .I(N__21744));
    InMux I__1917 (
            .O(N__21763),
            .I(N__21741));
    LocalMux I__1916 (
            .O(N__21758),
            .I(N__21736));
    Span4Mux_h I__1915 (
            .O(N__21755),
            .I(N__21736));
    InMux I__1914 (
            .O(N__21754),
            .I(N__21733));
    LocalMux I__1913 (
            .O(N__21751),
            .I(N__21728));
    LocalMux I__1912 (
            .O(N__21748),
            .I(N__21728));
    InMux I__1911 (
            .O(N__21747),
            .I(N__21725));
    Odrv4 I__1910 (
            .O(N__21744),
            .I(dds_state_0_adj_1510));
    LocalMux I__1909 (
            .O(N__21741),
            .I(dds_state_0_adj_1510));
    Odrv4 I__1908 (
            .O(N__21736),
            .I(dds_state_0_adj_1510));
    LocalMux I__1907 (
            .O(N__21733),
            .I(dds_state_0_adj_1510));
    Odrv4 I__1906 (
            .O(N__21728),
            .I(dds_state_0_adj_1510));
    LocalMux I__1905 (
            .O(N__21725),
            .I(dds_state_0_adj_1510));
    InMux I__1904 (
            .O(N__21712),
            .I(N__21709));
    LocalMux I__1903 (
            .O(N__21709),
            .I(n8_adj_1686));
    InMux I__1902 (
            .O(N__21706),
            .I(N__21701));
    InMux I__1901 (
            .O(N__21705),
            .I(N__21698));
    InMux I__1900 (
            .O(N__21704),
            .I(N__21695));
    LocalMux I__1899 (
            .O(N__21701),
            .I(N__21692));
    LocalMux I__1898 (
            .O(N__21698),
            .I(N__21687));
    LocalMux I__1897 (
            .O(N__21695),
            .I(N__21687));
    Odrv4 I__1896 (
            .O(N__21692),
            .I(read_buf_11));
    Odrv4 I__1895 (
            .O(N__21687),
            .I(read_buf_11));
    InMux I__1894 (
            .O(N__21682),
            .I(N__21678));
    CascadeMux I__1893 (
            .O(N__21681),
            .I(N__21674));
    LocalMux I__1892 (
            .O(N__21678),
            .I(N__21671));
    InMux I__1891 (
            .O(N__21677),
            .I(N__21666));
    InMux I__1890 (
            .O(N__21674),
            .I(N__21666));
    Odrv4 I__1889 (
            .O(N__21671),
            .I(read_buf_12));
    LocalMux I__1888 (
            .O(N__21666),
            .I(read_buf_12));
    CascadeMux I__1887 (
            .O(N__21661),
            .I(\RTD.n22632_cascade_ ));
    IoInMux I__1886 (
            .O(N__21658),
            .I(N__21655));
    LocalMux I__1885 (
            .O(N__21655),
            .I(N__21652));
    Span12Mux_s0_v I__1884 (
            .O(N__21652),
            .I(N__21649));
    Odrv12 I__1883 (
            .O(N__21649),
            .I(DDS_CS1));
    CEMux I__1882 (
            .O(N__21646),
            .I(N__21643));
    LocalMux I__1881 (
            .O(N__21643),
            .I(N__21640));
    Span4Mux_h I__1880 (
            .O(N__21640),
            .I(N__21637));
    Odrv4 I__1879 (
            .O(N__21637),
            .I(\CLK_DDS.n9_adj_1489 ));
    CascadeMux I__1878 (
            .O(N__21634),
            .I(N__21630));
    InMux I__1877 (
            .O(N__21633),
            .I(N__21625));
    InMux I__1876 (
            .O(N__21630),
            .I(N__21625));
    LocalMux I__1875 (
            .O(N__21625),
            .I(read_buf_15));
    InMux I__1874 (
            .O(N__21622),
            .I(\ADC_VAC.n20685 ));
    InMux I__1873 (
            .O(N__21619),
            .I(\ADC_VAC.n20686 ));
    InMux I__1872 (
            .O(N__21616),
            .I(\ADC_VAC.n20687 ));
    InMux I__1871 (
            .O(N__21613),
            .I(\ADC_VAC.n20688 ));
    InMux I__1870 (
            .O(N__21610),
            .I(\ADC_VAC.n20689 ));
    CEMux I__1869 (
            .O(N__21607),
            .I(N__21604));
    LocalMux I__1868 (
            .O(N__21604),
            .I(\ADC_VAC.n13784 ));
    CascadeMux I__1867 (
            .O(N__21601),
            .I(\ADC_VAC.n13784_cascade_ ));
    SRMux I__1866 (
            .O(N__21598),
            .I(N__21595));
    LocalMux I__1865 (
            .O(N__21595),
            .I(N__21592));
    Span4Mux_h I__1864 (
            .O(N__21592),
            .I(N__21589));
    Odrv4 I__1863 (
            .O(N__21589),
            .I(\ADC_VAC.n15660 ));
    CEMux I__1862 (
            .O(N__21586),
            .I(N__21582));
    CEMux I__1861 (
            .O(N__21585),
            .I(N__21579));
    LocalMux I__1860 (
            .O(N__21582),
            .I(N__21576));
    LocalMux I__1859 (
            .O(N__21579),
            .I(N__21573));
    Span4Mux_v I__1858 (
            .O(N__21576),
            .I(N__21570));
    Span4Mux_h I__1857 (
            .O(N__21573),
            .I(N__21567));
    Odrv4 I__1856 (
            .O(N__21570),
            .I(\CLK_DDS.n9 ));
    Odrv4 I__1855 (
            .O(N__21567),
            .I(\CLK_DDS.n9 ));
    InMux I__1854 (
            .O(N__21562),
            .I(N__21559));
    LocalMux I__1853 (
            .O(N__21559),
            .I(N__21556));
    Span4Mux_h I__1852 (
            .O(N__21556),
            .I(N__21551));
    InMux I__1851 (
            .O(N__21555),
            .I(N__21546));
    InMux I__1850 (
            .O(N__21554),
            .I(N__21546));
    Odrv4 I__1849 (
            .O(N__21551),
            .I(buf_adcdata_vac_4));
    LocalMux I__1848 (
            .O(N__21546),
            .I(buf_adcdata_vac_4));
    CascadeMux I__1847 (
            .O(N__21541),
            .I(N__21538));
    InMux I__1846 (
            .O(N__21538),
            .I(N__21534));
    InMux I__1845 (
            .O(N__21537),
            .I(N__21531));
    LocalMux I__1844 (
            .O(N__21534),
            .I(cmd_rdadctmp_1_adj_1547));
    LocalMux I__1843 (
            .O(N__21531),
            .I(cmd_rdadctmp_1_adj_1547));
    CascadeMux I__1842 (
            .O(N__21526),
            .I(N__21523));
    InMux I__1841 (
            .O(N__21523),
            .I(N__21520));
    LocalMux I__1840 (
            .O(N__21520),
            .I(N__21516));
    CascadeMux I__1839 (
            .O(N__21519),
            .I(N__21513));
    Span4Mux_h I__1838 (
            .O(N__21516),
            .I(N__21509));
    InMux I__1837 (
            .O(N__21513),
            .I(N__21504));
    InMux I__1836 (
            .O(N__21512),
            .I(N__21504));
    Odrv4 I__1835 (
            .O(N__21509),
            .I(cmd_rdadctmp_14_adj_1534));
    LocalMux I__1834 (
            .O(N__21504),
            .I(cmd_rdadctmp_14_adj_1534));
    InMux I__1833 (
            .O(N__21499),
            .I(bfn_2_14_0_));
    InMux I__1832 (
            .O(N__21496),
            .I(\ADC_VAC.n20683 ));
    InMux I__1831 (
            .O(N__21493),
            .I(\ADC_VAC.n20684 ));
    CEMux I__1830 (
            .O(N__21490),
            .I(N__21487));
    LocalMux I__1829 (
            .O(N__21487),
            .I(\RTD.n12262 ));
    CascadeMux I__1828 (
            .O(N__21484),
            .I(N__21481));
    InMux I__1827 (
            .O(N__21481),
            .I(N__21478));
    LocalMux I__1826 (
            .O(N__21478),
            .I(N__21475));
    Span4Mux_v I__1825 (
            .O(N__21475),
            .I(N__21472));
    Span4Mux_h I__1824 (
            .O(N__21472),
            .I(N__21469));
    Span4Mux_v I__1823 (
            .O(N__21469),
            .I(N__21466));
    Span4Mux_v I__1822 (
            .O(N__21466),
            .I(N__21463));
    Odrv4 I__1821 (
            .O(N__21463),
            .I(RTD_SDO));
    SRMux I__1820 (
            .O(N__21460),
            .I(N__21457));
    LocalMux I__1819 (
            .O(N__21457),
            .I(\CLK_DDS.n18366 ));
    InMux I__1818 (
            .O(N__21454),
            .I(N__21447));
    InMux I__1817 (
            .O(N__21453),
            .I(N__21440));
    InMux I__1816 (
            .O(N__21452),
            .I(N__21440));
    InMux I__1815 (
            .O(N__21451),
            .I(N__21440));
    InMux I__1814 (
            .O(N__21450),
            .I(N__21437));
    LocalMux I__1813 (
            .O(N__21447),
            .I(bit_cnt_0_adj_1512));
    LocalMux I__1812 (
            .O(N__21440),
            .I(bit_cnt_0_adj_1512));
    LocalMux I__1811 (
            .O(N__21437),
            .I(bit_cnt_0_adj_1512));
    InMux I__1810 (
            .O(N__21430),
            .I(N__21426));
    InMux I__1809 (
            .O(N__21429),
            .I(N__21423));
    LocalMux I__1808 (
            .O(N__21426),
            .I(bit_cnt_3));
    LocalMux I__1807 (
            .O(N__21423),
            .I(bit_cnt_3));
    InMux I__1806 (
            .O(N__21418),
            .I(N__21415));
    LocalMux I__1805 (
            .O(N__21415),
            .I(n22326));
    CascadeMux I__1804 (
            .O(N__21412),
            .I(N__21409));
    InMux I__1803 (
            .O(N__21409),
            .I(N__21406));
    LocalMux I__1802 (
            .O(N__21406),
            .I(N__21403));
    Span4Mux_v I__1801 (
            .O(N__21403),
            .I(N__21400));
    Span4Mux_h I__1800 (
            .O(N__21400),
            .I(N__21397));
    Odrv4 I__1799 (
            .O(N__21397),
            .I(VAC_MISO));
    CascadeMux I__1798 (
            .O(N__21394),
            .I(N__21391));
    InMux I__1797 (
            .O(N__21391),
            .I(N__21385));
    InMux I__1796 (
            .O(N__21390),
            .I(N__21385));
    LocalMux I__1795 (
            .O(N__21385),
            .I(cmd_rdadctmp_0_adj_1548));
    IoInMux I__1794 (
            .O(N__21382),
            .I(N__21379));
    LocalMux I__1793 (
            .O(N__21379),
            .I(N__21375));
    CascadeMux I__1792 (
            .O(N__21378),
            .I(N__21372));
    Span12Mux_s4_h I__1791 (
            .O(N__21375),
            .I(N__21369));
    InMux I__1790 (
            .O(N__21372),
            .I(N__21366));
    Odrv12 I__1789 (
            .O(N__21369),
            .I(VAC_SCLK));
    LocalMux I__1788 (
            .O(N__21366),
            .I(VAC_SCLK));
    CascadeMux I__1787 (
            .O(N__21361),
            .I(n14_cascade_));
    InMux I__1786 (
            .O(N__21358),
            .I(N__21355));
    LocalMux I__1785 (
            .O(N__21355),
            .I(n21889));
    IoInMux I__1784 (
            .O(N__21352),
            .I(N__21349));
    LocalMux I__1783 (
            .O(N__21349),
            .I(N__21345));
    CascadeMux I__1782 (
            .O(N__21348),
            .I(N__21342));
    Span12Mux_s4_h I__1781 (
            .O(N__21345),
            .I(N__21339));
    InMux I__1780 (
            .O(N__21342),
            .I(N__21336));
    Odrv12 I__1779 (
            .O(N__21339),
            .I(VAC_CS));
    LocalMux I__1778 (
            .O(N__21336),
            .I(VAC_CS));
    IoInMux I__1777 (
            .O(N__21331),
            .I(N__21328));
    LocalMux I__1776 (
            .O(N__21328),
            .I(N__21325));
    Span4Mux_s3_v I__1775 (
            .O(N__21325),
            .I(N__21322));
    Span4Mux_v I__1774 (
            .O(N__21322),
            .I(N__21318));
    CascadeMux I__1773 (
            .O(N__21321),
            .I(N__21315));
    Span4Mux_v I__1772 (
            .O(N__21318),
            .I(N__21312));
    InMux I__1771 (
            .O(N__21315),
            .I(N__21309));
    Odrv4 I__1770 (
            .O(N__21312),
            .I(DDS_SCK1));
    LocalMux I__1769 (
            .O(N__21309),
            .I(DDS_SCK1));
    IoInMux I__1768 (
            .O(N__21304),
            .I(N__21301));
    LocalMux I__1767 (
            .O(N__21301),
            .I(N__21298));
    Span4Mux_s2_h I__1766 (
            .O(N__21298),
            .I(N__21295));
    Span4Mux_v I__1765 (
            .O(N__21295),
            .I(N__21292));
    Odrv4 I__1764 (
            .O(N__21292),
            .I(RTD_SCLK));
    CEMux I__1763 (
            .O(N__21289),
            .I(N__21286));
    LocalMux I__1762 (
            .O(N__21286),
            .I(N__21283));
    Odrv12 I__1761 (
            .O(N__21283),
            .I(\RTD.n8 ));
    IoInMux I__1760 (
            .O(N__21280),
            .I(N__21277));
    LocalMux I__1759 (
            .O(N__21277),
            .I(N__21274));
    IoSpan4Mux I__1758 (
            .O(N__21274),
            .I(N__21271));
    IoSpan4Mux I__1757 (
            .O(N__21271),
            .I(N__21268));
    Span4Mux_s3_h I__1756 (
            .O(N__21268),
            .I(N__21265));
    Odrv4 I__1755 (
            .O(N__21265),
            .I(RTD_SDI));
    SRMux I__1754 (
            .O(N__21262),
            .I(N__21259));
    LocalMux I__1753 (
            .O(N__21259),
            .I(\RTD.n21253 ));
    IoInMux I__1752 (
            .O(N__21256),
            .I(N__21253));
    LocalMux I__1751 (
            .O(N__21253),
            .I(N__21250));
    IoSpan4Mux I__1750 (
            .O(N__21250),
            .I(N__21247));
    IoSpan4Mux I__1749 (
            .O(N__21247),
            .I(N__21244));
    Odrv4 I__1748 (
            .O(N__21244),
            .I(ICE_SYSCLK));
    IoInMux I__1747 (
            .O(N__21241),
            .I(N__21238));
    LocalMux I__1746 (
            .O(N__21238),
            .I(N__21235));
    IoSpan4Mux I__1745 (
            .O(N__21235),
            .I(N__21232));
    Span4Mux_s3_v I__1744 (
            .O(N__21232),
            .I(N__21229));
    Sp12to4 I__1743 (
            .O(N__21229),
            .I(N__21226));
    Span12Mux_h I__1742 (
            .O(N__21226),
            .I(N__21223));
    Odrv12 I__1741 (
            .O(N__21223),
            .I(ICE_GPMO_2));
    INV \INVADC_VDC.genclk.t0off_i8C  (
            .O(\INVADC_VDC.genclk.t0off_i8C_net ),
            .I(N__48417));
    INV \INVADC_VDC.genclk.t0off_i0C  (
            .O(\INVADC_VDC.genclk.t0off_i0C_net ),
            .I(N__48416));
    INV \INVADC_VDC.genclk.div_state_i0C  (
            .O(\INVADC_VDC.genclk.div_state_i0C_net ),
            .I(N__48415));
    INV \INVADC_VDC.genclk.div_state_i1C  (
            .O(\INVADC_VDC.genclk.div_state_i1C_net ),
            .I(N__48412));
    INV \INVcomm_spi.data_valid_85C  (
            .O(\INVcomm_spi.data_valid_85C_net ),
            .I(N__61891));
    INV INVdds0_mclk_297C (
            .O(INVdds0_mclk_297C_net),
            .I(N__48414));
    INV INVdds0_mclkcnt_i7_3792__i0C (
            .O(INVdds0_mclkcnt_i7_3792__i0C_net),
            .I(N__48413));
    INV \INVADC_VDC.genclk.t0on_i8C  (
            .O(\INVADC_VDC.genclk.t0on_i8C_net ),
            .I(N__48411));
    INV \INVADC_VDC.genclk.t0on_i0C  (
            .O(\INVADC_VDC.genclk.t0on_i0C_net ),
            .I(N__48409));
    INV INVdata_cntvec_i0_i8C (
            .O(INVdata_cntvec_i0_i8C_net),
            .I(N__61973));
    INV INVdata_cntvec_i0_i0C (
            .O(INVdata_cntvec_i0_i0C_net),
            .I(N__61956));
    INV \INVcomm_spi.bit_cnt_3787__i3C  (
            .O(\INVcomm_spi.bit_cnt_3787__i3C_net ),
            .I(N__53678));
    INV \INVADC_VDC.genclk.t_clk_24C  (
            .O(\INVADC_VDC.genclk.t_clk_24C_net ),
            .I(N__48402));
    INV \INVcomm_spi.MISO_48_12606_12607_setC  (
            .O(\INVcomm_spi.MISO_48_12606_12607_setC_net ),
            .I(N__61937));
    INV \INVcomm_spi.imiso_83_12612_12613_setC  (
            .O(\INVcomm_spi.imiso_83_12612_12613_setC_net ),
            .I(N__53706));
    INV \INVcomm_spi.MISO_48_12606_12607_resetC  (
            .O(\INVcomm_spi.MISO_48_12606_12607_resetC_net ),
            .I(N__61829));
    INV INVacadc_skipcnt_i0_i9C (
            .O(INVacadc_skipcnt_i0_i9C_net),
            .I(N__61969));
    INV INVacadc_skipcnt_i0_i1C (
            .O(INVacadc_skipcnt_i0_i1C_net),
            .I(N__61951));
    INV INVacadc_skipcnt_i0_i0C (
            .O(INVacadc_skipcnt_i0_i0C_net),
            .I(N__61935));
    INV INVeis_state_i0C (
            .O(INVeis_state_i0C_net),
            .I(N__61887));
    INV INVeis_state_i2C (
            .O(INVeis_state_i2C_net),
            .I(N__61900));
    INV INVeis_end_302C (
            .O(INVeis_end_302C_net),
            .I(N__61886));
    INV \INVcomm_spi.imiso_83_12612_12613_resetC  (
            .O(\INVcomm_spi.imiso_83_12612_12613_resetC_net ),
            .I(N__53638));
    INV INVdata_count_i0_i8C (
            .O(INVdata_count_i0_i8C_net),
            .I(N__61913));
    INV INVdata_count_i0_i0C (
            .O(INVdata_count_i0_i0C_net),
            .I(N__61899));
    INV INVacadc_trig_303C (
            .O(INVacadc_trig_303C_net),
            .I(N__61947));
    INV INViac_raw_buf_vac_raw_buf_merged2WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .I(N__61923));
    INV INViac_raw_buf_vac_raw_buf_merged7WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .I(N__62014));
    INV INViac_raw_buf_vac_raw_buf_merged1WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .I(N__61851));
    INV INViac_raw_buf_vac_raw_buf_merged6WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .I(N__62011));
    INV INViac_raw_buf_vac_raw_buf_merged0WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .I(N__61838));
    INV INViac_raw_buf_vac_raw_buf_merged5WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .I(N__62004));
    INV INViac_raw_buf_vac_raw_buf_merged9WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .I(N__61882));
    INV INViac_raw_buf_vac_raw_buf_merged4WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .I(N__61989));
    INV INViac_raw_buf_vac_raw_buf_merged8WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .I(N__61860));
    INV INViac_raw_buf_vac_raw_buf_merged10WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .I(N__61868));
    INV INViac_raw_buf_vac_raw_buf_merged3WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .I(N__61960));
    INV INViac_raw_buf_vac_raw_buf_merged11WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .I(N__61893));
    defparam IN_MUX_bfv_17_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_5_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(n20773),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(n20781),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(n20789),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(n20797),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(n20805),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(n20637_THRU_CRY_6_THRU_CO),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(n20645),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(n20629),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(n20620),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(n20668),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(n20659),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_23_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_5_0_));
    defparam IN_MUX_bfv_23_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_6_0_ (
            .carryinitin(\ADC_VDC.genclk.n20743 ),
            .carryinitout(bfn_23_6_0_));
    defparam IN_MUX_bfv_19_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_5_0_));
    defparam IN_MUX_bfv_19_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_6_0_ (
            .carryinitin(\ADC_VDC.genclk.n20758 ),
            .carryinitout(bfn_19_6_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\ADC_VDC.n20732 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\ADC_VDC.n20697 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\ADC_VDC.n20705 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\ADC_VDC.n20713 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\ADC_VDC.n20721 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_16_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \RTD.SCLK_51_LC_1_3_5 .C_ON=1'b0;
    defparam \RTD.SCLK_51_LC_1_3_5 .SEQ_MODE=4'b1000;
    defparam \RTD.SCLK_51_LC_1_3_5 .LUT_INIT=16'b0011100000011110;
    LogicCell40 \RTD.SCLK_51_LC_1_3_5  (
            .in0(N__26680),
            .in1(N__26864),
            .in2(N__26521),
            .in3(N__26249),
            .lcout(RTD_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35006),
            .ce(N__21289),
            .sr(_gnd_net_));
    defparam \RTD.i20152_4_lut_4_lut_LC_1_4_0 .C_ON=1'b0;
    defparam \RTD.i20152_4_lut_4_lut_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i20152_4_lut_4_lut_LC_1_4_0 .LUT_INIT=16'b1111011111011111;
    LogicCell40 \RTD.i20152_4_lut_4_lut_LC_1_4_0  (
            .in0(N__26837),
            .in1(N__26674),
            .in2(N__26503),
            .in3(N__26223),
            .lcout(\RTD.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_4_lut_LC_1_5_4 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_4_lut_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_4_lut_LC_1_5_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \RTD.i2_3_lut_4_lut_LC_1_5_4  (
            .in0(N__26866),
            .in1(N__26675),
            .in2(N__26519),
            .in3(N__26229),
            .lcout(\RTD.n21253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.MOSI_59_LC_1_6_3 .C_ON=1'b0;
    defparam \RTD.MOSI_59_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \RTD.MOSI_59_LC_1_6_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \RTD.MOSI_59_LC_1_6_3  (
            .in0(N__22657),
            .in1(N__26510),
            .in2(N__22768),
            .in3(N__26234),
            .lcout(RTD_SDI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35038),
            .ce(N__21490),
            .sr(N__21262));
    defparam \CLK_DDS.bit_cnt_i3_LC_1_7_0 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i3_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i3_LC_1_7_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \CLK_DDS.bit_cnt_i3_LC_1_7_0  (
            .in0(N__21453),
            .in1(N__21798),
            .in2(N__21823),
            .in3(N__21430),
            .lcout(bit_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61925),
            .ce(N__24640),
            .sr(N__21460));
    defparam \CLK_DDS.bit_cnt_i2_LC_1_7_1 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i2_LC_1_7_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i2_LC_1_7_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \CLK_DDS.bit_cnt_i2_LC_1_7_1  (
            .in0(N__21797),
            .in1(N__21452),
            .in2(_gnd_net_),
            .in3(N__21818),
            .lcout(bit_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61925),
            .ce(N__24640),
            .sr(N__21460));
    defparam \CLK_DDS.bit_cnt_i1_LC_1_7_2 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i1_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i1_LC_1_7_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \CLK_DDS.bit_cnt_i1_LC_1_7_2  (
            .in0(N__21451),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21796),
            .lcout(bit_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61925),
            .ce(N__24640),
            .sr(N__21460));
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_1_13_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_1_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_1_13_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i1_LC_1_13_1  (
            .in0(N__21537),
            .in1(N__33954),
            .in2(N__21394),
            .in3(N__35925),
            .lcout(cmd_rdadctmp_1_adj_1547),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62005),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_1_13_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_1_13_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i0_LC_1_13_3  (
            .in0(N__21390),
            .in1(N__33953),
            .in2(N__21412),
            .in3(N__35924),
            .lcout(cmd_rdadctmp_0_adj_1548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62005),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i1_LC_1_14_7 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i1_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i1_LC_1_14_7 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \ADC_VAC.adc_state_i1_LC_1_14_7  (
            .in0(N__32099),
            .in1(N__31992),
            .in2(_gnd_net_),
            .in3(N__35926),
            .lcout(adc_state_1_adj_1515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62009),
            .ce(N__22267),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_303_LC_1_15_0.C_ON=1'b0;
    defparam i1_2_lut_adj_303_LC_1_15_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_303_LC_1_15_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_303_LC_1_15_0 (
            .in0(_gnd_net_),
            .in1(N__31970),
            .in2(_gnd_net_),
            .in3(N__32093),
            .lcout(n21889),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.SCLK_35_LC_1_15_1 .C_ON=1'b0;
    defparam \ADC_VAC.SCLK_35_LC_1_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.SCLK_35_LC_1_15_1 .LUT_INIT=16'b1011000011100010;
    LogicCell40 \ADC_VAC.SCLK_35_LC_1_15_1  (
            .in0(N__32095),
            .in1(N__31972),
            .in2(N__21378),
            .in3(N__35913),
            .lcout(VAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62012),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_196_LC_1_15_3.C_ON=1'b0;
    defparam i1_4_lut_adj_196_LC_1_15_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_196_LC_1_15_3.LUT_INIT=16'b0000110100001110;
    LogicCell40 i1_4_lut_adj_196_LC_1_15_3 (
            .in0(N__32094),
            .in1(N__31971),
            .in2(N__21348),
            .in3(N__35911),
            .lcout(),
            .ltout(n14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.CS_37_LC_1_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.CS_37_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.CS_37_LC_1_15_4 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \ADC_VAC.CS_37_LC_1_15_4  (
            .in0(N__35912),
            .in1(N__22310),
            .in2(N__21361),
            .in3(N__21358),
            .lcout(VAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62012),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i0_LC_2_6_0 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i0_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i0_LC_2_6_0 .LUT_INIT=16'b0000111101000000;
    LogicCell40 \CLK_DDS.bit_cnt_i0_LC_2_6_0  (
            .in0(N__24704),
            .in1(N__21774),
            .in2(N__24639),
            .in3(N__21454),
            .lcout(bit_cnt_0_adj_1512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61894),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.SCLK_27_LC_2_6_1 .C_ON=1'b0;
    defparam \CLK_DDS.SCLK_27_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.SCLK_27_LC_2_6_1 .LUT_INIT=16'b0010000011111001;
    LogicCell40 \CLK_DDS.SCLK_27_LC_2_6_1  (
            .in0(N__21775),
            .in1(N__24614),
            .in2(N__21321),
            .in3(N__24703),
            .lcout(DDS_SCK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61894),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i27_4_lut_4_lut_LC_2_6_3 .C_ON=1'b0;
    defparam \RTD.i27_4_lut_4_lut_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i27_4_lut_4_lut_LC_2_6_3 .LUT_INIT=16'b1111000010010100;
    LogicCell40 \RTD.i27_4_lut_4_lut_LC_2_6_3  (
            .in0(N__26862),
            .in1(N__26676),
            .in2(N__26520),
            .in3(N__26233),
            .lcout(\RTD.n12262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i7_LC_2_6_5.C_ON=1'b0;
    defparam buf_cfgRTD_i7_LC_2_6_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i7_LC_2_6_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i7_LC_2_6_5 (
            .in0(N__57877),
            .in1(N__48800),
            .in2(N__46654),
            .in3(N__35337),
            .lcout(buf_cfgRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61894),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i0_LC_2_7_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i0_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i0_LC_2_7_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \RTD.read_buf_i0_LC_2_7_2  (
            .in0(N__22529),
            .in1(N__24083),
            .in2(N__21484),
            .in3(N__23976),
            .lcout(read_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35042),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i1_3_lut_LC_2_7_5 .C_ON=1'b0;
    defparam \CLK_DDS.i1_3_lut_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i1_3_lut_LC_2_7_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \CLK_DDS.i1_3_lut_LC_2_7_5  (
            .in0(N__24546),
            .in1(N__24691),
            .in2(_gnd_net_),
            .in3(N__21767),
            .lcout(\CLK_DDS.n18366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19900_2_lut_LC_2_7_6.C_ON=1'b0;
    defparam i19900_2_lut_LC_2_7_6.SEQ_MODE=4'b0000;
    defparam i19900_2_lut_LC_2_7_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i19900_2_lut_LC_2_7_6 (
            .in0(N__21450),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21429),
            .lcout(n22326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i1_LC_2_7_7 .C_ON=1'b0;
    defparam \RTD.read_buf_i1_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i1_LC_2_7_7 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \RTD.read_buf_i1_LC_2_7_7  (
            .in0(N__23975),
            .in1(N__22482),
            .in2(N__24091),
            .in3(N__22530),
            .lcout(read_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35042),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i0_LC_2_8_0 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i0_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i0_LC_2_8_0 .LUT_INIT=16'b1100010100000101;
    LogicCell40 \CLK_DDS.dds_state_i0_LC_2_8_0  (
            .in0(N__21763),
            .in1(N__21712),
            .in2(N__24609),
            .in3(N__21418),
            .lcout(dds_state_0_adj_1510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61926),
            .ce(N__21585),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i20153_4_lut_LC_2_9_5 .C_ON=1'b0;
    defparam \CLK_DDS.i20153_4_lut_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i20153_4_lut_LC_2_9_5 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \CLK_DDS.i20153_4_lut_LC_2_9_5  (
            .in0(N__24522),
            .in1(N__21754),
            .in2(N__56236),
            .in3(N__24706),
            .lcout(\CLK_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i6_LC_2_9_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i6_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i6_LC_2_9_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i6_LC_2_9_6  (
            .in0(N__35610),
            .in1(N__35946),
            .in2(N__21526),
            .in3(N__21861),
            .lcout(buf_adcdata_vac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61943),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i1_LC_2_10_0 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i1_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i1_LC_2_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLK_DDS.dds_state_i1_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__24707),
            .in2(_gnd_net_),
            .in3(N__21768),
            .lcout(dds_state_1_adj_1509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61961),
            .ce(N__21586),
            .sr(N__24635));
    defparam \ADC_VAC.ADC_DATA_i4_LC_2_11_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i4_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i4_LC_2_11_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i4_LC_2_11_2  (
            .in0(N__21555),
            .in1(N__35602),
            .in2(N__24321),
            .in3(N__35923),
            .lcout(buf_adcdata_vac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61977),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_4_i19_3_lut_LC_2_11_7.C_ON=1'b0;
    defparam mux_127_Mux_4_i19_3_lut_LC_2_11_7.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_4_i19_3_lut_LC_2_11_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_4_i19_3_lut_LC_2_11_7 (
            .in0(N__24985),
            .in1(N__21554),
            .in2(_gnd_net_),
            .in3(N__59112),
            .lcout(n19_adj_1700),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_2_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_2_12_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i2_LC_2_12_6  (
            .in0(N__35868),
            .in1(N__22698),
            .in2(N__21541),
            .in3(N__34001),
            .lcout(cmd_rdadctmp_2_adj_1546),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61990),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_2_13_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_2_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_2_13_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i14_LC_2_13_3  (
            .in0(N__21512),
            .in1(N__33979),
            .in2(N__22950),
            .in3(N__35777),
            .lcout(cmd_rdadctmp_14_adj_1534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61999),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_2_13_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_2_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_2_13_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i15_LC_2_13_5  (
            .in0(N__22205),
            .in1(N__33980),
            .in2(N__21519),
            .in3(N__35778),
            .lcout(cmd_rdadctmp_15_adj_1533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61999),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_2_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_2_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_2_13_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i13_LC_2_13_7  (
            .in0(N__22943),
            .in1(N__33978),
            .in2(N__24322),
            .in3(N__35776),
            .lcout(cmd_rdadctmp_13_adj_1535),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61999),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.bit_cnt_i0_LC_2_14_0 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i0_LC_2_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i0_LC_2_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i0_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__22375),
            .in2(_gnd_net_),
            .in3(N__21499),
            .lcout(\ADC_VAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\ADC_VAC.n20683 ),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.bit_cnt_i1_LC_2_14_1 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i1_LC_2_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i1_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i1_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__22120),
            .in2(_gnd_net_),
            .in3(N__21496),
            .lcout(\ADC_VAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC.n20683 ),
            .carryout(\ADC_VAC.n20684 ),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.bit_cnt_i2_LC_2_14_2 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i2_LC_2_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i2_LC_2_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i2_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__22132),
            .in2(_gnd_net_),
            .in3(N__21493),
            .lcout(\ADC_VAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC.n20684 ),
            .carryout(\ADC_VAC.n20685 ),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.bit_cnt_i3_LC_2_14_3 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i3_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i3_LC_2_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i3_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__22107),
            .in2(_gnd_net_),
            .in3(N__21622),
            .lcout(\ADC_VAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC.n20685 ),
            .carryout(\ADC_VAC.n20686 ),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.bit_cnt_i4_LC_2_14_4 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i4_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i4_LC_2_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i4_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__22093),
            .in2(_gnd_net_),
            .in3(N__21619),
            .lcout(\ADC_VAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC.n20686 ),
            .carryout(\ADC_VAC.n20687 ),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.bit_cnt_i5_LC_2_14_5 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i5_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i5_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i5_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__22345),
            .in2(_gnd_net_),
            .in3(N__21616),
            .lcout(\ADC_VAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC.n20687 ),
            .carryout(\ADC_VAC.n20688 ),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.bit_cnt_i6_LC_2_14_6 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i6_LC_2_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i6_LC_2_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i6_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__22387),
            .in2(_gnd_net_),
            .in3(N__21613),
            .lcout(\ADC_VAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC.n20688 ),
            .carryout(\ADC_VAC.n20689 ),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.bit_cnt_i7_LC_2_14_7 .C_ON=1'b0;
    defparam \ADC_VAC.bit_cnt_i7_LC_2_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i7_LC_2_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i7_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__22360),
            .in2(_gnd_net_),
            .in3(N__21610),
            .lcout(\ADC_VAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62006),
            .ce(N__21607),
            .sr(N__21598));
    defparam \ADC_VAC.i1_4_lut_adj_48_LC_2_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_adj_48_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_adj_48_LC_2_15_2 .LUT_INIT=16'b0000000001010010;
    LogicCell40 \ADC_VAC.i1_4_lut_adj_48_LC_2_15_2  (
            .in0(N__31963),
            .in1(N__22311),
            .in2(N__32092),
            .in3(N__35715),
            .lcout(\ADC_VAC.n13784 ),
            .ltout(\ADC_VAC.n13784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i12937_2_lut_LC_2_15_3 .C_ON=1'b0;
    defparam \ADC_VAC.i12937_2_lut_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i12937_2_lut_LC_2_15_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \ADC_VAC.i12937_2_lut_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21601),
            .in3(N__32071),
            .lcout(\ADC_VAC.n15660 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i20201_2_lut_LC_2_15_6 .C_ON=1'b0;
    defparam \ADC_VAC.i20201_2_lut_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i20201_2_lut_LC_2_15_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_VAC.i20201_2_lut_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__35716),
            .in2(_gnd_net_),
            .in3(N__22321),
            .lcout(\ADC_VAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i20130_4_lut_LC_3_4_0 .C_ON=1'b0;
    defparam \CLK_DDS.i20130_4_lut_LC_3_4_0 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i20130_4_lut_LC_3_4_0 .LUT_INIT=16'b1000100111001100;
    LogicCell40 \CLK_DDS.i20130_4_lut_LC_3_4_0  (
            .in0(N__24610),
            .in1(N__24684),
            .in2(N__56232),
            .in3(N__21777),
            .lcout(\CLK_DDS.n13376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i23_4_lut_LC_3_4_1 .C_ON=1'b0;
    defparam \CLK_DDS.i23_4_lut_LC_3_4_1 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i23_4_lut_LC_3_4_1 .LUT_INIT=16'b1111000010100111;
    LogicCell40 \CLK_DDS.i23_4_lut_LC_3_4_1  (
            .in0(N__21778),
            .in1(N__56228),
            .in2(N__24705),
            .in3(N__24611),
            .lcout(\CLK_DDS.n9_adj_1489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i2_LC_3_4_2 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i2_LC_3_4_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i2_LC_3_4_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \CLK_DDS.dds_state_i2_LC_3_4_2  (
            .in0(N__24612),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24688),
            .lcout(dds_state_2_adj_1508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61858),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i20043_3_lut_LC_3_4_5 .C_ON=1'b0;
    defparam \RTD.i20043_3_lut_LC_3_4_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i20043_3_lut_LC_3_4_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \RTD.i20043_3_lut_LC_3_4_5  (
            .in0(N__35131),
            .in1(N__26654),
            .in2(_gnd_net_),
            .in3(N__32875),
            .lcout(),
            .ltout(\RTD.n22632_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i17362_4_lut_LC_3_4_6 .C_ON=1'b0;
    defparam \RTD.i17362_4_lut_LC_3_4_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i17362_4_lut_LC_3_4_6 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \RTD.i17362_4_lut_LC_3_4_6  (
            .in0(N__23203),
            .in1(N__26838),
            .in2(N__21661),
            .in3(N__22429),
            .lcout(\RTD.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.CS_28_LC_3_5_2 .C_ON=1'b0;
    defparam \CLK_DDS.CS_28_LC_3_5_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.CS_28_LC_3_5_2 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \CLK_DDS.CS_28_LC_3_5_2  (
            .in0(N__24613),
            .in1(N__24689),
            .in2(_gnd_net_),
            .in3(N__21776),
            .lcout(DDS_CS1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61869),
            .ce(N__21646),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i15_LC_3_6_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i15_LC_3_6_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i15_LC_3_6_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \RTD.read_buf_i15_LC_3_6_0  (
            .in0(N__21943),
            .in1(N__24053),
            .in2(N__21634),
            .in3(N__23979),
            .lcout(read_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35013),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i15_LC_3_6_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i15_LC_3_6_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i15_LC_3_6_1 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \RTD.READ_DATA_i15_LC_3_6_1  (
            .in0(N__35298),
            .in1(N__21633),
            .in2(N__26518),
            .in3(N__23811),
            .lcout(buf_readRTD_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35013),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i10_LC_3_6_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i10_LC_3_6_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i10_LC_3_6_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i10_LC_3_6_3  (
            .in0(N__21838),
            .in1(N__23810),
            .in2(N__28740),
            .in3(N__26486),
            .lcout(buf_readRTD_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35013),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19153_2_lut_LC_3_6_4 .C_ON=1'b0;
    defparam \RTD.i19153_2_lut_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i19153_2_lut_LC_3_6_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i19153_2_lut_LC_3_6_4  (
            .in0(_gnd_net_),
            .in1(N__26222),
            .in2(_gnd_net_),
            .in3(N__26858),
            .lcout(\RTD.n22079 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i4_LC_3_6_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i4_LC_3_6_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i4_LC_3_6_6 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.read_buf_i4_LC_3_6_6  (
            .in0(N__22508),
            .in1(N__23980),
            .in2(N__21916),
            .in3(N__24054),
            .lcout(\RTD.read_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35013),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i10_LC_3_7_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i10_LC_3_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i10_LC_3_7_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \RTD.read_buf_i10_LC_3_7_1  (
            .in0(N__21836),
            .in1(N__24078),
            .in2(N__23722),
            .in3(N__23982),
            .lcout(read_buf_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35030),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i11_LC_3_7_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i11_LC_3_7_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i11_LC_3_7_2 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \RTD.read_buf_i11_LC_3_7_2  (
            .in0(N__23981),
            .in1(N__21837),
            .in2(N__24090),
            .in3(N__21704),
            .lcout(read_buf_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35030),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i3_LC_3_7_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i3_LC_3_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i3_LC_3_7_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \RTD.read_buf_i3_LC_3_7_3  (
            .in0(N__22471),
            .in1(N__24079),
            .in2(N__21915),
            .in3(N__23983),
            .lcout(read_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35030),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i14_LC_3_7_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i14_LC_3_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i14_LC_3_7_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i14_LC_3_7_4  (
            .in0(N__21942),
            .in1(N__23816),
            .in2(N__23403),
            .in3(N__26492),
            .lcout(buf_readRTD_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35030),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i12_LC_3_7_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i12_LC_3_7_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i12_LC_3_7_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i12_LC_3_7_5  (
            .in0(N__26490),
            .in1(N__21682),
            .in2(N__28851),
            .in3(N__23818),
            .lcout(buf_readRTD_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35030),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i11_LC_3_7_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i11_LC_3_7_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i11_LC_3_7_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i11_LC_3_7_6  (
            .in0(N__21705),
            .in1(N__23815),
            .in2(N__25242),
            .in3(N__26491),
            .lcout(buf_readRTD_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35030),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_7_7 .C_ON=1'b0;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_7_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \CLK_DDS.i3_3_lut_4_lut_LC_3_7_7  (
            .in0(N__21822),
            .in1(N__24690),
            .in2(N__21802),
            .in3(N__21747),
            .lcout(n8_adj_1686),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i12_LC_3_8_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i12_LC_3_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i12_LC_3_8_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \RTD.read_buf_i12_LC_3_8_1  (
            .in0(N__21706),
            .in1(N__24087),
            .in2(N__21681),
            .in3(N__23985),
            .lcout(read_buf_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35044),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i13_LC_3_8_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i13_LC_3_8_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i13_LC_3_8_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.read_buf_i13_LC_3_8_2  (
            .in0(N__23984),
            .in1(N__21677),
            .in2(N__21886),
            .in3(N__24089),
            .lcout(read_buf_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35044),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i14_LC_3_8_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i14_LC_3_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i14_LC_3_8_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \RTD.read_buf_i14_LC_3_8_3  (
            .in0(N__21885),
            .in1(N__24088),
            .in2(N__21941),
            .in3(N__23986),
            .lcout(read_buf_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35044),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i3_LC_3_8_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i3_LC_3_8_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i3_LC_3_8_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i3_LC_3_8_5  (
            .in0(N__26493),
            .in1(N__21914),
            .in2(N__44247),
            .in3(N__23817),
            .lcout(buf_readRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35044),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i13_LC_3_8_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i13_LC_3_8_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i13_LC_3_8_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i13_LC_3_8_6  (
            .in0(N__21884),
            .in1(N__23814),
            .in2(N__31227),
            .in3(N__26494),
            .lcout(buf_readRTD_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35044),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_7_i19_3_lut_LC_3_9_1.C_ON=1'b0;
    defparam mux_127_Mux_7_i19_3_lut_LC_3_9_1.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_7_i19_3_lut_LC_3_9_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_7_i19_3_lut_LC_3_9_1 (
            .in0(N__25027),
            .in1(N__21984),
            .in2(_gnd_net_),
            .in3(N__59509),
            .lcout(),
            .ltout(n19_adj_1690_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_7_i22_3_lut_LC_3_9_2.C_ON=1'b0;
    defparam mux_127_Mux_7_i22_3_lut_LC_3_9_2.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_7_i22_3_lut_LC_3_9_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_127_Mux_7_i22_3_lut_LC_3_9_2 (
            .in0(_gnd_net_),
            .in1(N__22040),
            .in2(N__21868),
            .in3(N__60100),
            .lcout(n22_adj_1691),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i21_LC_3_9_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i21_LC_3_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i21_LC_3_9_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i21_LC_3_9_4  (
            .in0(N__35609),
            .in1(N__35865),
            .in2(N__23145),
            .in3(N__31196),
            .lcout(buf_adcdata_vac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61927),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_3_9_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_3_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_3_9_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i29_LC_3_9_6  (
            .in0(N__23138),
            .in1(N__33902),
            .in2(N__23008),
            .in3(N__35866),
            .lcout(cmd_rdadctmp_29_adj_1519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61927),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_6_i19_3_lut_LC_3_10_0.C_ON=1'b0;
    defparam mux_127_Mux_6_i19_3_lut_LC_3_10_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_6_i19_3_lut_LC_3_10_0.LUT_INIT=16'b1100101011001010;
    LogicCell40 mux_127_Mux_6_i19_3_lut_LC_3_10_0 (
            .in0(N__21857),
            .in1(N__25183),
            .in2(N__59518),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n19_adj_1693_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_6_i22_3_lut_LC_3_10_1.C_ON=1'b0;
    defparam mux_127_Mux_6_i22_3_lut_LC_3_10_1.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_6_i22_3_lut_LC_3_10_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_127_Mux_6_i22_3_lut_LC_3_10_1 (
            .in0(_gnd_net_),
            .in1(N__22061),
            .in2(N__21841),
            .in3(N__60099),
            .lcout(n22_adj_1694),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_5_i30_3_lut_LC_3_10_3.C_ON=1'b0;
    defparam mux_127_Mux_5_i30_3_lut_LC_3_10_3.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_5_i30_3_lut_LC_3_10_3.LUT_INIT=16'b1010110010101100;
    LogicCell40 mux_127_Mux_5_i30_3_lut_LC_3_10_3 (
            .in0(N__22081),
            .in1(N__22225),
            .in2(N__61057),
            .in3(_gnd_net_),
            .lcout(n30_adj_1698),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i6_LC_3_10_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i6_LC_3_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i6_LC_3_10_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i6_LC_3_10_4  (
            .in0(N__22062),
            .in1(N__39406),
            .in2(N__22024),
            .in3(N__39780),
            .lcout(buf_adcdata_iac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61944),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i7_LC_3_10_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i7_LC_3_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i7_LC_3_10_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i7_LC_3_10_5  (
            .in0(N__39775),
            .in1(N__22968),
            .in2(N__39418),
            .in3(N__22044),
            .lcout(buf_adcdata_iac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61944),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_3_10_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_3_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_3_10_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i14_LC_3_10_6  (
            .in0(N__22019),
            .in1(N__39776),
            .in2(N__22189),
            .in3(N__37831),
            .lcout(cmd_rdadctmp_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61944),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_3_10_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_3_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_3_10_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i15_LC_3_10_7  (
            .in0(N__37830),
            .in1(N__22020),
            .in2(N__39809),
            .in3(N__22967),
            .lcout(cmd_rdadctmp_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61944),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_4_i22_3_lut_LC_3_11_0.C_ON=1'b0;
    defparam mux_127_Mux_4_i22_3_lut_LC_3_11_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_4_i22_3_lut_LC_3_11_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_127_Mux_4_i22_3_lut_LC_3_11_0 (
            .in0(N__60083),
            .in1(N__21956),
            .in2(_gnd_net_),
            .in3(N__22009),
            .lcout(),
            .ltout(n22_adj_1701_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_4_i30_3_lut_LC_3_11_1.C_ON=1'b0;
    defparam mux_127_Mux_4_i30_3_lut_LC_3_11_1.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_4_i30_3_lut_LC_3_11_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_127_Mux_4_i30_3_lut_LC_3_11_1 (
            .in0(_gnd_net_),
            .in1(N__22003),
            .in2(N__21991),
            .in3(N__61017),
            .lcout(n30_adj_1702),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i7_LC_3_11_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i7_LC_3_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i7_LC_3_11_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i7_LC_3_11_2  (
            .in0(N__35601),
            .in1(N__35881),
            .in2(N__22219),
            .in3(N__21983),
            .lcout(buf_adcdata_vac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61962),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i4_LC_3_11_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i4_LC_3_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i4_LC_3_11_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i4_LC_3_11_4  (
            .in0(N__39386),
            .in1(N__39781),
            .in2(N__22686),
            .in3(N__21957),
            .lcout(buf_adcdata_iac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61962),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_5_i22_3_lut_LC_3_11_7.C_ON=1'b0;
    defparam mux_127_Mux_5_i22_3_lut_LC_3_11_7.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_5_i22_3_lut_LC_3_11_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_127_Mux_5_i22_3_lut_LC_3_11_7 (
            .in0(N__22157),
            .in1(N__22855),
            .in2(_gnd_net_),
            .in3(N__60082),
            .lcout(n22_adj_1697),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_3_12_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_3_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_3_12_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i13_LC_3_12_2  (
            .in0(N__22178),
            .in1(N__39819),
            .in2(N__22687),
            .in3(N__37832),
            .lcout(cmd_rdadctmp_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61978),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_3_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_3_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_3_12_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i16_LC_3_12_4  (
            .in0(N__22808),
            .in1(N__35867),
            .in2(N__22212),
            .in3(N__33939),
            .lcout(cmd_rdadctmp_16_adj_1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61978),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i5_LC_3_12_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i5_LC_3_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i5_LC_3_12_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i5_LC_3_12_6  (
            .in0(N__39399),
            .in1(N__39818),
            .in2(N__22185),
            .in3(N__22161),
            .lcout(buf_adcdata_iac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61978),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i8_LC_3_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i8_LC_3_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i8_LC_3_13_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i8_LC_3_13_0  (
            .in0(N__35587),
            .in1(N__35775),
            .in2(N__22818),
            .in3(N__25283),
            .lcout(buf_adcdata_vac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61991),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_3_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_3_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_3_13_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i23_LC_3_13_7  (
            .in0(N__35774),
            .in1(N__23040),
            .in2(N__24262),
            .in3(N__33981),
            .lcout(cmd_rdadctmp_23_adj_1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61991),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i3_3_lut_LC_3_14_0 .C_ON=1'b0;
    defparam \ADC_VAC.i3_3_lut_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i3_3_lut_LC_3_14_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \ADC_VAC.i3_3_lut_LC_3_14_0  (
            .in0(N__25876),
            .in1(N__32089),
            .in2(_gnd_net_),
            .in3(N__35712),
            .lcout(),
            .ltout(\ADC_VAC.n13747_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_LC_3_14_1 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_LC_3_14_1 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \ADC_VAC.i1_4_lut_LC_3_14_1  (
            .in0(N__31999),
            .in1(N__22138),
            .in2(N__22141),
            .in3(N__32090),
            .lcout(\ADC_VAC.n22030 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_LC_3_14_2 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_LC_3_14_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \ADC_VAC.i1_2_lut_LC_3_14_2  (
            .in0(N__22294),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35711),
            .lcout(\ADC_VAC.n13842 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19182_4_lut_LC_3_14_3 .C_ON=1'b0;
    defparam \ADC_VAC.i19182_4_lut_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19182_4_lut_LC_3_14_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i19182_4_lut_LC_3_14_3  (
            .in0(N__22131),
            .in1(N__22119),
            .in2(N__22108),
            .in3(N__22092),
            .lcout(),
            .ltout(\ADC_VAC.n22109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19199_4_lut_LC_3_14_4 .C_ON=1'b0;
    defparam \ADC_VAC.i19199_4_lut_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19199_4_lut_LC_3_14_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i19199_4_lut_LC_3_14_4  (
            .in0(N__22386),
            .in1(N__22374),
            .in2(N__22363),
            .in3(N__22359),
            .lcout(),
            .ltout(\ADC_VAC.n22126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i20123_4_lut_LC_3_14_5 .C_ON=1'b0;
    defparam \ADC_VAC.i20123_4_lut_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i20123_4_lut_LC_3_14_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_VAC.i20123_4_lut_LC_3_14_5  (
            .in0(N__35713),
            .in1(N__31991),
            .in2(N__22348),
            .in3(N__22344),
            .lcout(),
            .ltout(\ADC_VAC.n22389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i0_LC_3_14_6 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i0_LC_3_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i0_LC_3_14_6 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \ADC_VAC.adc_state_i0_LC_3_14_6  (
            .in0(N__32091),
            .in1(N__32000),
            .in2(N__22333),
            .in3(N__35714),
            .lcout(adc_state_0_adj_1516),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62000),
            .ce(N__22330),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i30_4_lut_LC_3_14_7 .C_ON=1'b0;
    defparam \ADC_VAC.i30_4_lut_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i30_4_lut_LC_3_14_7 .LUT_INIT=16'b1010100000001101;
    LogicCell40 \ADC_VAC.i30_4_lut_LC_3_14_7  (
            .in0(N__31998),
            .in1(N__22295),
            .in2(N__32100),
            .in3(N__25875),
            .lcout(\ADC_VAC.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_4_lut_LC_3_15_0 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_4_lut_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_4_lut_LC_3_15_0 .LUT_INIT=16'b0010001000000010;
    LogicCell40 \ADC_VAC.i1_2_lut_4_lut_LC_3_15_0  (
            .in0(N__31996),
            .in1(N__32066),
            .in2(N__22315),
            .in3(N__35709),
            .lcout(n13847),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i2_LC_3_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i2_LC_3_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i2_LC_3_15_2 .LUT_INIT=16'b0110011000100010;
    LogicCell40 \ADC_VAC.adc_state_i2_LC_3_15_2  (
            .in0(N__31997),
            .in1(N__32067),
            .in2(_gnd_net_),
            .in3(N__35710),
            .lcout(DTRIG_N_1182_adj_1549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62007),
            .ce(N__22266),
            .sr(_gnd_net_));
    defparam \RTD.CS_52_LC_5_2_0 .C_ON=1'b0;
    defparam \RTD.CS_52_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \RTD.CS_52_LC_5_2_0 .LUT_INIT=16'b0000110001011111;
    LogicCell40 \RTD.CS_52_LC_5_2_0  (
            .in0(N__26672),
            .in1(N__22231),
            .in2(N__26855),
            .in3(N__26206),
            .lcout(RTD_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35014),
            .ce(N__23377),
            .sr(_gnd_net_));
    defparam \RTD.i19756_2_lut_LC_5_3_3 .C_ON=1'b0;
    defparam \RTD.i19756_2_lut_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i19756_2_lut_LC_5_3_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \RTD.i19756_2_lut_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__23345),
            .in2(_gnd_net_),
            .in3(N__23689),
            .lcout(\RTD.n22382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_rep_43_2_lut_3_lut_LC_5_4_1 .C_ON=1'b0;
    defparam \RTD.i1_rep_43_2_lut_3_lut_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_rep_43_2_lut_3_lut_LC_5_4_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \RTD.i1_rep_43_2_lut_3_lut_LC_5_4_1  (
            .in0(N__35128),
            .in1(N__26646),
            .in2(_gnd_net_),
            .in3(N__32872),
            .lcout(\RTD.n23689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_21_LC_5_4_2 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_21_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_21_LC_5_4_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \RTD.i1_2_lut_adj_21_LC_5_4_2  (
            .in0(N__32873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35129),
            .lcout(\RTD.n20051 ),
            .ltout(\RTD.n20051_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i20050_3_lut_4_lut_LC_5_4_3 .C_ON=1'b0;
    defparam \RTD.i20050_3_lut_4_lut_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i20050_3_lut_4_lut_LC_5_4_3 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \RTD.i20050_3_lut_4_lut_LC_5_4_3  (
            .in0(N__22402),
            .in1(N__23202),
            .in2(N__22447),
            .in3(N__26798),
            .lcout(),
            .ltout(\RTD.n22599_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i3_LC_5_4_4 .C_ON=1'b0;
    defparam \RTD.adc_state_i3_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i3_LC_5_4_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \RTD.adc_state_i3_LC_5_4_4  (
            .in0(N__22444),
            .in1(N__26393),
            .in2(N__22432),
            .in3(N__22428),
            .lcout(\RTD.adc_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34980),
            .ce(N__23272),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i2_LC_5_4_5 .C_ON=1'b0;
    defparam \RTD.adc_state_i2_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i2_LC_5_4_5 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \RTD.adc_state_i2_LC_5_4_5  (
            .in0(N__22393),
            .in1(N__23462),
            .in2(N__24940),
            .in3(N__26394),
            .lcout(adc_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34980),
            .ce(N__23272),
            .sr(_gnd_net_));
    defparam \RTD.i1_3_lut_4_lut_LC_5_4_6 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_4_lut_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_4_lut_LC_5_4_6 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \RTD.i1_3_lut_4_lut_LC_5_4_6  (
            .in0(N__32874),
            .in1(N__35130),
            .in2(N__26673),
            .in3(N__26799),
            .lcout(),
            .ltout(\RTD.n56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i0_LC_5_4_7 .C_ON=1'b0;
    defparam \RTD.adc_state_i0_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i0_LC_5_4_7 .LUT_INIT=16'b0101011100010011;
    LogicCell40 \RTD.adc_state_i0_LC_5_4_7  (
            .in0(N__26392),
            .in1(N__26165),
            .in2(N__22414),
            .in3(N__22411),
            .lcout(\RTD.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34980),
            .ce(N__23272),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_23_LC_5_5_2 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_23_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_23_LC_5_5_2 .LUT_INIT=16'b1100000010001101;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_23_LC_5_5_2  (
            .in0(N__26145),
            .in1(N__26785),
            .in2(N__26459),
            .in3(N__26605),
            .lcout(n13584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_26_LC_5_5_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_26_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_26_LC_5_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RTD.i1_2_lut_adj_26_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(N__26604),
            .in2(_gnd_net_),
            .in3(N__26144),
            .lcout(\RTD.n71 ),
            .ltout(\RTD.n71_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i20122_3_lut_4_lut_LC_5_5_6 .C_ON=1'b0;
    defparam \RTD.i20122_3_lut_4_lut_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i20122_3_lut_4_lut_LC_5_5_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \RTD.i20122_3_lut_4_lut_LC_5_5_6  (
            .in0(N__22546),
            .in1(N__23200),
            .in2(N__22396),
            .in3(N__26786),
            .lcout(\RTD.n22623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_LC_5_5_7 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_LC_5_5_7 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \RTD.i1_4_lut_LC_5_5_7  (
            .in0(N__26606),
            .in1(N__22545),
            .in2(N__26839),
            .in3(N__26146),
            .lcout(\RTD.n62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i4_LC_5_6_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i4_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i4_LC_5_6_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i4_LC_5_6_0  (
            .in0(N__23780),
            .in1(N__22515),
            .in2(N__30882),
            .in3(N__26437),
            .lcout(buf_readRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35021),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i0_LC_5_6_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i0_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i0_LC_5_6_1 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i0_LC_5_6_1  (
            .in0(N__26434),
            .in1(N__22537),
            .in2(N__25524),
            .in3(N__23781),
            .lcout(buf_readRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35021),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_adj_24_LC_5_6_2 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_adj_24_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_adj_24_LC_5_6_2 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \RTD.i1_2_lut_3_lut_adj_24_LC_5_6_2  (
            .in0(N__26181),
            .in1(N__26433),
            .in2(_gnd_net_),
            .in3(N__26817),
            .lcout(n21989),
            .ltout(n21989_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i5_LC_5_6_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i5_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i5_LC_5_6_3 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \RTD.read_buf_i5_LC_5_6_3  (
            .in0(N__23939),
            .in1(N__22516),
            .in2(N__22495),
            .in3(N__23291),
            .lcout(read_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35021),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i2_LC_5_6_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i2_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i2_LC_5_6_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \RTD.read_buf_i2_LC_5_6_4  (
            .in0(N__22492),
            .in1(N__24037),
            .in2(N__22467),
            .in3(N__23940),
            .lcout(read_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35021),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i1_LC_5_6_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i1_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i1_LC_5_6_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i1_LC_5_6_5  (
            .in0(N__26435),
            .in1(N__22491),
            .in2(N__22722),
            .in3(N__23782),
            .lcout(buf_readRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35021),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i6_LC_5_6_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i6_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i6_LC_5_6_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \RTD.read_buf_i6_LC_5_6_6  (
            .in0(N__23292),
            .in1(N__23941),
            .in2(N__24067),
            .in3(N__24107),
            .lcout(read_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35021),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i2_LC_5_6_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i2_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i2_LC_5_6_7 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i2_LC_5_6_7  (
            .in0(N__26436),
            .in1(N__22463),
            .in2(N__24339),
            .in3(N__23783),
            .lcout(buf_readRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35021),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i2_LC_5_7_0 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i2_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i2_LC_5_7_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i2_LC_5_7_0  (
            .in0(N__23459),
            .in1(N__23503),
            .in2(N__28965),
            .in3(N__22582),
            .lcout(\RTD.cfg_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35034),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i4_LC_5_7_1 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i4_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i4_LC_5_7_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.cfg_buf_i4_LC_5_7_1  (
            .in0(N__23505),
            .in1(N__23461),
            .in2(N__28924),
            .in3(N__22591),
            .lcout(\RTD.cfg_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35034),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_20_LC_5_7_2 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_20_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_20_LC_5_7_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \RTD.i1_2_lut_adj_20_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__26185),
            .in2(_gnd_net_),
            .in3(N__26818),
            .lcout(\RTD.n68 ),
            .ltout(\RTD.n68_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i0_LC_5_7_3 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i0_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i0_LC_5_7_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.cfg_buf_i0_LC_5_7_3  (
            .in0(N__23502),
            .in1(N__48719),
            .in2(N__22594),
            .in3(N__22573),
            .lcout(\RTD.cfg_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35034),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_4_lut_LC_5_7_4 .C_ON=1'b0;
    defparam \RTD.i2_4_lut_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_4_lut_LC_5_7_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i2_4_lut_LC_5_7_4  (
            .in0(N__22590),
            .in1(N__22581),
            .in2(N__28966),
            .in3(N__28922),
            .lcout(\RTD.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_30_LC_5_7_5 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_30_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_30_LC_5_7_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i1_4_lut_adj_30_LC_5_7_5  (
            .in0(N__48720),
            .in1(N__22554),
            .in2(N__25225),
            .in3(N__22572),
            .lcout(),
            .ltout(\RTD.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i7_4_lut_LC_5_7_6 .C_ON=1'b0;
    defparam \RTD.i7_4_lut_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i7_4_lut_LC_5_7_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \RTD.i7_4_lut_LC_5_7_6  (
            .in0(N__23536),
            .in1(N__22564),
            .in2(N__22558),
            .in3(N__23260),
            .lcout(\RTD.adress_7_N_1009_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i3_LC_5_7_7 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i3_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i3_LC_5_7_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.cfg_buf_i3_LC_5_7_7  (
            .in0(N__23504),
            .in1(N__23460),
            .in2(N__25224),
            .in3(N__22555),
            .lcout(\RTD.cfg_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35034),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i0_LC_5_8_0 .C_ON=1'b0;
    defparam \RTD.adress_i0_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i0_LC_5_8_0 .LUT_INIT=16'b1011000111110101;
    LogicCell40 \RTD.adress_i0_LC_5_8_0  (
            .in0(N__26670),
            .in1(N__26253),
            .in2(N__22653),
            .in3(N__23685),
            .lcout(\RTD.adress_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35022),
            .ce(N__24160),
            .sr(N__22630));
    defparam \RTD.adress_i7_LC_5_8_1 .C_ON=1'b0;
    defparam \RTD.adress_i7_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i7_LC_5_8_1 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.adress_i7_LC_5_8_1  (
            .in0(N__23686),
            .in1(N__23598),
            .in2(N__26257),
            .in3(N__26671),
            .lcout(\RTD.adress_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35022),
            .ce(N__24160),
            .sr(N__22630));
    defparam \RTD.i34_3_lut_4_lut_LC_5_8_2 .C_ON=1'b0;
    defparam \RTD.i34_3_lut_4_lut_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i34_3_lut_4_lut_LC_5_8_2 .LUT_INIT=16'b1101110110001101;
    LogicCell40 \RTD.i34_3_lut_4_lut_LC_5_8_2  (
            .in0(N__26668),
            .in1(N__26252),
            .in2(N__23363),
            .in3(N__23648),
            .lcout(),
            .ltout(\RTD.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i35_4_lut_LC_5_8_3 .C_ON=1'b0;
    defparam \RTD.i35_4_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i35_4_lut_LC_5_8_3 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \RTD.i35_4_lut_LC_5_8_3  (
            .in0(N__26431),
            .in1(N__22624),
            .in2(N__22633),
            .in3(N__26856),
            .lcout(\RTD.n13441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19113_2_lut_3_lut_4_lut_LC_5_8_4 .C_ON=1'b0;
    defparam \RTD.i19113_2_lut_3_lut_4_lut_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i19113_2_lut_3_lut_4_lut_LC_5_8_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \RTD.i19113_2_lut_3_lut_4_lut_LC_5_8_4  (
            .in0(N__26669),
            .in1(N__26432),
            .in2(N__26248),
            .in3(N__26854),
            .lcout(\RTD.n15396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_LC_5_8_6 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_LC_5_8_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \RTD.i1_2_lut_3_lut_LC_5_8_6  (
            .in0(N__26667),
            .in1(N__26430),
            .in2(_gnd_net_),
            .in3(N__26251),
            .lcout(\RTD.n1 ),
            .ltout(\RTD.n1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i22_4_lut_LC_5_8_7 .C_ON=1'b0;
    defparam \RTD.i22_4_lut_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i22_4_lut_LC_5_8_7 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \RTD.i22_4_lut_LC_5_8_7  (
            .in0(N__23649),
            .in1(N__23386),
            .in2(N__22618),
            .in3(N__26857),
            .lcout(\RTD.n13482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_tmp_i0_LC_5_9_0 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i0_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i0_LC_5_9_0 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \RTD.cfg_tmp_i0_LC_5_9_0  (
            .in0(N__26186),
            .in1(N__26499),
            .in2(N__48724),
            .in3(N__22758),
            .lcout(\RTD.cfg_tmp_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam \RTD.cfg_tmp_i1_LC_5_9_1 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i1_LC_5_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i1_LC_5_9_1 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \RTD.cfg_tmp_i1_LC_5_9_1  (
            .in0(N__22615),
            .in1(N__26190),
            .in2(N__38245),
            .in3(N__26495),
            .lcout(\RTD.cfg_tmp_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam \RTD.cfg_tmp_i2_LC_5_9_2 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i2_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i2_LC_5_9_2 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \RTD.cfg_tmp_i2_LC_5_9_2  (
            .in0(N__26187),
            .in1(N__26500),
            .in2(N__22609),
            .in3(N__28953),
            .lcout(\RTD.cfg_tmp_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam \RTD.cfg_tmp_i3_LC_5_9_3 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i3_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i3_LC_5_9_3 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.cfg_tmp_i3_LC_5_9_3  (
            .in0(N__26496),
            .in1(N__22600),
            .in2(N__25217),
            .in3(N__26193),
            .lcout(\RTD.cfg_tmp_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam \RTD.cfg_tmp_i4_LC_5_9_4 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i4_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i4_LC_5_9_4 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \RTD.cfg_tmp_i4_LC_5_9_4  (
            .in0(N__26188),
            .in1(N__26501),
            .in2(N__28923),
            .in3(N__22792),
            .lcout(\RTD.cfg_tmp_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam \RTD.cfg_tmp_i5_LC_5_9_5 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i5_LC_5_9_5 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i5_LC_5_9_5 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i5_LC_5_9_5  (
            .in0(N__26497),
            .in1(N__26191),
            .in2(N__31177),
            .in3(N__22786),
            .lcout(\RTD.cfg_tmp_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam \RTD.cfg_tmp_i6_LC_5_9_6 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i6_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i6_LC_5_9_6 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \RTD.cfg_tmp_i6_LC_5_9_6  (
            .in0(N__26189),
            .in1(N__26502),
            .in2(N__29011),
            .in3(N__22780),
            .lcout(\RTD.cfg_tmp_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam \RTD.cfg_tmp_i7_LC_5_9_7 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i7_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i7_LC_5_9_7 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i7_LC_5_9_7  (
            .in0(N__26498),
            .in1(N__26192),
            .in2(N__35362),
            .in3(N__22774),
            .lcout(\RTD.cfg_tmp_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35043),
            .ce(N__23632),
            .sr(N__23617));
    defparam mux_127_Mux_6_i30_3_lut_LC_5_10_0.C_ON=1'b0;
    defparam mux_127_Mux_6_i30_3_lut_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_6_i30_3_lut_LC_5_10_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_6_i30_3_lut_LC_5_10_0 (
            .in0(N__22747),
            .in1(N__22735),
            .in2(_gnd_net_),
            .in3(N__61051),
            .lcout(n30_adj_1695),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_5_10_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_5_10_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i26_LC_5_10_2  (
            .in0(N__33985),
            .in1(N__25124),
            .in2(N__31551),
            .in3(N__35964),
            .lcout(cmd_rdadctmp_26_adj_1522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61909),
            .ce(),
            .sr(_gnd_net_));
    defparam i19210_3_lut_LC_5_10_3.C_ON=1'b0;
    defparam i19210_3_lut_LC_5_10_3.SEQ_MODE=4'b0000;
    defparam i19210_3_lut_LC_5_10_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i19210_3_lut_LC_5_10_3 (
            .in0(N__22726),
            .in1(N__23842),
            .in2(_gnd_net_),
            .in3(N__60669),
            .lcout(n22137),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_5_10_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_5_10_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i3_LC_5_10_6  (
            .in0(N__33986),
            .in1(N__22705),
            .in2(N__31357),
            .in3(N__35965),
            .lcout(cmd_rdadctmp_3_adj_1545),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61909),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_5_11_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_5_11_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i12_LC_5_11_0  (
            .in0(N__39800),
            .in1(N__22670),
            .in2(N__35395),
            .in3(N__37801),
            .lcout(cmd_rdadctmp_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61928),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_5_11_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_5_11_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i19_LC_5_11_1  (
            .in0(N__28805),
            .in1(N__33988),
            .in2(N__22881),
            .in3(N__36007),
            .lcout(cmd_rdadctmp_19_adj_1529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61928),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i16_LC_5_11_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i16_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i16_LC_5_11_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i16_LC_5_11_2  (
            .in0(N__36003),
            .in1(N__35599),
            .in2(N__23029),
            .in3(N__43496),
            .lcout(buf_adcdata_vac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61928),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i10_LC_5_11_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i10_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i10_LC_5_11_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i10_LC_5_11_3  (
            .in0(N__35598),
            .in1(N__36005),
            .in2(N__22882),
            .in3(N__25077),
            .lcout(buf_adcdata_vac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61928),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i9_LC_5_11_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i9_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i9_LC_5_11_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i9_LC_5_11_4  (
            .in0(N__36004),
            .in1(N__35600),
            .in2(N__23868),
            .in3(N__22896),
            .lcout(buf_adcdata_vac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61928),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_5_i19_3_lut_LC_5_11_5.C_ON=1'b0;
    defparam mux_127_Mux_5_i19_3_lut_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_5_i19_3_lut_LC_5_11_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_5_i19_3_lut_LC_5_11_5 (
            .in0(N__28216),
            .in1(N__22926),
            .in2(_gnd_net_),
            .in3(N__59111),
            .lcout(n19_adj_1696),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_7_i30_3_lut_LC_5_11_6.C_ON=1'b0;
    defparam mux_127_Mux_7_i30_3_lut_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_7_i30_3_lut_LC_5_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_7_i30_3_lut_LC_5_11_6 (
            .in0(N__22846),
            .in1(N__22834),
            .in2(_gnd_net_),
            .in3(N__61052),
            .lcout(n30_adj_1692),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_5_11_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_5_11_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i17_LC_5_11_7  (
            .in0(N__22895),
            .in1(N__33987),
            .in2(N__22822),
            .in3(N__36006),
            .lcout(cmd_rdadctmp_17_adj_1531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61928),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_5_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_5_12_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i28_LC_5_12_0  (
            .in0(N__36010),
            .in1(N__22994),
            .in2(N__27861),
            .in3(N__33937),
            .lcout(cmd_rdadctmp_28_adj_1520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61945),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_5_12_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_5_12_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i27_LC_5_12_3  (
            .in0(N__33934),
            .in1(N__27854),
            .in2(N__25137),
            .in3(N__36012),
            .lcout(cmd_rdadctmp_27_adj_1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61945),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_5_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_5_12_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i24_LC_5_12_4  (
            .in0(N__36008),
            .in1(N__23021),
            .in2(N__23053),
            .in3(N__33935),
            .lcout(cmd_rdadctmp_24_adj_1524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61945),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i15_LC_5_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i15_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i15_LC_5_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i15_LC_5_12_5  (
            .in0(N__35567),
            .in1(N__36011),
            .in2(N__24228),
            .in3(N__23052),
            .lcout(buf_adcdata_vac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61945),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_5_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_5_12_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i25_LC_5_12_6  (
            .in0(N__36009),
            .in1(N__23022),
            .in2(N__31547),
            .in3(N__33936),
            .lcout(cmd_rdadctmp_25_adj_1523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61945),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i20_LC_5_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i20_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i20_LC_5_13_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i20_LC_5_13_0  (
            .in0(N__35565),
            .in1(N__35922),
            .in2(N__23004),
            .in3(N__25446),
            .lcout(buf_adcdata_vac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61963),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_5_13_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_5_13_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i16_LC_5_13_1  (
            .in0(N__34589),
            .in1(N__39728),
            .in2(N__22978),
            .in3(N__37810),
            .lcout(cmd_rdadctmp_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61963),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i5_LC_5_13_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i5_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i5_LC_5_13_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i5_LC_5_13_5  (
            .in0(N__35921),
            .in1(N__35566),
            .in2(N__22954),
            .in3(N__22925),
            .lcout(buf_adcdata_vac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61963),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_5_14_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_5_14_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i18_LC_5_14_0  (
            .in0(N__22869),
            .in1(N__33950),
            .in2(N__22903),
            .in3(N__35854),
            .lcout(cmd_rdadctmp_18_adj_1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61979),
            .ce(),
            .sr(_gnd_net_));
    defparam n23540_bdd_4_lut_LC_5_14_5.C_ON=1'b0;
    defparam n23540_bdd_4_lut_LC_5_14_5.SEQ_MODE=4'b0000;
    defparam n23540_bdd_4_lut_LC_5_14_5.LUT_INIT=16'b1100110010111000;
    LogicCell40 n23540_bdd_4_lut_LC_5_14_5 (
            .in0(N__25348),
            .in1(N__25411),
            .in2(N__32203),
            .in3(N__60670),
            .lcout(),
            .ltout(n23543_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19349_3_lut_LC_5_14_6.C_ON=1'b0;
    defparam i19349_3_lut_LC_5_14_6.SEQ_MODE=4'b0000;
    defparam i19349_3_lut_LC_5_14_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 i19349_3_lut_LC_5_14_6 (
            .in0(_gnd_net_),
            .in1(N__23215),
            .in2(N__22858),
            .in3(N__60096),
            .lcout(n22276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_5_15_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_5_15_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i31_LC_5_15_1  (
            .in0(N__23160),
            .in1(N__33952),
            .in2(N__23125),
            .in3(N__35917),
            .lcout(cmd_rdadctmp_31_adj_1517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61992),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i23_LC_5_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i23_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i23_LC_5_15_2 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i23_LC_5_15_2  (
            .in0(N__35914),
            .in1(N__23161),
            .in2(N__35571),
            .in3(N__23237),
            .lcout(buf_adcdata_vac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61992),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_5_15_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_5_15_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i30_LC_5_15_3  (
            .in0(N__23152),
            .in1(N__33951),
            .in2(N__23124),
            .in3(N__35916),
            .lcout(cmd_rdadctmp_30_adj_1518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61992),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_83_LC_5_15_4.C_ON=1'b0;
    defparam i1_2_lut_adj_83_LC_5_15_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_83_LC_5_15_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_83_LC_5_15_4 (
            .in0(_gnd_net_),
            .in1(N__32004),
            .in2(_gnd_net_),
            .in3(N__32072),
            .lcout(n21948),
            .ltout(n21948_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i22_LC_5_15_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i22_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i22_LC_5_15_5 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i22_LC_5_15_5  (
            .in0(N__23123),
            .in1(N__35915),
            .in2(N__23107),
            .in3(N__23091),
            .lcout(buf_adcdata_vac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61992),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_6_i19_3_lut_LC_5_16_5.C_ON=1'b0;
    defparam mux_125_Mux_6_i19_3_lut_LC_5_16_5.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_6_i19_3_lut_LC_5_16_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_6_i19_3_lut_LC_5_16_5 (
            .in0(N__25162),
            .in1(N__23087),
            .in2(_gnd_net_),
            .in3(N__59515),
            .lcout(n19_adj_1765),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_I_0_1_lut_LC_5_19_3.C_ON=1'b0;
    defparam acadc_rst_I_0_1_lut_LC_5_19_3.SEQ_MODE=4'b0000;
    defparam acadc_rst_I_0_1_lut_LC_5_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 acadc_rst_I_0_1_lut_LC_5_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39177),
            .lcout(AC_ADC_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_4_lut_LC_6_4_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_4_lut_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_4_lut_LC_6_4_5 .LUT_INIT=16'b1011011011000110;
    LogicCell40 \RTD.i1_2_lut_4_lut_LC_6_4_5  (
            .in0(N__26771),
            .in1(N__26653),
            .in2(N__26398),
            .in3(N__26174),
            .lcout(\RTD.n18274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_22_LC_6_5_0 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_22_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_22_LC_6_5_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \RTD.i1_2_lut_adj_22_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__26372),
            .in2(_gnd_net_),
            .in3(N__26117),
            .lcout(\RTD.n21988 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_2_lut_LC_6_5_1 .C_ON=1'b0;
    defparam \RTD.i2_2_lut_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_2_lut_LC_6_5_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i2_2_lut_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__26608),
            .in2(_gnd_net_),
            .in3(N__23688),
            .lcout(),
            .ltout(\RTD.n7_adj_1497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4_4_lut_LC_6_5_2 .C_ON=1'b0;
    defparam \RTD.i4_4_lut_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i4_4_lut_LC_6_5_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \RTD.i4_4_lut_LC_6_5_2  (
            .in0(N__23364),
            .in1(N__23305),
            .in2(N__23299),
            .in3(N__26791),
            .lcout(\RTD.n12274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i6_LC_6_5_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i6_LC_6_5_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i6_LC_6_5_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i6_LC_6_5_5  (
            .in0(N__26375),
            .in1(N__43671),
            .in2(N__24114),
            .in3(N__23779),
            .lcout(buf_readRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34956),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_LC_6_5_6 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_LC_6_5_6 .LUT_INIT=16'b1100100010000000;
    LogicCell40 \RTD.i1_4_lut_4_lut_LC_6_5_6  (
            .in0(N__26607),
            .in1(N__26790),
            .in2(N__26224),
            .in3(N__26373),
            .lcout(n13603),
            .ltout(n13603_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i5_LC_6_5_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i5_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i5_LC_6_5_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \RTD.READ_DATA_i5_LC_6_5_7  (
            .in0(N__26374),
            .in1(N__38004),
            .in2(N__23296),
            .in3(N__23293),
            .lcout(buf_readRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34956),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i1_LC_6_6_0 .C_ON=1'b0;
    defparam \RTD.adc_state_i1_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i1_LC_6_6_0 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \RTD.adc_state_i1_LC_6_6_0  (
            .in0(N__23458),
            .in1(N__23515),
            .in2(N__26517),
            .in3(N__23278),
            .lcout(\RTD.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35002),
            .ce(N__23271),
            .sr(_gnd_net_));
    defparam \RTD.i3_4_lut_LC_6_6_3 .C_ON=1'b0;
    defparam \RTD.i3_4_lut_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i3_4_lut_LC_6_6_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i3_4_lut_LC_6_6_3  (
            .in0(N__23526),
            .in1(N__23415),
            .in2(N__35354),
            .in3(N__38238),
            .lcout(\RTD.n11_adj_1500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23432_bdd_4_lut_LC_6_6_5.C_ON=1'b0;
    defparam n23432_bdd_4_lut_LC_6_6_5.SEQ_MODE=4'b0000;
    defparam n23432_bdd_4_lut_LC_6_6_5.LUT_INIT=16'b1100110011100010;
    LogicCell40 n23432_bdd_4_lut_LC_6_6_5 (
            .in0(N__23250),
            .in1(N__35287),
            .in2(N__25009),
            .in3(N__60649),
            .lcout(n23435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.mode_53_LC_6_7_0 .C_ON=1'b0;
    defparam \RTD.mode_53_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.mode_53_LC_6_7_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \RTD.mode_53_LC_6_7_0  (
            .in0(N__23464),
            .in1(N__23311),
            .in2(N__23201),
            .in3(N__23687),
            .lcout(\RTD.mode ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35029),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i6_LC_6_7_1 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i6_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i6_LC_6_7_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.cfg_buf_i6_LC_6_7_1  (
            .in0(N__23554),
            .in1(N__29009),
            .in2(N__23476),
            .in3(N__23509),
            .lcout(\RTD.cfg_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35029),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i5_LC_6_7_2 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i5_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i5_LC_6_7_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.cfg_buf_i5_LC_6_7_2  (
            .in0(N__23545),
            .in1(N__31159),
            .in2(N__23474),
            .in3(N__23507),
            .lcout(\RTD.cfg_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35029),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4_4_lut_adj_29_LC_6_7_3 .C_ON=1'b0;
    defparam \RTD.i4_4_lut_adj_29_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i4_4_lut_adj_29_LC_6_7_3 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i4_4_lut_adj_29_LC_6_7_3  (
            .in0(N__23553),
            .in1(N__29010),
            .in2(N__31169),
            .in3(N__23544),
            .lcout(\RTD.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i1_LC_6_7_4 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i1_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i1_LC_6_7_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \RTD.cfg_buf_i1_LC_6_7_4  (
            .in0(N__23463),
            .in1(N__23506),
            .in2(N__23530),
            .in3(N__38237),
            .lcout(\RTD.cfg_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35029),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i17375_3_lut_LC_6_7_5 .C_ON=1'b0;
    defparam \RTD.i17375_3_lut_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i17375_3_lut_LC_6_7_5 .LUT_INIT=16'b0101010100100010;
    LogicCell40 \RTD.i17375_3_lut_LC_6_7_5  (
            .in0(N__26609),
            .in1(N__26863),
            .in2(_gnd_net_),
            .in3(N__26225),
            .lcout(\RTD.n20093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i7_LC_6_7_6 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i7_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i7_LC_6_7_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \RTD.cfg_buf_i7_LC_6_7_6  (
            .in0(N__23416),
            .in1(N__23508),
            .in2(N__23475),
            .in3(N__35355),
            .lcout(\RTD.cfg_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35029),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i14786_3_lut_LC_6_7_7 .C_ON=1'b0;
    defparam \RTD.i14786_3_lut_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i14786_3_lut_LC_6_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \RTD.i14786_3_lut_LC_6_7_7  (
            .in0(N__23404),
            .in1(N__29008),
            .in2(_gnd_net_),
            .in3(N__59246),
            .lcout(n20_adj_1766),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_28_LC_6_8_0 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_28_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_28_LC_6_8_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \RTD.i1_2_lut_adj_28_LC_6_8_0  (
            .in0(N__26617),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26473),
            .lcout(\RTD.n68_adj_1498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i20131_3_lut_3_lut_LC_6_8_1 .C_ON=1'b0;
    defparam \RTD.i20131_3_lut_3_lut_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i20131_3_lut_3_lut_LC_6_8_1 .LUT_INIT=16'b1010000110100001;
    LogicCell40 \RTD.i20131_3_lut_3_lut_LC_6_8_1  (
            .in0(N__26474),
            .in1(N__26618),
            .in2(N__26865),
            .in3(_gnd_net_),
            .lcout(\RTD.n21954 ),
            .ltout(\RTD.n21954_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_3_lut_4_lut_adj_31_LC_6_8_2 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_4_lut_adj_31_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_4_lut_adj_31_LC_6_8_2 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \RTD.i1_3_lut_4_lut_adj_31_LC_6_8_2  (
            .in0(N__23365),
            .in1(N__26853),
            .in2(N__23314),
            .in3(N__23650),
            .lcout(\RTD.n21955 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i5_LC_6_8_3.C_ON=1'b0;
    defparam buf_cfgRTD_i5_LC_6_8_3.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i5_LC_6_8_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i5_LC_6_8_3 (
            .in0(N__57621),
            .in1(N__48810),
            .in2(N__45340),
            .in3(N__31158),
            .lcout(buf_cfgRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61861),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_25_LC_6_8_4 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_25_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_25_LC_6_8_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \RTD.i1_2_lut_adj_25_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__26250),
            .in2(_gnd_net_),
            .in3(N__23678),
            .lcout(\RTD.n11 ),
            .ltout(\RTD.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i30_4_lut_LC_6_8_5 .C_ON=1'b0;
    defparam \RTD.i30_4_lut_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i30_4_lut_LC_6_8_5 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \RTD.i30_4_lut_LC_6_8_5  (
            .in0(N__26475),
            .in1(N__24946),
            .in2(N__23635),
            .in3(N__23605),
            .lcout(\RTD.n13488 ),
            .ltout(\RTD.n13488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12862_2_lut_LC_6_8_6 .C_ON=1'b0;
    defparam \RTD.i12862_2_lut_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i12862_2_lut_LC_6_8_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \RTD.i12862_2_lut_LC_6_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23620),
            .in3(N__26852),
            .lcout(\RTD.n15585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19155_2_lut_LC_6_8_7 .C_ON=1'b0;
    defparam \RTD.i19155_2_lut_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i19155_2_lut_LC_6_8_7 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \RTD.i19155_2_lut_LC_6_8_7  (
            .in0(N__26848),
            .in1(N__26616),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RTD.n22081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i6_LC_6_9_0 .C_ON=1'b0;
    defparam \RTD.adress_i6_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i6_LC_6_9_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.adress_i6_LC_6_9_0  (
            .in0(N__24159),
            .in1(N__23583),
            .in2(N__23599),
            .in3(N__24929),
            .lcout(\RTD.adress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35000),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i5_LC_6_9_1 .C_ON=1'b0;
    defparam \RTD.adress_i5_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i5_LC_6_9_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i5_LC_6_9_1  (
            .in0(N__23584),
            .in1(N__24924),
            .in2(N__23575),
            .in3(N__24158),
            .lcout(\RTD.adress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35000),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i4_LC_6_9_2 .C_ON=1'b0;
    defparam \RTD.adress_i4_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i4_LC_6_9_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.adress_i4_LC_6_9_2  (
            .in0(N__24157),
            .in1(N__23574),
            .in2(N__24933),
            .in3(N__23563),
            .lcout(\RTD.adress_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35000),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i3_LC_6_9_3 .C_ON=1'b0;
    defparam \RTD.adress_i3_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i3_LC_6_9_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i3_LC_6_9_3  (
            .in0(N__23562),
            .in1(N__24923),
            .in2(N__24181),
            .in3(N__24156),
            .lcout(\RTD.adress_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35000),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i2_LC_6_9_4 .C_ON=1'b0;
    defparam \RTD.adress_i2_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i2_LC_6_9_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.adress_i2_LC_6_9_4  (
            .in0(N__24155),
            .in1(N__24180),
            .in2(N__24133),
            .in3(N__24928),
            .lcout(\RTD.adress_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35000),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i9_LC_6_9_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i9_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i9_LC_6_9_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \RTD.read_buf_i9_LC_6_9_6  (
            .in0(N__23835),
            .in1(N__24052),
            .in2(N__23714),
            .in3(N__23974),
            .lcout(read_buf_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35000),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i1_LC_6_9_7 .C_ON=1'b0;
    defparam \RTD.adress_i1_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i1_LC_6_9_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i1_LC_6_9_7  (
            .in0(N__24132),
            .in1(N__24922),
            .in2(N__24169),
            .in3(N__24154),
            .lcout(\RTD.adress_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35000),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i8_LC_6_10_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i8_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i8_LC_6_10_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.read_buf_i8_LC_6_10_0  (
            .in0(N__23977),
            .in1(N__23892),
            .in2(N__23836),
            .in3(N__24077),
            .lcout(read_buf_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35001),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i7_LC_6_10_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i7_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i7_LC_6_10_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \RTD.read_buf_i7_LC_6_10_1  (
            .in0(N__24118),
            .in1(N__24076),
            .in2(N__23893),
            .in3(N__23978),
            .lcout(read_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35001),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i7_LC_6_10_2 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i7_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i7_LC_6_10_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \RTD.READ_DATA_i7_LC_6_10_2  (
            .in0(N__24192),
            .in1(N__23891),
            .in2(N__23812),
            .in3(N__26515),
            .lcout(buf_readRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35001),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_1_i19_3_lut_LC_6_10_3.C_ON=1'b0;
    defparam mux_126_Mux_1_i19_3_lut_LC_6_10_3.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_1_i19_3_lut_LC_6_10_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_1_i19_3_lut_LC_6_10_3 (
            .in0(N__24961),
            .in1(N__23861),
            .in2(_gnd_net_),
            .in3(N__59466),
            .lcout(n19_adj_1752),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i8_LC_6_10_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i8_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i8_LC_6_10_5 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \RTD.READ_DATA_i8_LC_6_10_5  (
            .in0(N__26514),
            .in1(N__23834),
            .in2(N__23813),
            .in3(N__43305),
            .lcout(buf_readRTD_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35001),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i9_LC_6_10_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i9_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i9_LC_6_10_6 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i9_LC_6_10_6  (
            .in0(N__38256),
            .in1(N__23792),
            .in2(N__23715),
            .in3(N__26516),
            .lcout(buf_readRTD_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35001),
            .ce(),
            .sr(_gnd_net_));
    defparam i19222_3_lut_LC_6_11_1.C_ON=1'b0;
    defparam i19222_3_lut_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam i19222_3_lut_LC_6_11_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i19222_3_lut_LC_6_11_1 (
            .in0(N__60619),
            .in1(N__24343),
            .in2(_gnd_net_),
            .in3(N__25051),
            .lcout(n22149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_6_11_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_6_11_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i12_LC_6_11_2  (
            .in0(N__35896),
            .in1(N__33669),
            .in2(N__34000),
            .in3(N__24305),
            .lcout(cmd_rdadctmp_12_adj_1536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61896),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_6_11_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_6_11_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i11_LC_6_11_3  (
            .in0(N__33668),
            .in1(N__33973),
            .in2(N__36043),
            .in3(N__35897),
            .lcout(cmd_rdadctmp_11_adj_1537),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61896),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_6_11_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_6_11_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i22_LC_6_11_7  (
            .in0(N__24248),
            .in1(N__33974),
            .in2(N__31275),
            .in3(N__35898),
            .lcout(cmd_rdadctmp_22_adj_1526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61896),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.MOSI_31_LC_6_12_1 .C_ON=1'b0;
    defparam \CLK_DDS.MOSI_31_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.MOSI_31_LC_6_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CLK_DDS.MOSI_31_LC_6_12_1  (
            .in0(N__24273),
            .in1(N__24354),
            .in2(_gnd_net_),
            .in3(N__24618),
            .lcout(DDS_MOSI1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61911),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i14_LC_6_12_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i14_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i14_LC_6_12_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i14_LC_6_12_2  (
            .in0(N__35607),
            .in1(N__35909),
            .in2(N__24258),
            .in3(N__28664),
            .lcout(buf_adcdata_vac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61911),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_6_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_6_12_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i21_LC_6_12_4  (
            .in0(N__33938),
            .in1(N__31268),
            .in2(N__28788),
            .in3(N__35910),
            .lcout(cmd_rdadctmp_21_adj_1527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61911),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_7_i19_3_lut_LC_6_12_6.C_ON=1'b0;
    defparam mux_126_Mux_7_i19_3_lut_LC_6_12_6.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_7_i19_3_lut_LC_6_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_7_i19_3_lut_LC_6_12_6 (
            .in0(N__25045),
            .in1(N__24218),
            .in2(_gnd_net_),
            .in3(N__59475),
            .lcout(),
            .ltout(n19_adj_1714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19345_3_lut_LC_6_12_7.C_ON=1'b0;
    defparam i19345_3_lut_LC_6_12_7.SEQ_MODE=4'b0000;
    defparam i19345_3_lut_LC_6_12_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 i19345_3_lut_LC_6_12_7 (
            .in0(_gnd_net_),
            .in1(N__60665),
            .in2(N__24199),
            .in3(N__24196),
            .lcout(n22272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i10_LC_6_13_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i10_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i10_LC_6_13_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i10_LC_6_13_0  (
            .in0(N__24619),
            .in1(N__24748),
            .in2(N__24373),
            .in3(N__30638),
            .lcout(\CLK_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i11_LC_6_13_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i11_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i11_LC_6_13_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i11_LC_6_13_1  (
            .in0(N__24749),
            .in1(N__24620),
            .in2(N__24415),
            .in3(N__29734),
            .lcout(\CLK_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i12_LC_6_13_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i12_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i12_LC_6_13_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i12_LC_6_13_2  (
            .in0(N__24621),
            .in1(N__24750),
            .in2(N__24406),
            .in3(N__27970),
            .lcout(\CLK_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i13_LC_6_13_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i13_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i13_LC_6_13_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i13_LC_6_13_3  (
            .in0(N__24751),
            .in1(N__24622),
            .in2(N__24397),
            .in3(N__55237),
            .lcout(\CLK_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i14_LC_6_13_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i14_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i14_LC_6_13_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i14_LC_6_13_4  (
            .in0(N__24623),
            .in1(N__24752),
            .in2(N__24388),
            .in3(N__29066),
            .lcout(\CLK_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i15_LC_6_13_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i15_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i15_LC_6_13_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \CLK_DDS.tmp_buf_i15_LC_6_13_5  (
            .in0(N__24753),
            .in1(N__24624),
            .in2(N__25347),
            .in3(N__24379),
            .lcout(tmp_buf_15_adj_1511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i9_LC_6_13_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i9_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i9_LC_6_13_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i9_LC_6_13_6  (
            .in0(N__24626),
            .in1(N__24755),
            .in2(N__24364),
            .in3(N__31891),
            .lcout(\CLK_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i8_LC_6_13_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i8_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i8_LC_6_13_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i8_LC_6_13_7  (
            .in0(N__24754),
            .in1(N__24625),
            .in2(N__24478),
            .in3(N__34150),
            .lcout(\CLK_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61930),
            .ce(N__24465),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i0_LC_6_14_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i0_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i0_LC_6_14_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \CLK_DDS.tmp_buf_i0_LC_6_14_0  (
            .in0(N__24628),
            .in1(N__24756),
            .in2(N__37228),
            .in3(N__24355),
            .lcout(\CLK_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i1_LC_6_14_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i1_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i1_LC_6_14_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i1_LC_6_14_1  (
            .in0(N__24757),
            .in1(N__24629),
            .in2(N__24817),
            .in3(N__42133),
            .lcout(\CLK_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i2_LC_6_14_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i2_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i2_LC_6_14_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i2_LC_6_14_2  (
            .in0(N__24630),
            .in1(N__24758),
            .in2(N__24808),
            .in3(N__42095),
            .lcout(\CLK_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i3_LC_6_14_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i3_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i3_LC_6_14_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i3_LC_6_14_3  (
            .in0(N__24759),
            .in1(N__24631),
            .in2(N__24799),
            .in3(N__36868),
            .lcout(\CLK_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i4_LC_6_14_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i4_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i4_LC_6_14_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i4_LC_6_14_4  (
            .in0(N__24632),
            .in1(N__24760),
            .in2(N__24790),
            .in3(N__49462),
            .lcout(\CLK_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i5_LC_6_14_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i5_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i5_LC_6_14_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \CLK_DDS.tmp_buf_i5_LC_6_14_5  (
            .in0(N__24761),
            .in1(N__28722),
            .in2(N__24781),
            .in3(N__24633),
            .lcout(\CLK_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i6_LC_6_14_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i6_LC_6_14_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i6_LC_6_14_6 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \CLK_DDS.tmp_buf_i6_LC_6_14_6  (
            .in0(N__31327),
            .in1(N__24627),
            .in2(N__24772),
            .in3(N__24762),
            .lcout(\CLK_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i7_LC_6_14_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i7_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i7_LC_6_14_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i7_LC_6_14_7  (
            .in0(N__24763),
            .in1(N__24634),
            .in2(N__24487),
            .in3(N__27908),
            .lcout(\CLK_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61946),
            .ce(N__24469),
            .sr(_gnd_net_));
    defparam buf_dds1_i12_LC_6_15_2.C_ON=1'b0;
    defparam buf_dds1_i12_LC_6_15_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i12_LC_6_15_2.LUT_INIT=16'b1110010000000000;
    LogicCell40 buf_dds1_i12_LC_6_15_2 (
            .in0(N__55388),
            .in1(N__27968),
            .in2(N__44719),
            .in3(N__49518),
            .lcout(buf_dds1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61964),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20439_LC_6_16_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20439_LC_6_16_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20439_LC_6_16_4.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20439_LC_6_16_4 (
            .in0(N__24436),
            .in1(N__60098),
            .in2(N__24430),
            .in3(N__60648),
            .lcout(n23366),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i12899_2_lut_LC_6_16_7 .C_ON=1'b0;
    defparam \ADC_IAC.i12899_2_lut_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i12899_2_lut_LC_6_16_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ADC_IAC.i12899_2_lut_LC_6_16_7  (
            .in0(_gnd_net_),
            .in1(N__25677),
            .in2(_gnd_net_),
            .in3(N__30425),
            .lcout(\ADC_IAC.n15622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_adj_19_LC_6_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_adj_19_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_adj_19_LC_6_17_0 .LUT_INIT=16'b0000000001010010;
    LogicCell40 \ADC_IAC.i1_4_lut_adj_19_LC_6_17_0  (
            .in0(N__30342),
            .in1(N__25818),
            .in2(N__30432),
            .in3(N__39549),
            .lcout(\ADC_IAC.n13667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i2_LC_6_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i2_LC_6_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i2_LC_6_17_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_IAC.adc_state_i2_LC_6_17_1  (
            .in0(N__39551),
            .in1(N__30418),
            .in2(_gnd_net_),
            .in3(N__30345),
            .lcout(DTRIG_N_1182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61993),
            .ce(N__25840),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i1_LC_6_17_2 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i1_LC_6_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i1_LC_6_17_2 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \ADC_IAC.adc_state_i1_LC_6_17_2  (
            .in0(N__30344),
            .in1(_gnd_net_),
            .in2(N__30434),
            .in3(N__39552),
            .lcout(adc_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61993),
            .ce(N__25840),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_61_LC_6_17_3.C_ON=1'b0;
    defparam i1_2_lut_adj_61_LC_6_17_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_61_LC_6_17_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_61_LC_6_17_3 (
            .in0(_gnd_net_),
            .in1(N__30410),
            .in2(_gnd_net_),
            .in3(N__30340),
            .lcout(n21892),
            .ltout(n21892_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_3_lut_LC_6_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.i1_3_lut_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_3_lut_LC_6_17_4 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \ADC_IAC.i1_3_lut_LC_6_17_4  (
            .in0(_gnd_net_),
            .in1(N__25817),
            .in2(N__24853),
            .in3(N__39548),
            .lcout(n13746),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_198_LC_6_17_6.C_ON=1'b0;
    defparam i1_4_lut_adj_198_LC_6_17_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_198_LC_6_17_6.LUT_INIT=16'b0010001100110010;
    LogicCell40 i1_4_lut_adj_198_LC_6_17_6 (
            .in0(N__30343),
            .in1(N__25764),
            .in2(N__30433),
            .in3(N__39550),
            .lcout(n14_adj_1578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_74_LC_6_17_7.C_ON=1'b0;
    defparam i1_2_lut_adj_74_LC_6_17_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_74_LC_6_17_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_74_LC_6_17_7 (
            .in0(_gnd_net_),
            .in1(N__30411),
            .in2(_gnd_net_),
            .in3(N__30341),
            .lcout(n21951),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_2  (
            .in0(N__25719),
            .in1(N__39630),
            .in2(N__24850),
            .in3(N__37748),
            .lcout(cmd_rdadctmp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62001),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_DDS_MCLK1_THRU_LUT4_0_LC_7_1_1.C_ON=1'b0;
    defparam GB_BUFFER_DDS_MCLK1_THRU_LUT4_0_LC_7_1_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_DDS_MCLK1_THRU_LUT4_0_LC_7_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_DDS_MCLK1_THRU_LUT4_0_LC_7_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48421),
            .lcout(GB_BUFFER_DDS_MCLK1_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i8_4_lut_LC_7_2_4 .C_ON=1'b0;
    defparam \ADC_VDC.i8_4_lut_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i8_4_lut_LC_7_2_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \ADC_VDC.i8_4_lut_LC_7_2_4  (
            .in0(N__25950),
            .in1(N__25917),
            .in2(N__26884),
            .in3(N__26904),
            .lcout(\ADC_VDC.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i9_4_lut_LC_7_2_5 .C_ON=1'b0;
    defparam \ADC_VDC.i9_4_lut_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i9_4_lut_LC_7_2_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i9_4_lut_LC_7_2_5  (
            .in0(N__25902),
            .in1(N__25983),
            .in2(N__25969),
            .in3(N__25935),
            .lcout(\ADC_VDC.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12594_12595_reset_LC_7_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12594_12595_reset_LC_7_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i0_12594_12595_reset_LC_7_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.data_tx_i0_12594_12595_reset_LC_7_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64557),
            .lcout(\comm_spi.n15323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53689),
            .ce(),
            .sr(N__35272));
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_18_LC_7_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_18_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_18_LC_7_4_0 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_adj_18_LC_7_4_0  (
            .in0(N__32497),
            .in1(N__33582),
            .in2(N__33432),
            .in3(N__32731),
            .lcout(n13925),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20024_2_lut_LC_7_5_4.C_ON=1'b0;
    defparam i20024_2_lut_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam i20024_2_lut_LC_7_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 i20024_2_lut_LC_7_5_4 (
            .in0(_gnd_net_),
            .in1(N__33380),
            .in2(_gnd_net_),
            .in3(N__32732),
            .lcout(n22388),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_6_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_6_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.SCLK_46_LC_7_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.SCLK_46_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.SCLK_46_LC_7_6_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.SCLK_46_LC_7_6_1  (
            .in0(N__24886),
            .in1(N__24864),
            .in2(N__24895),
            .in3(N__32505),
            .lcout(VDC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42739),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_7_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_7_6_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i12_LC_7_6_2  (
            .in0(N__27054),
            .in1(N__28391),
            .in2(N__27502),
            .in3(N__32723),
            .lcout(cmd_rdadctmp_12_adj_1562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42739),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_7_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_7_6_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i7_LC_7_6_3  (
            .in0(N__32722),
            .in1(N__27129),
            .in2(N__28401),
            .in3(N__27159),
            .lcout(cmd_rdadctmp_7_adj_1567),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42739),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_7_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_7_6_4 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i11_LC_7_6_4  (
            .in0(N__27053),
            .in1(N__27084),
            .in2(N__32733),
            .in3(N__28390),
            .lcout(cmd_rdadctmp_11_adj_1563),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42739),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_7_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_7_6_5 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i2_LC_7_6_5  (
            .in0(N__28386),
            .in1(N__32715),
            .in2(N__27007),
            .in3(N__26970),
            .lcout(cmd_rdadctmp_2_adj_1572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42739),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_7_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_7_6_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i8_LC_7_6_6  (
            .in0(N__27128),
            .in1(N__28421),
            .in2(N__32734),
            .in3(N__28392),
            .lcout(cmd_rdadctmp_8_adj_1566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42739),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_7_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_7_6_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i1_LC_7_6_7  (
            .in0(N__28385),
            .in1(N__32714),
            .in2(N__27006),
            .in3(N__27033),
            .lcout(cmd_rdadctmp_1_adj_1573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42739),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_0  (
            .in0(N__27459),
            .in1(N__27437),
            .in2(N__28394),
            .in3(N__32712),
            .lcout(cmd_rdadctmp_14_adj_1560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42719),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i1_LC_7_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i1_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i1_LC_7_7_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i1_LC_7_7_1  (
            .in0(N__31083),
            .in1(N__33436),
            .in2(N__33627),
            .in3(N__27475),
            .lcout(buf_adcdata_vdc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42719),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_7_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_7_7_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i16_LC_7_7_2  (
            .in0(N__27359),
            .in1(N__27412),
            .in2(N__28395),
            .in3(N__32713),
            .lcout(cmd_rdadctmp_16_adj_1558),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42719),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3  (
            .in0(N__32710),
            .in1(N__28372),
            .in2(N__27601),
            .in3(N__27636),
            .lcout(cmd_rdadctmp_21_adj_1553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42719),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_7_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_7_7_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i10_LC_7_7_4  (
            .in0(N__27083),
            .in1(N__28285),
            .in2(N__28393),
            .in3(N__32711),
            .lcout(cmd_rdadctmp_10_adj_1564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42719),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_7_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_7_7_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i13_LC_7_7_5  (
            .in0(N__32708),
            .in1(N__27458),
            .in2(N__27501),
            .in3(N__28370),
            .lcout(cmd_rdadctmp_13_adj_1561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42719),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i20132_4_lut_4_lut_LC_7_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.i20132_4_lut_4_lut_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i20132_4_lut_4_lut_LC_7_7_6 .LUT_INIT=16'b1111111111100001;
    LogicCell40 \ADC_VDC.i20132_4_lut_4_lut_LC_7_7_6  (
            .in0(N__32506),
            .in1(N__33586),
            .in2(N__33448),
            .in3(N__32707),
            .lcout(n12356),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_7  (
            .in0(N__32709),
            .in1(N__27635),
            .in2(N__27262),
            .in3(N__28371),
            .lcout(cmd_rdadctmp_20_adj_1554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42719),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_7_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_7_8_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i22_LC_7_8_0  (
            .in0(N__32725),
            .in1(N__28380),
            .in2(N__30795),
            .in3(N__27599),
            .lcout(cmd_rdadctmp_22_adj_1552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42757),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i31_3_lut_LC_7_8_2 .C_ON=1'b0;
    defparam \RTD.i31_3_lut_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i31_3_lut_LC_7_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \RTD.i31_3_lut_LC_7_8_2  (
            .in0(N__26846),
            .in1(N__26650),
            .in2(_gnd_net_),
            .in3(N__26235),
            .lcout(\RTD.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_LC_7_8_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_LC_7_8_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \RTD.i1_2_lut_LC_7_8_3  (
            .in0(N__26651),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26847),
            .lcout(\RTD.n79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_7_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_7_8_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i18_LC_7_8_4  (
            .in0(N__32724),
            .in1(N__27294),
            .in2(N__27337),
            .in3(N__28379),
            .lcout(cmd_rdadctmp_18_adj_1556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42757),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_7_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_7_8_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i17_LC_7_8_5  (
            .in0(N__27332),
            .in1(N__27360),
            .in2(N__28396),
            .in3(N__32726),
            .lcout(cmd_rdadctmp_17_adj_1557),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42757),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_7_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_7_8_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i19_LC_7_8_7  (
            .in0(N__27293),
            .in1(N__27260),
            .in2(N__28397),
            .in3(N__32727),
            .lcout(cmd_rdadctmp_19_adj_1555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42757),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i12_LC_7_9_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i12_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i12_LC_7_9_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i12_LC_7_9_0  (
            .in0(N__31074),
            .in1(N__33443),
            .in2(N__30945),
            .in3(N__27553),
            .lcout(buf_adcdata_vdc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i17_LC_7_9_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i17_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i17_LC_7_9_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i17_LC_7_9_1  (
            .in0(N__33440),
            .in1(N__31078),
            .in2(N__48561),
            .in3(N__27718),
            .lcout(buf_adcdata_vdc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i15_LC_7_9_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i15_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i15_LC_7_9_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i15_LC_7_9_2  (
            .in0(N__31076),
            .in1(N__33445),
            .in2(N__25044),
            .in3(N__27520),
            .lcout(buf_adcdata_vdc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i19_LC_7_9_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i19_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i19_LC_7_9_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i19_LC_7_9_3  (
            .in0(N__33441),
            .in1(N__31079),
            .in2(N__27753),
            .in3(N__27688),
            .lcout(buf_adcdata_vdc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i7_LC_7_9_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i7_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i7_LC_7_9_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i7_LC_7_9_4  (
            .in0(N__31077),
            .in1(N__33446),
            .in2(N__25026),
            .in3(N__27277),
            .lcout(buf_adcdata_vdc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i23_LC_7_9_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i23_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i23_LC_7_9_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i23_LC_7_9_5  (
            .in0(N__33442),
            .in1(N__31080),
            .in2(N__25002),
            .in3(N__28474),
            .lcout(buf_adcdata_vdc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i14_LC_7_9_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i14_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i14_LC_7_9_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i14_LC_7_9_6  (
            .in0(N__31075),
            .in1(N__33444),
            .in2(N__28692),
            .in3(N__27535),
            .lcout(buf_adcdata_vdc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i4_LC_7_9_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i4_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i4_LC_7_9_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ADC_VDC.ADC_DATA_i4_LC_7_9_7  (
            .in0(N__27379),
            .in1(N__31081),
            .in2(N__24978),
            .in3(N__33447),
            .lcout(buf_adcdata_vdc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42721),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i10_LC_7_10_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i10_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i10_LC_7_10_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i10_LC_7_10_0  (
            .in0(N__33394),
            .in1(N__31066),
            .in2(N__25104),
            .in3(N__27577),
            .lcout(buf_adcdata_vdc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42748),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i18_LC_7_10_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i18_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i18_LC_7_10_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i18_LC_7_10_2  (
            .in0(N__33395),
            .in1(N__31067),
            .in2(N__31512),
            .in3(N__27703),
            .lcout(buf_adcdata_vdc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42748),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i9_LC_7_10_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i9_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i9_LC_7_10_3 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.ADC_DATA_i9_LC_7_10_3  (
            .in0(N__27619),
            .in1(N__24957),
            .in2(N__31084),
            .in3(N__33402),
            .lcout(buf_adcdata_vdc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42748),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i8_LC_7_10_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i8_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i8_LC_7_10_4 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i8_LC_7_10_4  (
            .in0(N__27238),
            .in1(N__25311),
            .in2(N__33437),
            .in3(N__31072),
            .lcout(buf_adcdata_vdc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42748),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i6_LC_7_10_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i6_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i6_LC_7_10_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i6_LC_7_10_5  (
            .in0(N__31065),
            .in1(N__33398),
            .in2(N__25179),
            .in3(N__27313),
            .lcout(buf_adcdata_vdc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42748),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i22_LC_7_10_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i22_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i22_LC_7_10_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i22_LC_7_10_6  (
            .in0(N__33396),
            .in1(N__31068),
            .in2(N__25158),
            .in3(N__27655),
            .lcout(buf_adcdata_vdc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42748),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i20_LC_7_10_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i20_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i20_LC_7_10_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i20_LC_7_10_7  (
            .in0(N__31064),
            .in1(N__33397),
            .in2(N__25476),
            .in3(N__27673),
            .lcout(buf_adcdata_vdc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42748),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i18_LC_7_11_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i18_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i18_LC_7_11_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i18_LC_7_11_0  (
            .in0(N__35992),
            .in1(N__35597),
            .in2(N__25141),
            .in3(N__31484),
            .lcout(buf_adcdata_vac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61884),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_4_i112_3_lut_LC_7_11_1.C_ON=1'b0;
    defparam mux_125_Mux_4_i112_3_lut_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i112_3_lut_LC_7_11_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_125_Mux_4_i112_3_lut_LC_7_11_1 (
            .in0(N__60543),
            .in1(N__34098),
            .in2(_gnd_net_),
            .in3(N__31405),
            .lcout(),
            .ltout(n112_adj_1786_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_4_i127_3_lut_LC_7_11_2.C_ON=1'b0;
    defparam mux_125_Mux_4_i127_3_lut_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i127_3_lut_LC_7_11_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 mux_125_Mux_4_i127_3_lut_LC_7_11_2 (
            .in0(_gnd_net_),
            .in1(N__61412),
            .in2(N__25108),
            .in3(N__27802),
            .lcout(comm_buf_0_7_N_543_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i11_LC_7_11_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i11_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i11_LC_7_11_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i11_LC_7_11_3  (
            .in0(N__35596),
            .in1(N__35993),
            .in2(N__28821),
            .in3(N__41208),
            .lcout(buf_adcdata_vac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61884),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_2_i19_3_lut_LC_7_11_5.C_ON=1'b0;
    defparam mux_126_Mux_2_i19_3_lut_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_2_i19_3_lut_LC_7_11_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_2_i19_3_lut_LC_7_11_5 (
            .in0(N__25105),
            .in1(N__25076),
            .in2(_gnd_net_),
            .in3(N__59335),
            .lcout(n19_adj_1747),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_6_i111_3_lut_LC_7_11_6.C_ON=1'b0;
    defparam mux_125_Mux_6_i111_3_lut_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_6_i111_3_lut_LC_7_11_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_125_Mux_6_i111_3_lut_LC_7_11_6 (
            .in0(N__59336),
            .in1(N__25356),
            .in2(_gnd_net_),
            .in3(N__34321),
            .lcout(n111_adj_1771),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i22_LC_7_11_7.C_ON=1'b0;
    defparam comm_test_buf_24_i22_LC_7_11_7.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i22_LC_7_11_7.LUT_INIT=16'b0000110010101010;
    LogicCell40 comm_test_buf_24_i22_LC_7_11_7 (
            .in0(N__25357),
            .in1(N__40526),
            .in2(N__57869),
            .in3(N__45422),
            .lcout(comm_test_buf_24_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61884),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i12_LC_7_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i12_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i12_LC_7_12_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i12_LC_7_12_0  (
            .in0(N__35608),
            .in1(N__36013),
            .in2(N__28789),
            .in3(N__30911),
            .lcout(buf_adcdata_vac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61897),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i15_LC_7_12_1.C_ON=1'b0;
    defparam buf_dds1_i15_LC_7_12_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i15_LC_7_12_1.LUT_INIT=16'b1010000010001000;
    LogicCell40 buf_dds1_i15_LC_7_12_1 (
            .in0(N__49561),
            .in1(N__25340),
            .in2(N__46662),
            .in3(N__55432),
            .lcout(buf_dds1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61897),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_6_i112_3_lut_LC_7_12_2.C_ON=1'b0;
    defparam mux_125_Mux_6_i112_3_lut_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_6_i112_3_lut_LC_7_12_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_125_Mux_6_i112_3_lut_LC_7_12_2 (
            .in0(N__34299),
            .in1(N__60615),
            .in2(_gnd_net_),
            .in3(N__25321),
            .lcout(n112_adj_1772),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i3_LC_7_12_3.C_ON=1'b0;
    defparam buf_cfgRTD_i3_LC_7_12_3.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i3_LC_7_12_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i3_LC_7_12_3 (
            .in0(N__56850),
            .in1(N__48814),
            .in2(_gnd_net_),
            .in3(N__25197),
            .lcout(buf_cfgRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61897),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i14_LC_7_12_4.C_ON=1'b0;
    defparam buf_dds1_i14_LC_7_12_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i14_LC_7_12_4.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i14_LC_7_12_4 (
            .in0(N__29067),
            .in1(N__55371),
            .in2(N__40570),
            .in3(N__49560),
            .lcout(buf_dds1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61897),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_0_i19_3_lut_LC_7_12_5.C_ON=1'b0;
    defparam mux_126_Mux_0_i19_3_lut_LC_7_12_5.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_0_i19_3_lut_LC_7_12_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_0_i19_3_lut_LC_7_12_5 (
            .in0(N__25315),
            .in1(N__25290),
            .in2(_gnd_net_),
            .in3(N__59467),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_6_i127_3_lut_LC_7_12_6.C_ON=1'b0;
    defparam mux_127_Mux_6_i127_3_lut_LC_7_12_6.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_6_i127_3_lut_LC_7_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_6_i127_3_lut_LC_7_12_6 (
            .in0(N__34300),
            .in1(N__25261),
            .in2(_gnd_net_),
            .in3(N__61394),
            .lcout(comm_buf_2_7_N_575_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i20_3_lut_LC_7_12_7.C_ON=1'b0;
    defparam mux_125_Mux_3_i20_3_lut_LC_7_12_7.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i20_3_lut_LC_7_12_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_3_i20_3_lut_LC_7_12_7 (
            .in0(N__25249),
            .in1(N__25196),
            .in2(_gnd_net_),
            .in3(N__59468),
            .lcout(n20_adj_1790),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20543_LC_7_13_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20543_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20543_LC_7_13_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20543_LC_7_13_0 (
            .in0(N__27736),
            .in1(N__60080),
            .in2(N__25489),
            .in3(N__60611),
            .lcout(),
            .ltout(n23498_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23498_bdd_4_lut_LC_7_13_1.C_ON=1'b0;
    defparam n23498_bdd_4_lut_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam n23498_bdd_4_lut_LC_7_13_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n23498_bdd_4_lut_LC_7_13_1 (
            .in0(N__60081),
            .in1(N__25423),
            .in2(N__25480),
            .in3(N__25417),
            .lcout(n23501),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_4_i19_3_lut_LC_7_13_4.C_ON=1'b0;
    defparam mux_125_Mux_4_i19_3_lut_LC_7_13_4.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i19_3_lut_LC_7_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_125_Mux_4_i19_3_lut_LC_7_13_4 (
            .in0(N__59490),
            .in1(N__25477),
            .in2(_gnd_net_),
            .in3(N__25445),
            .lcout(n19_adj_1780),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i16_3_lut_LC_7_13_6.C_ON=1'b0;
    defparam mux_125_Mux_3_i16_3_lut_LC_7_13_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i16_3_lut_LC_7_13_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_125_Mux_3_i16_3_lut_LC_7_13_6 (
            .in0(N__59488),
            .in1(N__29733),
            .in2(_gnd_net_),
            .in3(N__32903),
            .lcout(n16_adj_1787),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i17_3_lut_LC_7_13_7.C_ON=1'b0;
    defparam mux_125_Mux_3_i17_3_lut_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i17_3_lut_LC_7_13_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_3_i17_3_lut_LC_7_13_7 (
            .in0(N__27993),
            .in1(N__29799),
            .in2(_gnd_net_),
            .in3(N__59489),
            .lcout(n17_adj_1788),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_LC_7_14_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_LC_7_14_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_LC_7_14_0.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_LC_7_14_0 (
            .in0(N__59491),
            .in1(N__31602),
            .in2(N__25392),
            .in3(N__60610),
            .lcout(n23540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i10_LC_7_14_1.C_ON=1'b0;
    defparam buf_dds1_i10_LC_7_14_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i10_LC_7_14_1.LUT_INIT=16'b1010000010001000;
    LogicCell40 buf_dds1_i10_LC_7_14_1 (
            .in0(N__49567),
            .in1(N__30639),
            .in2(N__40947),
            .in3(N__55369),
            .lcout(buf_dds1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61931),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i23_LC_7_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i23_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i23_LC_7_14_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i23_LC_7_14_3  (
            .in0(N__39351),
            .in1(N__39651),
            .in2(N__25372),
            .in3(N__25388),
            .lcout(buf_adcdata_iac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61931),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i7_LC_7_14_4.C_ON=1'b0;
    defparam buf_dds1_i7_LC_7_14_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i7_LC_7_14_4.LUT_INIT=16'b1110010000000000;
    LogicCell40 buf_dds1_i7_LC_7_14_4 (
            .in0(N__55368),
            .in1(N__27909),
            .in2(N__55849),
            .in3(N__49569),
            .lcout(buf_dds1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61931),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_7_14_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_7_14_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i31_LC_7_14_5  (
            .in0(N__31797),
            .in1(N__39652),
            .in2(N__25371),
            .in3(N__37772),
            .lcout(cmd_rdadctmp_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61931),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20377_LC_7_14_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20377_LC_7_14_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20377_LC_7_14_6.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20377_LC_7_14_6 (
            .in0(N__25543),
            .in1(N__60076),
            .in2(N__25534),
            .in3(N__60609),
            .lcout(n23300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i2_LC_7_14_7.C_ON=1'b0;
    defparam buf_dds1_i2_LC_7_14_7.SEQ_MODE=4'b1000;
    defparam buf_dds1_i2_LC_7_14_7.LUT_INIT=16'b1010000010001000;
    LogicCell40 buf_dds1_i2_LC_7_14_7 (
            .in0(N__49568),
            .in1(N__42096),
            .in2(N__52935),
            .in3(N__55370),
            .lcout(buf_dds1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61931),
            .ce(),
            .sr(_gnd_net_));
    defparam i19116_4_lut_LC_7_15_3.C_ON=1'b0;
    defparam i19116_4_lut_LC_7_15_3.SEQ_MODE=4'b0000;
    defparam i19116_4_lut_LC_7_15_3.LUT_INIT=16'b1111111111100100;
    LogicCell40 i19116_4_lut_LC_7_15_3 (
            .in0(N__45809),
            .in1(N__34700),
            .in2(N__34798),
            .in3(N__39170),
            .lcout(),
            .ltout(n22041_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_trig_303_LC_7_15_4.C_ON=1'b0;
    defparam acadc_trig_303_LC_7_15_4.SEQ_MODE=4'b1000;
    defparam acadc_trig_303_LC_7_15_4.LUT_INIT=16'b1111010000000100;
    LogicCell40 acadc_trig_303_LC_7_15_4 (
            .in0(N__34701),
            .in1(N__45810),
            .in2(N__25507),
            .in3(N__25867),
            .lcout(acadc_trig),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_trig_303C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.bit_cnt_i0_LC_7_16_0 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i0_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i0_LC_7_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i0_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__25585),
            .in2(_gnd_net_),
            .in3(N__25504),
            .lcout(\ADC_IAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\ADC_IAC.n20676 ),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.bit_cnt_i1_LC_7_16_1 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i1_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i1_LC_7_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i1_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__25623),
            .in2(_gnd_net_),
            .in3(N__25501),
            .lcout(\ADC_IAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_IAC.n20676 ),
            .carryout(\ADC_IAC.n20677 ),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.bit_cnt_i2_LC_7_16_2 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i2_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i2_LC_7_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i2_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__25609),
            .in2(_gnd_net_),
            .in3(N__25498),
            .lcout(\ADC_IAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_IAC.n20677 ),
            .carryout(\ADC_IAC.n20678 ),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.bit_cnt_i3_LC_7_16_3 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i3_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i3_LC_7_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i3_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__25636),
            .in2(_gnd_net_),
            .in3(N__25495),
            .lcout(\ADC_IAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_IAC.n20678 ),
            .carryout(\ADC_IAC.n20679 ),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.bit_cnt_i4_LC_7_16_4 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i4_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i4_LC_7_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i4_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__25648),
            .in2(_gnd_net_),
            .in3(N__25492),
            .lcout(\ADC_IAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_IAC.n20679 ),
            .carryout(\ADC_IAC.n20680 ),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.bit_cnt_i5_LC_7_16_5 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i5_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i5_LC_7_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i5_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__25558),
            .in2(_gnd_net_),
            .in3(N__25696),
            .lcout(\ADC_IAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_IAC.n20680 ),
            .carryout(\ADC_IAC.n20681 ),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.bit_cnt_i6_LC_7_16_6 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i6_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i6_LC_7_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i6_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__25597),
            .in2(_gnd_net_),
            .in3(N__25693),
            .lcout(\ADC_IAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_IAC.n20681 ),
            .carryout(\ADC_IAC.n20682 ),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.bit_cnt_i7_LC_7_16_7 .C_ON=1'b0;
    defparam \ADC_IAC.bit_cnt_i7_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i7_LC_7_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i7_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__25570),
            .in2(_gnd_net_),
            .in3(N__25690),
            .lcout(\ADC_IAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61965),
            .ce(N__25687),
            .sr(N__25666));
    defparam \ADC_IAC.i1_2_lut_LC_7_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.i1_2_lut_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_2_lut_LC_7_17_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \ADC_IAC.i1_2_lut_LC_7_17_0  (
            .in0(N__30365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25654),
            .lcout(\ADC_IAC.n22032 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_LC_7_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_LC_7_17_1 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_IAC.i1_4_lut_LC_7_17_1  (
            .in0(N__30422),
            .in1(N__39553),
            .in2(N__25819),
            .in3(N__25868),
            .lcout(\ADC_IAC.n22031 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19186_4_lut_LC_7_17_2 .C_ON=1'b0;
    defparam \ADC_IAC.i19186_4_lut_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19186_4_lut_LC_7_17_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_IAC.i19186_4_lut_LC_7_17_2  (
            .in0(N__25647),
            .in1(N__25635),
            .in2(N__25624),
            .in3(N__25608),
            .lcout(),
            .ltout(\ADC_IAC.n22113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19201_4_lut_LC_7_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.i19201_4_lut_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19201_4_lut_LC_7_17_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_IAC.i19201_4_lut_LC_7_17_3  (
            .in0(N__25596),
            .in1(N__25584),
            .in2(N__25573),
            .in3(N__25569),
            .lcout(),
            .ltout(\ADC_IAC.n22128_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19757_4_lut_LC_7_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.i19757_4_lut_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19757_4_lut_LC_7_17_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_IAC.i19757_4_lut_LC_7_17_4  (
            .in0(N__39555),
            .in1(N__25557),
            .in2(N__25546),
            .in3(N__30367),
            .lcout(),
            .ltout(\ADC_IAC.n22384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i0_LC_7_17_5 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i0_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i0_LC_7_17_5 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \ADC_IAC.adc_state_i0_LC_7_17_5  (
            .in0(N__30424),
            .in1(N__30366),
            .in2(N__25888),
            .in3(N__39556),
            .lcout(adc_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61980),
            .ce(N__25885),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i30_4_lut_LC_7_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.i30_4_lut_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i30_4_lut_LC_7_17_6 .LUT_INIT=16'b1011000110000001;
    LogicCell40 \ADC_IAC.i30_4_lut_LC_7_17_6  (
            .in0(N__25869),
            .in1(N__30423),
            .in2(N__30372),
            .in3(N__25816),
            .lcout(),
            .ltout(\ADC_IAC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i20195_2_lut_LC_7_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.i20195_2_lut_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i20195_2_lut_LC_7_17_7 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \ADC_IAC.i20195_2_lut_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25843),
            .in3(N__39554),
            .lcout(\ADC_IAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.CS_37_LC_7_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.CS_37_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.CS_37_LC_7_18_0 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \ADC_IAC.CS_37_LC_7_18_0  (
            .in0(N__25831),
            .in1(N__25825),
            .in2(N__39715),
            .in3(N__25812),
            .lcout(IAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61994),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_7_18_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_7_18_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i2_LC_7_18_2  (
            .in0(N__25752),
            .in1(N__39622),
            .in2(N__25708),
            .in3(N__37746),
            .lcout(cmd_rdadctmp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61994),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_3  (
            .in0(N__37743),
            .in1(N__25743),
            .in2(N__39713),
            .in3(N__25753),
            .lcout(cmd_rdadctmp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61994),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_4  (
            .in0(N__25744),
            .in1(N__39623),
            .in2(N__25735),
            .in3(N__37747),
            .lcout(cmd_rdadctmp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61994),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_5  (
            .in0(N__37744),
            .in1(N__30480),
            .in2(N__39714),
            .in3(N__25734),
            .lcout(cmd_rdadctmp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61994),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_7_18_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_7_18_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i1_LC_7_18_6  (
            .in0(N__25704),
            .in1(N__39621),
            .in2(N__25723),
            .in3(N__37745),
            .lcout(cmd_rdadctmp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61994),
            .ce(),
            .sr(_gnd_net_));
    defparam EIS_SYNCCLK_I_0_1_lut_LC_8_1_2.C_ON=1'b0;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_8_1_2.SEQ_MODE=4'b0000;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_8_1_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 EIS_SYNCCLK_I_0_1_lut_LC_8_1_2 (
            .in0(N__26038),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(IAC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.avg_cnt_i0_LC_8_2_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i0_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i0_LC_8_2_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i0_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__28045),
            .in2(_gnd_net_),
            .in3(N__25987),
            .lcout(\ADC_VDC.avg_cnt_0 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\ADC_VDC.n20725 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i1_LC_8_2_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i1_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i1_LC_8_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i1_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__25984),
            .in2(_gnd_net_),
            .in3(N__25972),
            .lcout(\ADC_VDC.avg_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n20725 ),
            .carryout(\ADC_VDC.n20726 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i2_LC_8_2_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i2_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i2_LC_8_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i2_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__25968),
            .in2(_gnd_net_),
            .in3(N__25954),
            .lcout(\ADC_VDC.avg_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n20726 ),
            .carryout(\ADC_VDC.n20727 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i3_LC_8_2_3 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i3_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i3_LC_8_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i3_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__25951),
            .in2(_gnd_net_),
            .in3(N__25939),
            .lcout(\ADC_VDC.avg_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n20727 ),
            .carryout(\ADC_VDC.n20728 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i4_LC_8_2_4 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i4_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i4_LC_8_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i4_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(N__25936),
            .in2(_gnd_net_),
            .in3(N__25924),
            .lcout(\ADC_VDC.avg_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n20728 ),
            .carryout(\ADC_VDC.n20729 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i5_LC_8_2_5 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i5_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i5_LC_8_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i5_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__28033),
            .in2(_gnd_net_),
            .in3(N__25921),
            .lcout(\ADC_VDC.avg_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n20729 ),
            .carryout(\ADC_VDC.n20730 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i6_LC_8_2_6 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i6_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i6_LC_8_2_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i6_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(N__25918),
            .in2(_gnd_net_),
            .in3(N__25906),
            .lcout(\ADC_VDC.avg_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n20730 ),
            .carryout(\ADC_VDC.n20731 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i7_LC_8_2_7 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i7_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i7_LC_8_2_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i7_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__25903),
            .in2(_gnd_net_),
            .in3(N__25891),
            .lcout(\ADC_VDC.avg_cnt_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n20731 ),
            .carryout(\ADC_VDC.n20732 ),
            .clk(N__42747),
            .ce(N__28637),
            .sr(N__28563));
    defparam \ADC_VDC.avg_cnt_i8_LC_8_3_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i8_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i8_LC_8_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i8_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__28017),
            .in2(_gnd_net_),
            .in3(N__26908),
            .lcout(\ADC_VDC.avg_cnt_8 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\ADC_VDC.n20733 ),
            .clk(N__42737),
            .ce(N__28636),
            .sr(N__28562));
    defparam \ADC_VDC.avg_cnt_i9_LC_8_3_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i9_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i9_LC_8_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i9_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__26905),
            .in2(_gnd_net_),
            .in3(N__26893),
            .lcout(\ADC_VDC.avg_cnt_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n20733 ),
            .carryout(\ADC_VDC.n20734 ),
            .clk(N__42737),
            .ce(N__28636),
            .sr(N__28562));
    defparam \ADC_VDC.avg_cnt_i10_LC_8_3_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i10_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i10_LC_8_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i10_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__28180),
            .in2(_gnd_net_),
            .in3(N__26890),
            .lcout(\ADC_VDC.avg_cnt_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n20734 ),
            .carryout(\ADC_VDC.n20735 ),
            .clk(N__42737),
            .ce(N__28636),
            .sr(N__28562));
    defparam \ADC_VDC.avg_cnt_i11_LC_8_3_3 .C_ON=1'b0;
    defparam \ADC_VDC.avg_cnt_i11_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i11_LC_8_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i11_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__26880),
            .in2(_gnd_net_),
            .in3(N__26887),
            .lcout(\ADC_VDC.avg_cnt_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42737),
            .ce(N__28636),
            .sr(N__28562));
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_8_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_8_4_3 .LUT_INIT=16'b1111011111110010;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_LC_8_4_3  (
            .in0(N__32607),
            .in1(N__28123),
            .in2(N__33381),
            .in3(N__30673),
            .lcout(\ADC_VDC.n13865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_27_LC_8_4_5 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_27_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_27_LC_8_4_5 .LUT_INIT=16'b1011000010000110;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_27_LC_8_4_5  (
            .in0(N__26822),
            .in1(N__26652),
            .in2(N__26472),
            .in3(N__26213),
            .lcout(\RTD.n18275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19145_2_lut_3_lut_LC_8_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.i19145_2_lut_3_lut_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19145_2_lut_3_lut_LC_8_4_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ADC_VDC.i19145_2_lut_3_lut_LC_8_4_6  (
            .in0(N__32828),
            .in1(N__32486),
            .in2(_gnd_net_),
            .in3(N__33516),
            .lcout(\ADC_VDC.n22071 ),
            .ltout(\ADC_VDC.n22071_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i34_3_lut_4_lut_LC_8_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i34_3_lut_4_lut_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i34_3_lut_4_lut_LC_8_4_7 .LUT_INIT=16'b0001101100001010;
    LogicCell40 \ADC_VDC.i34_3_lut_4_lut_LC_8_4_7  (
            .in0(N__32606),
            .in1(N__33552),
            .in2(N__26041),
            .in3(N__32829),
            .lcout(\ADC_VDC.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_8_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_8_5_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i4_LC_8_5_0  (
            .in0(N__32619),
            .in1(N__27218),
            .in2(N__26941),
            .in3(N__28344),
            .lcout(cmd_rdadctmp_4_adj_1570),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42663),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_1  (
            .in0(N__27219),
            .in1(N__27188),
            .in2(N__28381),
            .in3(N__32622),
            .lcout(cmd_rdadctmp_5_adj_1569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42663),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_2  (
            .in0(N__32617),
            .in1(N__27439),
            .in2(N__27410),
            .in3(N__28342),
            .lcout(cmd_rdadctmp_15_adj_1559),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42663),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4  (
            .in0(N__32620),
            .in1(N__28338),
            .in2(N__27193),
            .in3(N__27158),
            .lcout(cmd_rdadctmp_6_adj_1568),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42663),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5  (
            .in0(N__28337),
            .in1(N__27032),
            .in2(N__32800),
            .in3(N__32621),
            .lcout(cmd_rdadctmp_0_adj_1574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42663),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_6  (
            .in0(N__32618),
            .in1(N__26969),
            .in2(N__26940),
            .in3(N__28343),
            .lcout(cmd_rdadctmp_3_adj_1571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42663),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__27013),
            .in2(N__27034),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.cmd_rdadcbuf_0 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\ADC_VDC.n20690 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__26983),
            .in2(N__27005),
            .in3(N__26977),
            .lcout(\ADC_VDC.cmd_rdadcbuf_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n20690 ),
            .carryout(\ADC_VDC.n20691 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__26950),
            .in2(N__26974),
            .in3(N__26944),
            .lcout(\ADC_VDC.cmd_rdadcbuf_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n20691 ),
            .carryout(\ADC_VDC.n20692 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__26917),
            .in2(N__26939),
            .in3(N__26911),
            .lcout(\ADC_VDC.cmd_rdadcbuf_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n20692 ),
            .carryout(\ADC_VDC.n20693 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__27202),
            .in2(N__27220),
            .in3(N__27196),
            .lcout(\ADC_VDC.cmd_rdadcbuf_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n20693 ),
            .carryout(\ADC_VDC.n20694 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__27172),
            .in2(N__27192),
            .in3(N__27163),
            .lcout(\ADC_VDC.cmd_rdadcbuf_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n20694 ),
            .carryout(\ADC_VDC.n20695 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__27139),
            .in2(N__27160),
            .in3(N__27133),
            .lcout(\ADC_VDC.cmd_rdadcbuf_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n20695 ),
            .carryout(\ADC_VDC.n20696 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__27112),
            .in2(N__27130),
            .in3(N__27106),
            .lcout(\ADC_VDC.cmd_rdadcbuf_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n20696 ),
            .carryout(\ADC_VDC.n20697 ),
            .clk(N__42738),
            .ce(N__28626),
            .sr(N__28557));
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__27103),
            .in2(N__28425),
            .in3(N__27097),
            .lcout(\ADC_VDC.cmd_rdadcbuf_8 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\ADC_VDC.n20698 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__27094),
            .in2(N__28281),
            .in3(N__27088),
            .lcout(\ADC_VDC.cmd_rdadcbuf_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n20698 ),
            .carryout(\ADC_VDC.n20699 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__27064),
            .in2(N__27085),
            .in3(N__27058),
            .lcout(\ADC_VDC.cmd_rdadcbuf_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n20699 ),
            .carryout(\ADC_VDC.n20700 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__30957),
            .in2(N__27055),
            .in3(N__27037),
            .lcout(cmd_rdadcbuf_11),
            .ltout(),
            .carryin(\ADC_VDC.n20700 ),
            .carryout(\ADC_VDC.n20701 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__27474),
            .in2(N__27500),
            .in3(N__27463),
            .lcout(cmd_rdadcbuf_12),
            .ltout(),
            .carryin(\ADC_VDC.n20701 ),
            .carryout(\ADC_VDC.n20702 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__28242),
            .in2(N__27460),
            .in3(N__27442),
            .lcout(cmd_rdadcbuf_13),
            .ltout(),
            .carryin(\ADC_VDC.n20702 ),
            .carryout(\ADC_VDC.n20703 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__28437),
            .in2(N__27438),
            .in3(N__27415),
            .lcout(cmd_rdadcbuf_14),
            .ltout(),
            .carryin(\ADC_VDC.n20703 ),
            .carryout(\ADC_VDC.n20704 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__27375),
            .in2(N__27411),
            .in3(N__27364),
            .lcout(cmd_rdadcbuf_15),
            .ltout(),
            .carryin(\ADC_VDC.n20704 ),
            .carryout(\ADC_VDC.n20705 ),
            .clk(N__42718),
            .ce(N__28625),
            .sr(N__28553));
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__28227),
            .in2(N__27361),
            .in3(N__27340),
            .lcout(cmd_rdadcbuf_16),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\ADC_VDC.n20706 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__27309),
            .in2(N__27336),
            .in3(N__27298),
            .lcout(cmd_rdadcbuf_17),
            .ltout(),
            .carryin(\ADC_VDC.n20706 ),
            .carryout(\ADC_VDC.n20707 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__27276),
            .in2(N__27295),
            .in3(N__27265),
            .lcout(cmd_rdadcbuf_18),
            .ltout(),
            .carryin(\ADC_VDC.n20707 ),
            .carryout(\ADC_VDC.n20708 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__27234),
            .in2(N__27261),
            .in3(N__27223),
            .lcout(cmd_rdadcbuf_19),
            .ltout(),
            .carryin(\ADC_VDC.n20708 ),
            .carryout(\ADC_VDC.n20709 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__27615),
            .in2(N__27637),
            .in3(N__27604),
            .lcout(cmd_rdadcbuf_20),
            .ltout(),
            .carryin(\ADC_VDC.n20709 ),
            .carryout(\ADC_VDC.n20710 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__27576),
            .in2(N__27600),
            .in3(N__27559),
            .lcout(cmd_rdadcbuf_21),
            .ltout(),
            .carryin(\ADC_VDC.n20710 ),
            .carryout(\ADC_VDC.n20711 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__28254),
            .in2(N__30794),
            .in3(N__27556),
            .lcout(cmd_rdadcbuf_22),
            .ltout(),
            .carryin(\ADC_VDC.n20711 ),
            .carryout(\ADC_VDC.n20712 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__27552),
            .in2(N__30760),
            .in3(N__27541),
            .lcout(cmd_rdadcbuf_23),
            .ltout(),
            .carryin(\ADC_VDC.n20712 ),
            .carryout(\ADC_VDC.n20713 ),
            .clk(N__42740),
            .ce(N__28638),
            .sr(N__28549));
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__31095),
            .in2(_gnd_net_),
            .in3(N__27538),
            .lcout(cmd_rdadcbuf_24),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\ADC_VDC.n20714 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__27534),
            .in2(_gnd_net_),
            .in3(N__27523),
            .lcout(cmd_rdadcbuf_25),
            .ltout(),
            .carryin(\ADC_VDC.n20714 ),
            .carryout(\ADC_VDC.n20715 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__27519),
            .in2(_gnd_net_),
            .in3(N__27508),
            .lcout(cmd_rdadcbuf_26),
            .ltout(),
            .carryin(\ADC_VDC.n20715 ),
            .carryout(\ADC_VDC.n20716 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__28191),
            .in2(_gnd_net_),
            .in3(N__27505),
            .lcout(cmd_rdadcbuf_27),
            .ltout(),
            .carryin(\ADC_VDC.n20716 ),
            .carryout(\ADC_VDC.n20717 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__27717),
            .in2(_gnd_net_),
            .in3(N__27706),
            .lcout(cmd_rdadcbuf_28),
            .ltout(),
            .carryin(\ADC_VDC.n20717 ),
            .carryout(\ADC_VDC.n20718 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__27702),
            .in2(_gnd_net_),
            .in3(N__27691),
            .lcout(cmd_rdadcbuf_29),
            .ltout(),
            .carryin(\ADC_VDC.n20718 ),
            .carryout(\ADC_VDC.n20719 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__27687),
            .in2(_gnd_net_),
            .in3(N__27676),
            .lcout(cmd_rdadcbuf_30),
            .ltout(),
            .carryin(\ADC_VDC.n20719 ),
            .carryout(\ADC_VDC.n20720 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__27672),
            .in2(_gnd_net_),
            .in3(N__27661),
            .lcout(cmd_rdadcbuf_31),
            .ltout(),
            .carryin(\ADC_VDC.n20720 ),
            .carryout(\ADC_VDC.n20721 ),
            .clk(N__42720),
            .ce(N__28621),
            .sr(N__28561));
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__31125),
            .in2(_gnd_net_),
            .in3(N__27658),
            .lcout(cmd_rdadcbuf_32),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\ADC_VDC.n20722 ),
            .clk(N__42758),
            .ce(N__28642),
            .sr(N__28564));
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__27654),
            .in2(_gnd_net_),
            .in3(N__27643),
            .lcout(cmd_rdadcbuf_33),
            .ltout(),
            .carryin(\ADC_VDC.n20722 ),
            .carryout(\ADC_VDC.n20723 ),
            .clk(N__42758),
            .ce(N__28642),
            .sr(N__28564));
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .C_ON=1'b0;
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.add_23_36_lut_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__28466),
            .in2(_gnd_net_),
            .in3(N__27640),
            .lcout(\ADC_VDC.cmd_rdadcbuf_35_N_1344_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_12640_12641_reset_LC_8_11_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12640_12641_reset_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i6_12640_12641_reset_LC_8_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.data_tx_i6_12640_12641_reset_LC_8_11_0  (
            .in0(N__36615),
            .in1(N__36591),
            .in2(_gnd_net_),
            .in3(N__36564),
            .lcout(\comm_spi.n15369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53665),
            .ce(),
            .sr(N__34114));
    defparam comm_cmd_1__bdd_4_lut_20533_LC_8_12_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20533_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20533_LC_8_12_0.LUT_INIT=16'b1110101001001010;
    LogicCell40 comm_cmd_1__bdd_4_lut_20533_LC_8_12_0 (
            .in0(N__60642),
            .in1(N__49705),
            .in2(N__60091),
            .in3(N__53026),
            .lcout(),
            .ltout(n23474_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23474_bdd_4_lut_LC_8_12_1.C_ON=1'b0;
    defparam n23474_bdd_4_lut_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam n23474_bdd_4_lut_LC_8_12_1.LUT_INIT=16'b1111000011001010;
    LogicCell40 n23474_bdd_4_lut_LC_8_12_1 (
            .in0(N__39835),
            .in1(N__27763),
            .in2(N__27808),
            .in3(N__60052),
            .lcout(),
            .ltout(n23477_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1662065_i1_3_lut_LC_8_12_2.C_ON=1'b0;
    defparam i1662065_i1_3_lut_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam i1662065_i1_3_lut_LC_8_12_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1662065_i1_3_lut_LC_8_12_2 (
            .in0(_gnd_net_),
            .in1(N__27724),
            .in2(N__27805),
            .in3(N__61053),
            .lcout(n30_adj_1784),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1662668_i1_3_lut_LC_8_12_3.C_ON=1'b0;
    defparam i1662668_i1_3_lut_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam i1662668_i1_3_lut_LC_8_12_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 i1662668_i1_3_lut_LC_8_12_3 (
            .in0(N__61054),
            .in1(N__29032),
            .in2(_gnd_net_),
            .in3(N__28756),
            .lcout(),
            .ltout(n30_adj_1768_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_6_i127_3_lut_LC_8_12_4.C_ON=1'b0;
    defparam mux_125_Mux_6_i127_3_lut_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_6_i127_3_lut_LC_8_12_4.LUT_INIT=16'b1101100011011000;
    LogicCell40 mux_125_Mux_6_i127_3_lut_LC_8_12_4 (
            .in0(N__61390),
            .in1(N__27796),
            .in2(N__27787),
            .in3(_gnd_net_),
            .lcout(comm_buf_0_7_N_543_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20483_LC_8_12_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20483_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20483_LC_8_12_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20483_LC_8_12_5 (
            .in0(N__27784),
            .in1(N__60048),
            .in2(N__28834),
            .in3(N__60641),
            .lcout(n23426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_4_i127_3_lut_LC_8_12_6.C_ON=1'b0;
    defparam mux_127_Mux_4_i127_3_lut_LC_8_12_6.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_4_i127_3_lut_LC_8_12_6.LUT_INIT=16'b1010110010101100;
    LogicCell40 mux_127_Mux_4_i127_3_lut_LC_8_12_6 (
            .in0(N__34102),
            .in1(N__27778),
            .in2(N__61413),
            .in3(_gnd_net_),
            .lcout(comm_buf_2_7_N_575_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20034_2_lut_LC_8_12_7.C_ON=1'b0;
    defparam i20034_2_lut_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam i20034_2_lut_LC_8_12_7.LUT_INIT=16'b0011001100000000;
    LogicCell40 i20034_2_lut_LC_8_12_7 (
            .in0(_gnd_net_),
            .in1(N__59350),
            .in2(_gnd_net_),
            .in3(N__38698),
            .lcout(n22358),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i19_3_lut_LC_8_13_0.C_ON=1'b0;
    defparam mux_125_Mux_3_i19_3_lut_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i19_3_lut_LC_8_13_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_125_Mux_3_i19_3_lut_LC_8_13_0 (
            .in0(N__27824),
            .in1(N__27757),
            .in2(_gnd_net_),
            .in3(N__59483),
            .lcout(n19_adj_1789),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23426_bdd_4_lut_LC_8_13_1.C_ON=1'b0;
    defparam n23426_bdd_4_lut_LC_8_13_1.SEQ_MODE=4'b0000;
    defparam n23426_bdd_4_lut_LC_8_13_1.LUT_INIT=16'b1010101011011000;
    LogicCell40 n23426_bdd_4_lut_LC_8_13_1 (
            .in0(N__27730),
            .in1(N__36814),
            .in2(N__27946),
            .in3(N__60094),
            .lcout(n23429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_337_LC_8_13_3.C_ON=1'b0;
    defparam i1_4_lut_adj_337_LC_8_13_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_337_LC_8_13_3.LUT_INIT=16'b1110010000000000;
    LogicCell40 i1_4_lut_adj_337_LC_8_13_3 (
            .in0(N__59484),
            .in1(N__52927),
            .in2(N__40978),
            .in3(N__37403),
            .lcout(n11983),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i9_LC_8_13_4.C_ON=1'b0;
    defparam buf_dds1_i9_LC_8_13_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i9_LC_8_13_4.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i9_LC_8_13_4 (
            .in0(N__31877),
            .in1(N__55431),
            .in2(N__44646),
            .in3(N__49562),
            .lcout(buf_dds1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61898),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i11_LC_8_13_6.C_ON=1'b0;
    defparam buf_dds0_i11_LC_8_13_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i11_LC_8_13_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 buf_dds0_i11_LC_8_13_6 (
            .in0(N__32904),
            .in1(N__56854),
            .in2(_gnd_net_),
            .in3(N__50753),
            .lcout(buf_dds0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61898),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_8_13_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_8_13_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i27_LC_8_13_7  (
            .in0(N__30287),
            .in1(N__39754),
            .in2(N__27934),
            .in3(N__37814),
            .lcout(cmd_rdadctmp_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61898),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i5_LC_8_14_0.C_ON=1'b0;
    defparam buf_dds1_i5_LC_8_14_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i5_LC_8_14_0.LUT_INIT=16'b1110001011101110;
    LogicCell40 buf_dds1_i5_LC_8_14_0 (
            .in0(N__28718),
            .in1(N__55403),
            .in2(N__47113),
            .in3(N__63783),
            .lcout(buf_dds1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61912),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i14_LC_8_14_1.C_ON=1'b0;
    defparam buf_dds0_i14_LC_8_14_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i14_LC_8_14_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_dds0_i14_LC_8_14_1 (
            .in0(N__57870),
            .in1(N__50764),
            .in2(N__40564),
            .in3(N__32231),
            .lcout(buf_dds0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i19_LC_8_14_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i19_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i19_LC_8_14_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i19_LC_8_14_2  (
            .in0(N__35988),
            .in1(N__35603),
            .in2(N__27868),
            .in3(N__27828),
            .lcout(buf_adcdata_vac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61912),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i0_LC_8_14_3.C_ON=1'b0;
    defparam buf_dds1_i0_LC_8_14_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i0_LC_8_14_3.LUT_INIT=16'b1110010000000000;
    LogicCell40 buf_dds1_i0_LC_8_14_3 (
            .in0(N__55402),
            .in1(N__37220),
            .in2(N__49150),
            .in3(N__49563),
            .lcout(buf_dds1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i13_LC_8_14_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i13_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i13_LC_8_14_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i13_LC_8_14_6  (
            .in0(N__39341),
            .in1(N__39753),
            .in2(N__28096),
            .in3(N__52319),
            .lcout(buf_adcdata_iac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61912),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i6_LC_8_15_1.C_ON=1'b0;
    defparam buf_dds0_i6_LC_8_15_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i6_LC_8_15_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_dds0_i6_LC_8_15_1 (
            .in0(N__47077),
            .in1(N__50763),
            .in2(_gnd_net_),
            .in3(N__31829),
            .lcout(buf_dds0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61932),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i1_LC_8_15_2.C_ON=1'b0;
    defparam buf_dds1_i1_LC_8_15_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i1_LC_8_15_2.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i1_LC_8_15_2 (
            .in0(N__42125),
            .in1(N__55423),
            .in2(N__52134),
            .in3(N__49570),
            .lcout(buf_dds1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61932),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i19_LC_8_15_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i19_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i19_LC_8_15_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i19_LC_8_15_5  (
            .in0(N__39402),
            .in1(N__39745),
            .in2(N__30303),
            .in3(N__27992),
            .lcout(buf_adcdata_iac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61932),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_4_i16_3_lut_LC_8_15_6.C_ON=1'b0;
    defparam mux_125_Mux_4_i16_3_lut_LC_8_15_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i16_3_lut_LC_8_15_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_125_Mux_4_i16_3_lut_LC_8_15_6 (
            .in0(N__32283),
            .in1(N__27969),
            .in2(_gnd_net_),
            .in3(N__59492),
            .lcout(n16_adj_1778),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_15_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_15_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i22_LC_8_15_7  (
            .in0(N__39403),
            .in1(N__39746),
            .in2(N__31801),
            .in3(N__31676),
            .lcout(buf_adcdata_iac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61932),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_16_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_16_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i14_LC_8_16_3  (
            .in0(N__39360),
            .in1(N__39618),
            .in2(N__41297),
            .in3(N__28075),
            .lcout(buf_adcdata_iac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61948),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i18_LC_8_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i18_LC_8_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i18_LC_8_16_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i18_LC_8_16_4  (
            .in0(N__39617),
            .in1(N__39361),
            .in2(N__30603),
            .in3(N__27927),
            .lcout(buf_adcdata_iac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61948),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_8_16_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_8_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_8_16_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i26_LC_8_16_7  (
            .in0(N__27926),
            .in1(N__39619),
            .in2(N__30460),
            .in3(N__37815),
            .lcout(cmd_rdadctmp_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61948),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_7_i16_3_lut_LC_8_17_0.C_ON=1'b0;
    defparam mux_126_Mux_7_i16_3_lut_LC_8_17_0.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_7_i16_3_lut_LC_8_17_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_7_i16_3_lut_LC_8_17_0 (
            .in0(N__27913),
            .in1(N__32314),
            .in2(_gnd_net_),
            .in3(N__59516),
            .lcout(n16_adj_1713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.SCLK_35_LC_8_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.SCLK_35_LC_8_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.SCLK_35_LC_8_17_1 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_IAC.SCLK_35_LC_8_17_1  (
            .in0(N__39608),
            .in1(N__30436),
            .in2(N__27885),
            .in3(N__30371),
            .lcout(IAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61966),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_17_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i23_LC_8_17_3  (
            .in0(N__37790),
            .in1(N__28055),
            .in2(N__39712),
            .in3(N__28074),
            .lcout(cmd_rdadctmp_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61966),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_8_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_8_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_8_17_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i21_LC_8_17_4  (
            .in0(N__28088),
            .in1(N__39609),
            .in2(N__37258),
            .in3(N__37791),
            .lcout(cmd_rdadctmp_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61966),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_8_17_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_8_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_8_17_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i22_LC_8_17_5  (
            .in0(N__37789),
            .in1(N__28073),
            .in2(N__39711),
            .in3(N__28089),
            .lcout(cmd_rdadctmp_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61966),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_8_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_8_17_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i24_LC_8_17_6  (
            .in0(N__30506),
            .in1(N__39610),
            .in2(N__28060),
            .in3(N__37792),
            .lcout(cmd_rdadctmp_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61966),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i15_LC_8_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i15_LC_8_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i15_LC_8_17_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i15_LC_8_17_7  (
            .in0(N__39334),
            .in1(N__39620),
            .in2(N__46910),
            .in3(N__28059),
            .lcout(buf_adcdata_iac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61966),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_8_18_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_8_18_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i18_LC_8_18_1  (
            .in0(N__29750),
            .in1(N__39632),
            .in2(N__39216),
            .in3(N__37823),
            .lcout(cmd_rdadctmp_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61981),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_8_18_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_8_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_8_18_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i25_LC_8_18_2  (
            .in0(N__37821),
            .in1(N__30452),
            .in2(N__30511),
            .in3(N__39636),
            .lcout(cmd_rdadctmp_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61981),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_8_18_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_8_18_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i17_LC_8_18_5  (
            .in0(N__39209),
            .in1(N__39631),
            .in2(N__34614),
            .in3(N__37822),
            .lcout(cmd_rdadctmp_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61981),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_19_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_19_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_19_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i19_LC_8_19_7  (
            .in0(N__37269),
            .in1(N__39675),
            .in2(N__29757),
            .in3(N__37824),
            .lcout(cmd_rdadctmp_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61995),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7_4_lut_LC_9_2_1 .C_ON=1'b0;
    defparam \ADC_VDC.i7_4_lut_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7_4_lut_LC_9_2_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i7_4_lut_LC_9_2_1  (
            .in0(N__28044),
            .in1(N__28032),
            .in2(N__28021),
            .in3(N__28179),
            .lcout(),
            .ltout(\ADC_VDC.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i11_3_lut_LC_9_2_2 .C_ON=1'b0;
    defparam \ADC_VDC.i11_3_lut_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i11_3_lut_LC_9_2_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \ADC_VDC.i11_3_lut_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__28168),
            .in2(N__28159),
            .in3(N__28156),
            .lcout(\ADC_VDC.adc_state_3_N_1316_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19130_2_lut_LC_9_2_5 .C_ON=1'b0;
    defparam \ADC_VDC.i19130_2_lut_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19130_2_lut_LC_9_2_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i19130_2_lut_LC_9_2_5  (
            .in0(_gnd_net_),
            .in1(N__32849),
            .in2(_gnd_net_),
            .in3(N__32495),
            .lcout(\ADC_VDC.n22055 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i2_LC_9_2_6 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i2_LC_9_2_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i2_LC_9_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ADC_VDC.adc_state_i2_LC_9_2_6  (
            .in0(N__32496),
            .in1(N__33273),
            .in2(_gnd_net_),
            .in3(N__33576),
            .lcout(adc_state_2_adj_1550),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42753),
            .ce(N__28141),
            .sr(N__28108));
    defparam \ADC_VDC.i1_4_lut_LC_9_3_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_LC_9_3_7 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \ADC_VDC.i1_4_lut_LC_9_3_7  (
            .in0(N__28147),
            .in1(N__33575),
            .in2(N__33348),
            .in3(N__30517),
            .lcout(\ADC_VDC.n21871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i3_LC_9_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i3_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i3_LC_9_4_1 .LUT_INIT=16'b0000011110000000;
    LogicCell40 \ADC_VDC.adc_state_i3_LC_9_4_1  (
            .in0(N__33532),
            .in1(N__32485),
            .in2(N__33368),
            .in3(N__32599),
            .lcout(adc_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42717),
            .ce(N__28132),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i14825_3_lut_LC_9_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.i14825_3_lut_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i14825_3_lut_LC_9_4_4 .LUT_INIT=16'b1101110110101010;
    LogicCell40 \ADC_VDC.i14825_3_lut_LC_9_4_4  (
            .in0(N__32833),
            .in1(N__32450),
            .in2(_gnd_net_),
            .in3(N__33531),
            .lcout(),
            .ltout(\ADC_VDC.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_15_LC_9_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_15_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_15_LC_9_4_5 .LUT_INIT=16'b1011101111111010;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_15_LC_9_4_5  (
            .in0(N__33290),
            .in1(N__28121),
            .in2(N__28126),
            .in3(N__32597),
            .lcout(\ADC_VDC.n44_adj_1487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i20180_3_lut_LC_9_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i20180_3_lut_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i20180_3_lut_LC_9_4_7 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \ADC_VDC.i20180_3_lut_LC_9_4_7  (
            .in0(N__33291),
            .in1(N__28122),
            .in2(_gnd_net_),
            .in3(N__32598),
            .lcout(\ADC_VDC.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i0_LC_9_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i0_LC_9_5_0 .LUT_INIT=16'b0001000100110010;
    LogicCell40 \ADC_VDC.adc_state_i0_LC_9_5_0  (
            .in0(N__33314),
            .in1(N__33550),
            .in2(N__32848),
            .in3(N__32700),
            .lcout(\ADC_VDC.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42696),
            .ce(N__30841),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i3_LC_9_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i3_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i3_LC_9_6_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i3_LC_9_6_3  (
            .in0(N__33393),
            .in1(N__31082),
            .in2(N__33741),
            .in3(N__28438),
            .lcout(buf_adcdata_vdc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42749),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_7  (
            .in0(N__28277),
            .in1(N__28426),
            .in2(N__28402),
            .in3(N__32701),
            .lcout(cmd_rdadctmp_9_adj_1565),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42749),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_7_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \ADC_VDC.ADC_DATA_i11_LC_9_7_0  (
            .in0(N__31060),
            .in1(N__33354),
            .in2(N__28258),
            .in3(N__41241),
            .lcout(buf_adcdata_vdc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42694),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_12_LC_9_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_12_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_12_LC_9_7_1 .LUT_INIT=16'b1111001010000000;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_adj_12_LC_9_7_1  (
            .in0(N__32490),
            .in1(N__33551),
            .in2(N__33403),
            .in3(N__32688),
            .lcout(\ADC_VDC.n14120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_7_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i2_LC_9_7_2  (
            .in0(N__31061),
            .in1(N__33355),
            .in2(N__35214),
            .in3(N__28243),
            .lcout(buf_adcdata_vdc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42694),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i5_LC_9_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i5_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i5_LC_9_7_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.ADC_DATA_i5_LC_9_7_5  (
            .in0(N__33353),
            .in1(N__31063),
            .in2(N__28231),
            .in3(N__28206),
            .lcout(buf_adcdata_vdc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42694),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_7_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i16_LC_9_7_7  (
            .in0(N__33352),
            .in1(N__31062),
            .in2(N__43536),
            .in3(N__28195),
            .lcout(buf_adcdata_vdc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42694),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i7_12609_12610_set_LC_9_8_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12609_12610_set_LC_9_8_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i7_12609_12610_set_LC_9_8_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.data_tx_i7_12609_12610_set_LC_9_8_0  (
            .in0(N__36553),
            .in1(_gnd_net_),
            .in2(N__36187),
            .in3(N__31251),
            .lcout(\comm_spi.n15337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53691),
            .ce(),
            .sr(N__41903));
    defparam mux_126_Mux_5_i111_3_lut_LC_9_8_1.C_ON=1'b0;
    defparam mux_126_Mux_5_i111_3_lut_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_5_i111_3_lut_LC_9_8_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_126_Mux_5_i111_3_lut_LC_9_8_1 (
            .in0(N__36919),
            .in1(N__36940),
            .in2(_gnd_net_),
            .in3(N__59326),
            .lcout(n111_adj_1732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_5_i16_3_lut_LC_9_8_2.C_ON=1'b0;
    defparam mux_126_Mux_5_i16_3_lut_LC_9_8_2.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_5_i16_3_lut_LC_9_8_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_126_Mux_5_i16_3_lut_LC_9_8_2 (
            .in0(N__59325),
            .in1(N__28723),
            .in2(_gnd_net_),
            .in3(N__32372),
            .lcout(n16_adj_1728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_6_i16_3_lut_LC_9_8_4.C_ON=1'b0;
    defparam mux_126_Mux_6_i16_3_lut_LC_9_8_4.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_6_i16_3_lut_LC_9_8_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_126_Mux_6_i16_3_lut_LC_9_8_4 (
            .in0(N__59324),
            .in1(N__31323),
            .in2(_gnd_net_),
            .in3(N__31839),
            .lcout(n16_adj_1721),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_6_i19_3_lut_LC_9_8_5.C_ON=1'b0;
    defparam mux_126_Mux_6_i19_3_lut_LC_9_8_5.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_6_i19_3_lut_LC_9_8_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_6_i19_3_lut_LC_9_8_5 (
            .in0(N__28696),
            .in1(N__28671),
            .in2(_gnd_net_),
            .in3(N__59323),
            .lcout(n19_adj_1722),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i13037_2_lut_LC_9_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.i13037_2_lut_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i13037_2_lut_LC_9_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i13037_2_lut_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__32696),
            .in2(_gnd_net_),
            .in3(N__28589),
            .lcout(\ADC_VDC.n15721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i5_12636_12637_reset_LC_9_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12636_12637_reset_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i5_12636_12637_reset_LC_9_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_12636_12637_reset_LC_9_9_0  (
            .in0(N__28879),
            .in1(N__31456),
            .in2(_gnd_net_),
            .in3(N__33771),
            .lcout(\comm_spi.n15365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53690),
            .ce(),
            .sr(N__35236));
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_9_10_0 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_9_10_0 .LUT_INIT=16'b1111001110000000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_LC_9_10_0  (
            .in0(N__32509),
            .in1(N__33574),
            .in2(N__33439),
            .in3(N__32729),
            .lcout(\ADC_VDC.n14092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_LC_9_10_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_LC_9_10_1 .LUT_INIT=16'b1101110111101110;
    LogicCell40 \ADC_VDC.i1_3_lut_LC_9_10_1  (
            .in0(N__28467),
            .in1(N__32508),
            .in2(_gnd_net_),
            .in3(N__30535),
            .lcout(),
            .ltout(\ADC_VDC.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_10_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_10_2 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i34_LC_9_10_2  (
            .in0(N__33410),
            .in1(N__28483),
            .in2(N__28477),
            .in3(N__32730),
            .lcout(cmd_rdadcbuf_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42759),
            .ce(N__28450),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_17_LC_9_10_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_17_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_17_LC_9_10_6 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_adj_17_LC_9_10_6  (
            .in0(N__32507),
            .in1(N__33573),
            .in2(N__33438),
            .in3(N__32728),
            .lcout(n12352),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_9_11_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_9_11_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \comm_spi.RESET_I_0_95_2_lut_LC_9_11_0  (
            .in0(N__36294),
            .in1(_gnd_net_),
            .in2(N__57147),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_857 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20238_4_lut_3_lut_LC_9_11_1 .C_ON=1'b0;
    defparam \comm_spi.i20238_4_lut_3_lut_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20238_4_lut_3_lut_LC_9_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i20238_4_lut_3_lut_LC_9_11_1  (
            .in0(N__28875),
            .in1(N__36295),
            .in2(_gnd_net_),
            .in3(N__57135),
            .lcout(\comm_spi.n24028 ),
            .ltout(\comm_spi.n24028_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i5_12636_12637_set_LC_9_11_2 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12636_12637_set_LC_9_11_2 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i5_12636_12637_set_LC_9_11_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.data_tx_i5_12636_12637_set_LC_9_11_2  (
            .in0(N__31452),
            .in1(_gnd_net_),
            .in2(N__28864),
            .in3(N__33772),
            .lcout(\comm_spi.n15364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53699),
            .ce(),
            .sr(N__36157));
    defparam \comm_spi.i20243_4_lut_3_lut_LC_9_11_3 .C_ON=1'b0;
    defparam \comm_spi.i20243_4_lut_3_lut_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20243_4_lut_3_lut_LC_9_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i20243_4_lut_3_lut_LC_9_11_3  (
            .in0(N__36590),
            .in1(N__45657),
            .in2(_gnd_net_),
            .in3(N__57136),
            .lcout(\comm_spi.n24025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_9_11_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_9_11_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \comm_spi.RESET_I_0_92_2_lut_LC_9_11_4  (
            .in0(N__57131),
            .in1(N__40657),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_854 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_4_i20_3_lut_LC_9_11_7.C_ON=1'b0;
    defparam mux_125_Mux_4_i20_3_lut_LC_9_11_7.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i20_3_lut_LC_9_11_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_4_i20_3_lut_LC_9_11_7 (
            .in0(N__28861),
            .in1(N__28901),
            .in2(_gnd_net_),
            .in3(N__59327),
            .lcout(n20_adj_1781),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_0  (
            .in0(N__35958),
            .in1(N__28769),
            .in2(N__28825),
            .in3(N__33972),
            .lcout(cmd_rdadctmp_20_adj_1528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61871),
            .ce(),
            .sr(_gnd_net_));
    defparam n23306_bdd_4_lut_LC_9_12_1.C_ON=1'b0;
    defparam n23306_bdd_4_lut_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam n23306_bdd_4_lut_LC_9_12_1.LUT_INIT=16'b1100110010111000;
    LogicCell40 n23306_bdd_4_lut_LC_9_12_1 (
            .in0(N__45601),
            .in1(N__43444),
            .in2(N__37462),
            .in3(N__60047),
            .lcout(n23309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19237_3_lut_LC_9_12_2.C_ON=1'b0;
    defparam i19237_3_lut_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam i19237_3_lut_LC_9_12_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 i19237_3_lut_LC_9_12_2 (
            .in0(N__28750),
            .in1(N__28940),
            .in2(_gnd_net_),
            .in3(N__59371),
            .lcout(),
            .ltout(n22164_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20513_LC_9_12_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20513_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20513_LC_9_12_3.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20513_LC_9_12_3 (
            .in0(N__31462),
            .in1(N__60045),
            .in2(N__29071),
            .in3(N__60640),
            .lcout(n23468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_6_i16_3_lut_LC_9_12_4.C_ON=1'b0;
    defparam mux_125_Mux_6_i16_3_lut_LC_9_12_4.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_6_i16_3_lut_LC_9_12_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_6_i16_3_lut_LC_9_12_4 (
            .in0(N__29068),
            .in1(N__32235),
            .in2(_gnd_net_),
            .in3(N__59372),
            .lcout(),
            .ltout(n16_adj_1763_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23366_bdd_4_lut_LC_9_12_5.C_ON=1'b0;
    defparam n23366_bdd_4_lut_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam n23366_bdd_4_lut_LC_9_12_5.LUT_INIT=16'b1100110010111000;
    LogicCell40 n23366_bdd_4_lut_LC_9_12_5 (
            .in0(N__31630),
            .in1(N__29047),
            .in2(N__29035),
            .in3(N__60046),
            .lcout(n23369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_5_i127_3_lut_LC_9_12_6.C_ON=1'b0;
    defparam mux_127_Mux_5_i127_3_lut_LC_9_12_6.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_5_i127_3_lut_LC_9_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_5_i127_3_lut_LC_9_12_6 (
            .in0(N__36918),
            .in1(N__29026),
            .in2(_gnd_net_),
            .in3(N__61395),
            .lcout(comm_buf_2_7_N_575_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i6_LC_9_13_0.C_ON=1'b0;
    defparam buf_cfgRTD_i6_LC_9_13_0.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i6_LC_9_13_0.LUT_INIT=16'b0111001001010000;
    LogicCell40 buf_cfgRTD_i6_LC_9_13_0 (
            .in0(N__48808),
            .in1(N__57861),
            .in2(N__28994),
            .in3(N__40562),
            .lcout(buf_cfgRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i2_LC_9_13_1.C_ON=1'b0;
    defparam buf_cfgRTD_i2_LC_9_13_1.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i2_LC_9_13_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i2_LC_9_13_1 (
            .in0(N__47452),
            .in1(N__48809),
            .in2(_gnd_net_),
            .in3(N__28941),
            .lcout(buf_cfgRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i4_LC_9_13_2.C_ON=1'b0;
    defparam buf_cfgRTD_i4_LC_9_13_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i4_LC_9_13_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 buf_cfgRTD_i4_LC_9_13_2 (
            .in0(N__48807),
            .in1(N__47373),
            .in2(_gnd_net_),
            .in3(N__28900),
            .lcout(buf_cfgRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i12_LC_9_13_3.C_ON=1'b0;
    defparam buf_dds0_i12_LC_9_13_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i12_LC_9_13_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_dds0_i12_LC_9_13_3 (
            .in0(N__47374),
            .in1(N__50722),
            .in2(_gnd_net_),
            .in3(N__32282),
            .lcout(buf_dds0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i5_LC_9_13_4.C_ON=1'b0;
    defparam buf_dds0_i5_LC_9_13_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i5_LC_9_13_4.LUT_INIT=16'b0101000011011000;
    LogicCell40 buf_dds0_i5_LC_9_13_4 (
            .in0(N__50723),
            .in1(N__56569),
            .in2(N__32376),
            .in3(N__57862),
            .lcout(buf_dds0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i19_LC_9_13_5.C_ON=1'b0;
    defparam comm_test_buf_24_i19_LC_9_13_5.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i19_LC_9_13_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_test_buf_24_i19_LC_9_13_5 (
            .in0(N__57860),
            .in1(N__31431),
            .in2(N__62100),
            .in3(N__45421),
            .lcout(comm_test_buf_24_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i10_LC_9_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i10_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i10_LC_9_13_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i10_LC_9_13_6  (
            .in0(N__39421),
            .in1(N__39732),
            .in2(N__29764),
            .in3(N__42056),
            .lcout(buf_adcdata_iac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i11_LC_9_13_7.C_ON=1'b0;
    defparam buf_dds1_i11_LC_9_13_7.SEQ_MODE=4'b1000;
    defparam buf_dds1_i11_LC_9_13_7.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i11_LC_9_13_7 (
            .in0(N__29732),
            .in1(N__55401),
            .in2(N__62101),
            .in3(N__49559),
            .lcout(buf_dds1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61885),
            .ce(),
            .sr(_gnd_net_));
    defparam data_count_i0_i0_LC_9_14_0.C_ON=1'b1;
    defparam data_count_i0_i0_LC_9_14_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i0_LC_9_14_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i0_LC_9_14_0 (
            .in0(_gnd_net_),
            .in1(N__29630),
            .in2(N__49437),
            .in3(_gnd_net_),
            .lcout(data_count_0),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(n20613),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i1_LC_9_14_1.C_ON=1'b1;
    defparam data_count_i0_i1_LC_9_14_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i1_LC_9_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i1_LC_9_14_1 (
            .in0(_gnd_net_),
            .in1(N__29522),
            .in2(_gnd_net_),
            .in3(N__29500),
            .lcout(data_count_1),
            .ltout(),
            .carryin(n20613),
            .carryout(n20614),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i2_LC_9_14_2.C_ON=1'b1;
    defparam data_count_i0_i2_LC_9_14_2.SEQ_MODE=4'b1000;
    defparam data_count_i0_i2_LC_9_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i2_LC_9_14_2 (
            .in0(_gnd_net_),
            .in1(N__29414),
            .in2(_gnd_net_),
            .in3(N__29392),
            .lcout(data_count_2),
            .ltout(),
            .carryin(n20614),
            .carryout(n20615),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i3_LC_9_14_3.C_ON=1'b1;
    defparam data_count_i0_i3_LC_9_14_3.SEQ_MODE=4'b1000;
    defparam data_count_i0_i3_LC_9_14_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i3_LC_9_14_3 (
            .in0(_gnd_net_),
            .in1(N__29309),
            .in2(_gnd_net_),
            .in3(N__29287),
            .lcout(data_count_3),
            .ltout(),
            .carryin(n20615),
            .carryout(n20616),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i4_LC_9_14_4.C_ON=1'b1;
    defparam data_count_i0_i4_LC_9_14_4.SEQ_MODE=4'b1000;
    defparam data_count_i0_i4_LC_9_14_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i4_LC_9_14_4 (
            .in0(_gnd_net_),
            .in1(N__29198),
            .in2(_gnd_net_),
            .in3(N__29179),
            .lcout(data_count_4),
            .ltout(),
            .carryin(n20616),
            .carryout(n20617),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i5_LC_9_14_5.C_ON=1'b1;
    defparam data_count_i0_i5_LC_9_14_5.SEQ_MODE=4'b1000;
    defparam data_count_i0_i5_LC_9_14_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i5_LC_9_14_5 (
            .in0(_gnd_net_),
            .in1(N__29096),
            .in2(_gnd_net_),
            .in3(N__29074),
            .lcout(data_count_5),
            .ltout(),
            .carryin(n20617),
            .carryout(n20618),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i6_LC_9_14_6.C_ON=1'b1;
    defparam data_count_i0_i6_LC_9_14_6.SEQ_MODE=4'b1000;
    defparam data_count_i0_i6_LC_9_14_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i6_LC_9_14_6 (
            .in0(_gnd_net_),
            .in1(N__30161),
            .in2(_gnd_net_),
            .in3(N__30142),
            .lcout(data_count_6),
            .ltout(),
            .carryin(n20618),
            .carryout(n20619),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i7_LC_9_14_7.C_ON=1'b1;
    defparam data_count_i0_i7_LC_9_14_7.SEQ_MODE=4'b1000;
    defparam data_count_i0_i7_LC_9_14_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i7_LC_9_14_7 (
            .in0(_gnd_net_),
            .in1(N__30053),
            .in2(_gnd_net_),
            .in3(N__30034),
            .lcout(data_count_7),
            .ltout(),
            .carryin(n20619),
            .carryout(n20620),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__50013),
            .sr(N__49956));
    defparam data_count_i0_i8_LC_9_15_0.C_ON=1'b1;
    defparam data_count_i0_i8_LC_9_15_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i8_LC_9_15_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i8_LC_9_15_0 (
            .in0(_gnd_net_),
            .in1(N__29951),
            .in2(_gnd_net_),
            .in3(N__29929),
            .lcout(data_count_8),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(n20621),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__50019),
            .sr(N__49957));
    defparam data_count_i0_i9_LC_9_15_1.C_ON=1'b0;
    defparam data_count_i0_i9_LC_9_15_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i9_LC_9_15_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i9_LC_9_15_1 (
            .in0(_gnd_net_),
            .in1(N__29846),
            .in2(_gnd_net_),
            .in3(N__29926),
            .lcout(data_count_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__50019),
            .sr(N__49957));
    defparam i1_2_lut_4_lut_adj_270_LC_9_16_0.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_270_LC_9_16_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_270_LC_9_16_0.LUT_INIT=16'b1100110011000100;
    LogicCell40 i1_2_lut_4_lut_adj_270_LC_9_16_0 (
            .in0(N__55635),
            .in1(N__30560),
            .in2(N__38775),
            .in3(N__50887),
            .lcout(),
            .ltout(n24_adj_1598_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i3_LC_9_16_1.C_ON=1'b0;
    defparam buf_device_acadc_i3_LC_9_16_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i3_LC_9_16_1.LUT_INIT=16'b1111111011111100;
    LogicCell40 buf_device_acadc_i3_LC_9_16_1 (
            .in0(N__40940),
            .in1(N__29824),
            .in2(N__29815),
            .in3(N__43618),
            .lcout(IAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61933),
            .ce(N__36799),
            .sr(N__37141));
    defparam i1_2_lut_4_lut_adj_271_LC_9_16_2.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_271_LC_9_16_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_271_LC_9_16_2.LUT_INIT=16'b1100110011000100;
    LogicCell40 i1_2_lut_4_lut_adj_271_LC_9_16_2 (
            .in0(N__55636),
            .in1(N__29789),
            .in2(N__38776),
            .in3(N__50888),
            .lcout(),
            .ltout(n24_adj_1506_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i4_LC_9_16_3.C_ON=1'b0;
    defparam buf_device_acadc_i4_LC_9_16_3.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i4_LC_9_16_3.LUT_INIT=16'b1111111011111100;
    LogicCell40 buf_device_acadc_i4_LC_9_16_3 (
            .in0(N__62093),
            .in1(N__29770),
            .in2(N__29812),
            .in3(N__43423),
            .lcout(IAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61933),
            .ce(N__36799),
            .sr(N__37141));
    defparam i1_4_lut_LC_9_16_5.C_ON=1'b0;
    defparam i1_4_lut_LC_9_16_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_9_16_5.LUT_INIT=16'b1110010000000000;
    LogicCell40 i1_4_lut_LC_9_16_5 (
            .in0(N__59431),
            .in1(N__49322),
            .in2(N__46123),
            .in3(N__37394),
            .lcout(n11982),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_276_LC_9_16_6.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_276_LC_9_16_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_276_LC_9_16_6.LUT_INIT=16'b1100110011000100;
    LogicCell40 i1_2_lut_4_lut_adj_276_LC_9_16_6 (
            .in0(N__55634),
            .in1(N__38657),
            .in2(N__38774),
            .in3(N__50886),
            .lcout(n24_adj_1503),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_17_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i16_LC_9_17_0  (
            .in0(N__39377),
            .in1(N__39767),
            .in2(N__34385),
            .in3(N__30510),
            .lcout(buf_adcdata_iac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61949),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_9_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_9_17_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i6_LC_9_17_1  (
            .in0(N__39766),
            .in1(N__32160),
            .in2(N__30490),
            .in3(N__37794),
            .lcout(cmd_rdadctmp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61949),
            .ce(),
            .sr(_gnd_net_));
    defparam n23468_bdd_4_lut_LC_9_17_2.C_ON=1'b0;
    defparam n23468_bdd_4_lut_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam n23468_bdd_4_lut_LC_9_17_2.LUT_INIT=16'b1010101011011000;
    LogicCell40 n23468_bdd_4_lut_LC_9_17_2 (
            .in0(N__30469),
            .in1(N__30541),
            .in2(N__30619),
            .in3(N__60095),
            .lcout(n23471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i17_LC_9_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i17_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i17_LC_9_17_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i17_LC_9_17_3  (
            .in0(N__39764),
            .in1(N__39378),
            .in2(N__30267),
            .in3(N__30456),
            .lcout(buf_adcdata_iac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61949),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_264_LC_9_17_4.C_ON=1'b0;
    defparam i1_2_lut_adj_264_LC_9_17_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_264_LC_9_17_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_264_LC_9_17_4 (
            .in0(_gnd_net_),
            .in1(N__31911),
            .in2(_gnd_net_),
            .in3(N__32147),
            .lcout(n13_adj_1591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.DTRIG_39_LC_9_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.DTRIG_39_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.DTRIG_39_LC_9_17_6 .LUT_INIT=16'b1100110011101000;
    LogicCell40 \ADC_IAC.DTRIG_39_LC_9_17_6  (
            .in0(N__30435),
            .in1(N__32148),
            .in2(N__30373),
            .in3(N__39768),
            .lcout(acadc_dtrig_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61949),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_9_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_9_17_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i28_LC_9_17_7  (
            .in0(N__39765),
            .in1(N__37187),
            .in2(N__30304),
            .in3(N__37793),
            .lcout(cmd_rdadctmp_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61949),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_20567_LC_9_18_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20567_LC_9_18_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20567_LC_9_18_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_20567_LC_9_18_0 (
            .in0(N__37047),
            .in1(N__60620),
            .in2(N__30263),
            .in3(N__59428),
            .lcout(n23534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i10_LC_9_18_1.C_ON=1'b0;
    defparam buf_dds0_i10_LC_9_18_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i10_LC_9_18_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 buf_dds0_i10_LC_9_18_1 (
            .in0(N__31854),
            .in1(_gnd_net_),
            .in2(N__47453),
            .in3(N__50770),
            .lcout(buf_dds0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61967),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i15_LC_9_18_4.C_ON=1'b0;
    defparam buf_dds0_i15_LC_9_18_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i15_LC_9_18_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i15_LC_9_18_4 (
            .in0(N__50771),
            .in1(N__57876),
            .in2(N__46663),
            .in3(N__32195),
            .lcout(buf_dds0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61967),
            .ce(),
            .sr(_gnd_net_));
    defparam i19233_3_lut_LC_9_18_6.C_ON=1'b0;
    defparam i19233_3_lut_LC_9_18_6.SEQ_MODE=4'b0000;
    defparam i19233_3_lut_LC_9_18_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i19233_3_lut_LC_9_18_6 (
            .in0(N__30643),
            .in1(N__31853),
            .in2(_gnd_net_),
            .in3(N__59430),
            .lcout(n22160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19234_3_lut_LC_9_18_7.C_ON=1'b0;
    defparam i19234_3_lut_LC_9_18_7.SEQ_MODE=4'b0000;
    defparam i19234_3_lut_LC_9_18_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i19234_3_lut_LC_9_18_7 (
            .in0(N__59429),
            .in1(N__30599),
            .in2(_gnd_net_),
            .in3(N__30564),
            .lcout(n22161),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_9_LC_10_3_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_9_LC_10_3_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_9_LC_10_3_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_9_LC_10_3_3  (
            .in0(_gnd_net_),
            .in1(N__33249),
            .in2(_gnd_net_),
            .in3(N__32590),
            .lcout(\ADC_VDC.n21991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_LC_10_3_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_LC_10_3_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ADC_VDC.i1_2_lut_LC_10_3_4  (
            .in0(N__32591),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33266),
            .lcout(\ADC_VDC.n21707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_3__I_0_56_Mux_1_i10_3_lut_LC_10_3_5 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_3__I_0_56_Mux_1_i10_3_lut_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.adc_state_3__I_0_56_Mux_1_i10_3_lut_LC_10_3_5 .LUT_INIT=16'b0111011101100110;
    LogicCell40 \ADC_VDC.adc_state_3__I_0_56_Mux_1_i10_3_lut_LC_10_3_5  (
            .in0(N__32484),
            .in1(N__33581),
            .in2(_gnd_net_),
            .in3(N__30531),
            .lcout(\ADC_VDC.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i20026_4_lut_LC_10_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.i20026_4_lut_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i20026_4_lut_LC_10_4_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \ADC_VDC.i20026_4_lut_LC_10_4_2  (
            .in0(N__33086),
            .in1(N__30685),
            .in2(N__32641),
            .in3(N__32881),
            .lcout(),
            .ltout(\ADC_VDC.n22404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i35_4_lut_LC_10_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i35_4_lut_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i35_4_lut_LC_10_4_3 .LUT_INIT=16'b1100000001010101;
    LogicCell40 \ADC_VDC.i35_4_lut_LC_10_4_3  (
            .in0(N__32853),
            .in1(N__33151),
            .in2(N__30520),
            .in3(N__32457),
            .lcout(\ADC_VDC.n17 ),
            .ltout(\ADC_VDC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i33_3_lut_LC_10_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.i33_3_lut_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i33_3_lut_LC_10_4_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ADC_VDC.i33_3_lut_LC_10_4_4  (
            .in0(_gnd_net_),
            .in1(N__32852),
            .in2(N__30715),
            .in3(N__33549),
            .lcout(),
            .ltout(\ADC_VDC.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_14_LC_10_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_14_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_14_LC_10_4_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_14_LC_10_4_5  (
            .in0(N__30712),
            .in1(N__33318),
            .in2(N__30703),
            .in3(N__32595),
            .lcout(\ADC_VDC.n21869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i1_LC_10_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i1_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i1_LC_10_4_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.adc_state_i1_LC_10_4_7  (
            .in0(N__30700),
            .in1(N__33319),
            .in2(N__30661),
            .in3(N__32596),
            .lcout(adc_state_1_adj_1551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42698),
            .ce(N__30694),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_6_LC_10_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_6_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_6_LC_10_5_0 .LUT_INIT=16'b1111000001100000;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_6_LC_10_5_0  (
            .in0(N__33534),
            .in1(N__32472),
            .in2(N__33429),
            .in3(N__32605),
            .lcout(\ADC_VDC.n13957 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_13_LC_10_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_13_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_13_LC_10_5_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_13_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__33115),
            .in2(_gnd_net_),
            .in3(N__30819),
            .lcout(\ADC_VDC.n11923 ),
            .ltout(\ADC_VDC.n11923_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_adj_11_LC_10_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_adj_11_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_adj_11_LC_10_5_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.i4_4_lut_adj_11_LC_10_5_2  (
            .in0(N__30832),
            .in1(N__33146),
            .in2(N__30679),
            .in3(N__33008),
            .lcout(\ADC_VDC.n20869 ),
            .ltout(\ADC_VDC.n20869_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i5307_4_lut_LC_10_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.i5307_4_lut_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i5307_4_lut_LC_10_5_3 .LUT_INIT=16'b0011101101001100;
    LogicCell40 \ADC_VDC.i5307_4_lut_LC_10_5_3  (
            .in0(N__32470),
            .in1(N__33533),
            .in2(N__30676),
            .in3(N__32850),
            .lcout(\ADC_VDC.n8031 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.n23528_bdd_4_lut_4_lut_LC_10_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.n23528_bdd_4_lut_4_lut_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.n23528_bdd_4_lut_4_lut_LC_10_5_4 .LUT_INIT=16'b1111010100001100;
    LogicCell40 \ADC_VDC.n23528_bdd_4_lut_4_lut_LC_10_5_4  (
            .in0(N__33536),
            .in1(N__30808),
            .in2(N__33430),
            .in3(N__33157),
            .lcout(\ADC_VDC.n23531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19149_2_lut_LC_10_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i19149_2_lut_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19149_2_lut_LC_10_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i19149_2_lut_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__33535),
            .in2(_gnd_net_),
            .in3(N__30649),
            .lcout(),
            .ltout(\ADC_VDC.n22075_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_16_LC_10_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_16_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_16_LC_10_5_6 .LUT_INIT=16'b1011111100000000;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_16_LC_10_5_6  (
            .in0(N__30862),
            .in1(N__32471),
            .in2(N__30850),
            .in3(N__30847),
            .lcout(\ADC_VDC.n39_adj_1488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_10_LC_10_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_10_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_10_LC_10_5_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_10_LC_10_5_7  (
            .in0(_gnd_net_),
            .in1(N__33066),
            .in2(_gnd_net_),
            .in3(N__33039),
            .lcout(\ADC_VDC.n6_adj_1485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i2_3_lut_LC_10_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.i2_3_lut_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i2_3_lut_LC_10_6_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ADC_VDC.i2_3_lut_LC_10_6_1  (
            .in0(N__32961),
            .in1(N__32976),
            .in2(_gnd_net_),
            .in3(N__32943),
            .lcout(\ADC_VDC.n21859 ),
            .ltout(\ADC_VDC.n21859_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_10_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_10_6_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \ADC_VDC.i1_2_lut_3_lut_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__33116),
            .in2(N__30826),
            .in3(N__33144),
            .lcout(\ADC_VDC.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i20014_4_lut_LC_10_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.i20014_4_lut_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i20014_4_lut_LC_10_6_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \ADC_VDC.i20014_4_lut_LC_10_6_3  (
            .in0(N__33145),
            .in1(N__33117),
            .in2(N__33088),
            .in3(N__33040),
            .lcout(),
            .ltout(\ADC_VDC.n22628_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i20101_4_lut_LC_10_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.i20101_4_lut_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i20101_4_lut_LC_10_6_4 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \ADC_VDC.i20101_4_lut_LC_10_6_4  (
            .in0(N__33548),
            .in1(N__33007),
            .in2(N__30823),
            .in3(N__30820),
            .lcout(\ADC_VDC.n22625 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_LC_10_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_LC_10_6_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \ADC_VDC.i4_4_lut_LC_10_6_6  (
            .in0(N__33041),
            .in1(N__33006),
            .in2(N__33087),
            .in3(N__30802),
            .lcout(\ADC_VDC.n11183 ),
            .ltout(\ADC_VDC.n11183_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_7 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_7  (
            .in0(N__30753),
            .in1(N__30796),
            .in2(N__30763),
            .in3(N__32494),
            .lcout(\ADC_VDC.cmd_rdadctmp_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42697),
            .ce(N__30739),
            .sr(N__30724));
    defparam \comm_spi.imiso_83_12612_12613_reset_LC_10_7_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12612_12613_reset_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imiso_83_12612_12613_reset_LC_10_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.imiso_83_12612_12613_reset_LC_10_7_0  (
            .in0(N__38181),
            .in1(N__38436),
            .in2(_gnd_net_),
            .in3(N__41986),
            .lcout(\comm_spi.n15341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12612_12613_resetC_net ),
            .ce(),
            .sr(N__40629));
    defparam \comm_spi.data_tx_i7_12609_12610_reset_LC_10_8_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12609_12610_reset_LC_10_8_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i7_12609_12610_reset_LC_10_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.data_tx_i7_12609_12610_reset_LC_10_8_0  (
            .in0(N__36183),
            .in1(N__31252),
            .in2(_gnd_net_),
            .in3(N__36552),
            .lcout(\comm_spi.n15338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53666),
            .ce(),
            .sr(N__40630));
    defparam comm_cmd_1__bdd_4_lut_20473_LC_10_9_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20473_LC_10_9_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20473_LC_10_9_0.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20473_LC_10_9_0 (
            .in0(N__59328),
            .in1(N__31234),
            .in2(N__31114),
            .in3(N__60544),
            .lcout(),
            .ltout(n23384_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23384_bdd_4_lut_LC_10_9_1.C_ON=1'b0;
    defparam n23384_bdd_4_lut_LC_10_9_1.SEQ_MODE=4'b0000;
    defparam n23384_bdd_4_lut_LC_10_9_1.LUT_INIT=16'b1111000011001010;
    LogicCell40 n23384_bdd_4_lut_LC_10_9_1 (
            .in0(N__31197),
            .in1(N__31170),
            .in2(N__31135),
            .in3(N__59330),
            .lcout(n23387),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i21_LC_10_9_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i21_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i21_LC_10_9_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i21_LC_10_9_2  (
            .in0(N__31033),
            .in1(N__33387),
            .in2(N__31113),
            .in3(N__31132),
            .lcout(buf_adcdata_vdc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42695),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i13_LC_10_9_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i13_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i13_LC_10_9_3 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ADC_VDC.ADC_DATA_i13_LC_10_9_3  (
            .in0(N__33385),
            .in1(N__31099),
            .in2(N__31073),
            .in3(N__38061),
            .lcout(buf_adcdata_vdc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42695),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i0_LC_10_9_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i0_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i0_LC_10_9_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i0_LC_10_9_4  (
            .in0(N__31032),
            .in1(N__33386),
            .in2(N__37899),
            .in3(N__30964),
            .lcout(buf_adcdata_vdc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42695),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_4_i19_3_lut_LC_10_9_5.C_ON=1'b0;
    defparam mux_126_Mux_4_i19_3_lut_LC_10_9_5.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_4_i19_3_lut_LC_10_9_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_4_i19_3_lut_LC_10_9_5 (
            .in0(N__30946),
            .in1(N__30918),
            .in2(_gnd_net_),
            .in3(N__59329),
            .lcout(),
            .ltout(n19_adj_1734_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20498_LC_10_9_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20498_LC_10_9_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20498_LC_10_9_6.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20498_LC_10_9_6 (
            .in0(N__30889),
            .in1(N__60036),
            .in2(N__30865),
            .in3(N__60545),
            .lcout(n23438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_124_Mux_1_i30_4_lut_4_lut_LC_10_9_7.C_ON=1'b0;
    defparam mux_124_Mux_1_i30_4_lut_4_lut_LC_10_9_7.SEQ_MODE=4'b0000;
    defparam mux_124_Mux_1_i30_4_lut_4_lut_LC_10_9_7.LUT_INIT=16'b1111011111011001;
    LogicCell40 mux_124_Mux_1_i30_4_lut_4_lut_LC_10_9_7 (
            .in0(N__60546),
            .in1(N__61032),
            .in2(N__60090),
            .in3(N__59331),
            .lcout(n30_adj_1805),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_10_10_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_10_10_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i8_LC_10_10_0  (
            .in0(N__35999),
            .in1(N__36113),
            .in2(N__31393),
            .in3(N__34002),
            .lcout(cmd_rdadctmp_8_adj_1540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61845),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_10_10_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_10_10_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i7_LC_10_10_1  (
            .in0(N__33990),
            .in1(N__31389),
            .in2(N__31381),
            .in3(N__36001),
            .lcout(cmd_rdadctmp_7_adj_1541),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61845),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_10_10_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_10_10_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i6_LC_10_10_2  (
            .in0(N__35998),
            .in1(N__33991),
            .in2(N__31369),
            .in3(N__31377),
            .lcout(cmd_rdadctmp_6_adj_1542),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61845),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_10_10_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_10_10_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i5_LC_10_10_3  (
            .in0(N__33989),
            .in1(N__31365),
            .in2(N__31339),
            .in3(N__36000),
            .lcout(cmd_rdadctmp_5_adj_1543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61845),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_10_10_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_10_10_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i4_LC_10_10_4  (
            .in0(N__35997),
            .in1(N__31335),
            .in2(N__34006),
            .in3(N__31356),
            .lcout(cmd_rdadctmp_4_adj_1544),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61845),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i6_LC_10_10_5.C_ON=1'b0;
    defparam buf_dds1_i6_LC_10_10_5.SEQ_MODE=4'b1000;
    defparam buf_dds1_i6_LC_10_10_5.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i6_LC_10_10_5 (
            .in0(N__31322),
            .in1(N__55399),
            .in2(N__49243),
            .in3(N__49503),
            .lcout(buf_dds1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61845),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_10_10_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_10_10_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i9_LC_10_10_6  (
            .in0(N__35421),
            .in1(N__38128),
            .in2(N__39807),
            .in3(N__37840),
            .lcout(cmd_rdadctmp_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61845),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_0_i30_3_lut_LC_10_11_0.C_ON=1'b0;
    defparam mux_127_Mux_0_i30_3_lut_LC_10_11_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_0_i30_3_lut_LC_10_11_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_127_Mux_0_i30_3_lut_LC_10_11_0 (
            .in0(N__31300),
            .in1(N__60989),
            .in2(_gnd_net_),
            .in3(N__37855),
            .lcout(n30_adj_1588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i13_LC_10_11_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i13_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i13_LC_10_11_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i13_LC_10_11_1  (
            .in0(N__35616),
            .in1(N__35962),
            .in2(N__31282),
            .in3(N__38036),
            .lcout(buf_adcdata_vac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61853),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_7_i127_3_lut_LC_10_11_2.C_ON=1'b0;
    defparam mux_127_Mux_7_i127_3_lut_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_7_i127_3_lut_LC_10_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_127_Mux_7_i127_3_lut_LC_10_11_2 (
            .in0(N__61396),
            .in1(N__38352),
            .in2(_gnd_net_),
            .in3(N__31567),
            .lcout(comm_buf_2_7_N_575_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i17_LC_10_11_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i17_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i17_LC_10_11_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i17_LC_10_11_3  (
            .in0(N__35617),
            .in1(N__35963),
            .in2(N__31555),
            .in3(N__48602),
            .lcout(buf_adcdata_vac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61853),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i20_LC_10_11_5.C_ON=1'b0;
    defparam comm_test_buf_24_i20_LC_10_11_5.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i20_LC_10_11_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_test_buf_24_i20_LC_10_11_5 (
            .in0(N__57863),
            .in1(N__31417),
            .in2(N__44707),
            .in3(N__45414),
            .lcout(comm_test_buf_24_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61853),
            .ce(),
            .sr(_gnd_net_));
    defparam i19236_3_lut_LC_10_11_7.C_ON=1'b0;
    defparam i19236_3_lut_LC_10_11_7.SEQ_MODE=4'b0000;
    defparam i19236_3_lut_LC_10_11_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i19236_3_lut_LC_10_11_7 (
            .in0(N__31516),
            .in1(N__31485),
            .in2(_gnd_net_),
            .in3(N__59020),
            .lcout(n22163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i4_12632_12633_set_LC_10_12_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12632_12633_set_LC_10_12_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i4_12632_12633_set_LC_10_12_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_tx_i4_12632_12633_set_LC_10_12_0  (
            .in0(N__36238),
            .in1(N__34045),
            .in2(_gnd_net_),
            .in3(N__51052),
            .lcout(\comm_spi.n15360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53710),
            .ce(),
            .sr(N__31441));
    defparam mux_125_Mux_3_i111_3_lut_LC_10_12_1.C_ON=1'b0;
    defparam mux_125_Mux_3_i111_3_lut_LC_10_12_1.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i111_3_lut_LC_10_12_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_3_i111_3_lut_LC_10_12_1 (
            .in0(N__31432),
            .in1(N__34257),
            .in2(_gnd_net_),
            .in3(N__59261),
            .lcout(n111_adj_1794),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_3_i111_3_lut_LC_10_12_2.C_ON=1'b0;
    defparam mux_126_Mux_3_i111_3_lut_LC_10_12_2.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_3_i111_3_lut_LC_10_12_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_126_Mux_3_i111_3_lut_LC_10_12_2 (
            .in0(N__59262),
            .in1(N__34178),
            .in2(_gnd_net_),
            .in3(N__34258),
            .lcout(n111_adj_1744),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_4_i111_3_lut_LC_10_12_4.C_ON=1'b0;
    defparam mux_125_Mux_4_i111_3_lut_LC_10_12_4.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i111_3_lut_LC_10_12_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_125_Mux_4_i111_3_lut_LC_10_12_4 (
            .in0(N__59263),
            .in1(N__31416),
            .in2(_gnd_net_),
            .in3(N__34245),
            .lcout(n111_adj_1785),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_4_i111_3_lut_LC_10_12_6.C_ON=1'b0;
    defparam mux_126_Mux_4_i111_3_lut_LC_10_12_6.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_4_i111_3_lut_LC_10_12_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_126_Mux_4_i111_3_lut_LC_10_12_6 (
            .in0(N__59264),
            .in1(N__34091),
            .in2(_gnd_net_),
            .in3(N__34246),
            .lcout(n111_adj_1737),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_289_LC_10_13_0.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_289_LC_10_13_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_289_LC_10_13_0.LUT_INIT=16'b1100110010001100;
    LogicCell40 i1_2_lut_4_lut_adj_289_LC_10_13_0 (
            .in0(N__50893),
            .in1(N__31644),
            .in2(N__55651),
            .in3(N__38757),
            .lcout(),
            .ltout(n24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i7_LC_10_13_1.C_ON=1'b0;
    defparam buf_device_acadc_i7_LC_10_13_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i7_LC_10_13_1.LUT_INIT=16'b1111111011111010;
    LogicCell40 buf_device_acadc_i7_LC_10_13_1 (
            .in0(N__31573),
            .in1(N__40561),
            .in2(N__31693),
            .in3(N__43611),
            .lcout(VAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61872),
            .ce(N__36798),
            .sr(N__37126));
    defparam mux_125_Mux_6_i17_3_lut_LC_10_13_2.C_ON=1'b0;
    defparam mux_125_Mux_6_i17_3_lut_LC_10_13_2.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_6_i17_3_lut_LC_10_13_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_6_i17_3_lut_LC_10_13_2 (
            .in0(N__31683),
            .in1(N__31643),
            .in2(_gnd_net_),
            .in3(N__59265),
            .lcout(n17_adj_1764),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_64_LC_10_13_3.C_ON=1'b0;
    defparam i1_4_lut_adj_64_LC_10_13_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_64_LC_10_13_3.LUT_INIT=16'b1110010000000000;
    LogicCell40 i1_4_lut_adj_64_LC_10_13_3 (
            .in0(N__59267),
            .in1(N__55822),
            .in2(N__40429),
            .in3(N__37405),
            .lcout(),
            .ltout(n11981_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i8_LC_10_13_4.C_ON=1'b0;
    defparam buf_device_acadc_i8_LC_10_13_4.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i8_LC_10_13_4.LUT_INIT=16'b1111111011111100;
    LogicCell40 buf_device_acadc_i8_LC_10_13_4 (
            .in0(N__46621),
            .in1(N__31579),
            .in2(N__31621),
            .in3(N__43422),
            .lcout(VAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61872),
            .ce(N__36798),
            .sr(N__37126));
    defparam i1_2_lut_4_lut_adj_292_LC_10_13_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_292_LC_10_13_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_292_LC_10_13_5.LUT_INIT=16'b1111110100000000;
    LogicCell40 i1_2_lut_4_lut_adj_292_LC_10_13_5 (
            .in0(N__55626),
            .in1(N__50892),
            .in2(N__38772),
            .in3(N__31595),
            .lcout(n24_adj_1576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_57_LC_10_13_6.C_ON=1'b0;
    defparam i1_4_lut_adj_57_LC_10_13_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_57_LC_10_13_6.LUT_INIT=16'b1010000010001000;
    LogicCell40 i1_4_lut_adj_57_LC_10_13_6 (
            .in0(N__37404),
            .in1(N__49214),
            .in2(N__36346),
            .in3(N__59266),
            .lcout(n11986),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10511_3_lut_LC_10_13_7.C_ON=1'b0;
    defparam i10511_3_lut_LC_10_13_7.SEQ_MODE=4'b0000;
    defparam i10511_3_lut_LC_10_13_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i10511_3_lut_LC_10_13_7 (
            .in0(N__40425),
            .in1(N__46620),
            .in2(_gnd_net_),
            .in3(N__46202),
            .lcout(n13237),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20548_LC_10_14_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20548_LC_10_14_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20548_LC_10_14_0.LUT_INIT=16'b1110011011000100;
    LogicCell40 comm_cmd_1__bdd_4_lut_20548_LC_10_14_0 (
            .in0(N__60041),
            .in1(N__60587),
            .in2(N__50221),
            .in3(N__31723),
            .lcout(),
            .ltout(n23510_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23510_bdd_4_lut_LC_10_14_1.C_ON=1'b0;
    defparam n23510_bdd_4_lut_LC_10_14_1.SEQ_MODE=4'b0000;
    defparam n23510_bdd_4_lut_LC_10_14_1.LUT_INIT=16'b1111000011001010;
    LogicCell40 n23510_bdd_4_lut_LC_10_14_1 (
            .in0(N__41482),
            .in1(N__44365),
            .in2(N__31741),
            .in3(N__60042),
            .lcout(),
            .ltout(n23513_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1663271_i1_3_lut_LC_10_14_2.C_ON=1'b0;
    defparam i1663271_i1_3_lut_LC_10_14_2.SEQ_MODE=4'b0000;
    defparam i1663271_i1_3_lut_LC_10_14_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1663271_i1_3_lut_LC_10_14_2 (
            .in0(_gnd_net_),
            .in1(N__31738),
            .in2(N__31729),
            .in3(N__61055),
            .lcout(),
            .ltout(n30_adj_1759_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_7_i127_3_lut_LC_10_14_3.C_ON=1'b0;
    defparam mux_125_Mux_7_i127_3_lut_LC_10_14_3.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_7_i127_3_lut_LC_10_14_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_125_Mux_7_i127_3_lut_LC_10_14_3 (
            .in0(_gnd_net_),
            .in1(N__31708),
            .in2(N__31726),
            .in3(N__61397),
            .lcout(comm_buf_0_7_N_543_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_7_i26_3_lut_LC_10_14_4.C_ON=1'b0;
    defparam mux_125_Mux_7_i26_3_lut_LC_10_14_4.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_7_i26_3_lut_LC_10_14_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_125_Mux_7_i26_3_lut_LC_10_14_4 (
            .in0(N__47293),
            .in1(N__59268),
            .in2(_gnd_net_),
            .in3(N__31716),
            .lcout(n26_adj_1758),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_end_302_LC_10_14_5.C_ON=1'b0;
    defparam eis_end_302_LC_10_14_5.SEQ_MODE=4'b1000;
    defparam eis_end_302_LC_10_14_5.LUT_INIT=16'b1011100010101010;
    LogicCell40 eis_end_302_LC_10_14_5 (
            .in0(N__31717),
            .in1(N__39173),
            .in2(N__34705),
            .in3(N__31699),
            .lcout(eis_end),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_end_302C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_7_i112_3_lut_LC_10_14_6.C_ON=1'b0;
    defparam mux_125_Mux_7_i112_3_lut_LC_10_14_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_7_i112_3_lut_LC_10_14_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_125_Mux_7_i112_3_lut_LC_10_14_6 (
            .in0(N__38351),
            .in1(N__36880),
            .in2(_gnd_net_),
            .in3(N__60588),
            .lcout(n112_adj_1762),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_10_15_0.C_ON=1'b0;
    defparam i24_4_lut_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_10_15_0.LUT_INIT=16'b0111110000101100;
    LogicCell40 i24_4_lut_LC_10_15_0 (
            .in0(N__45787),
            .in1(N__34782),
            .in2(N__34699),
            .in3(N__49435),
            .lcout(n17_adj_1742),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_272_LC_10_15_1.C_ON=1'b0;
    defparam i2_4_lut_adj_272_LC_10_15_1.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_272_LC_10_15_1.LUT_INIT=16'b0000001000000000;
    LogicCell40 i2_4_lut_adj_272_LC_10_15_1 (
            .in0(N__45781),
            .in1(N__31762),
            .in2(N__34796),
            .in3(N__34274),
            .lcout(),
            .ltout(n21946_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20133_3_lut_4_lut_LC_10_15_2.C_ON=1'b0;
    defparam i20133_3_lut_4_lut_LC_10_15_2.SEQ_MODE=4'b0000;
    defparam i20133_3_lut_4_lut_LC_10_15_2.LUT_INIT=16'b1111000001110111;
    LogicCell40 i20133_3_lut_4_lut_LC_10_15_2 (
            .in0(N__34783),
            .in1(N__45782),
            .in2(N__31702),
            .in3(N__34685),
            .lcout(n21880),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i34_3_lut_LC_10_15_3.C_ON=1'b0;
    defparam i34_3_lut_LC_10_15_3.SEQ_MODE=4'b0000;
    defparam i34_3_lut_LC_10_15_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 i34_3_lut_LC_10_15_3 (
            .in0(N__49436),
            .in1(N__34784),
            .in2(_gnd_net_),
            .in3(N__41370),
            .lcout(),
            .ltout(n13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i2_LC_10_15_4.C_ON=1'b0;
    defparam eis_state_i2_LC_10_15_4.SEQ_MODE=4'b1010;
    defparam eis_state_i2_LC_10_15_4.LUT_INIT=16'b1110110001100100;
    LogicCell40 eis_state_i2_LC_10_15_4 (
            .in0(N__45790),
            .in1(N__34686),
            .in2(N__31810),
            .in3(N__31807),
            .lcout(eis_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i2C_net),
            .ce(N__34423),
            .sr(N__39178));
    defparam i19812_2_lut_LC_10_15_5.C_ON=1'b0;
    defparam i19812_2_lut_LC_10_15_5.SEQ_MODE=4'b0000;
    defparam i19812_2_lut_LC_10_15_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 i19812_2_lut_LC_10_15_5 (
            .in0(N__34781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34275),
            .lcout(n22395),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20187_2_lut_3_lut_LC_10_15_6.C_ON=1'b0;
    defparam i20187_2_lut_3_lut_LC_10_15_6.SEQ_MODE=4'b0000;
    defparam i20187_2_lut_3_lut_LC_10_15_6.LUT_INIT=16'b0000000000000101;
    LogicCell40 i20187_2_lut_3_lut_LC_10_15_6 (
            .in0(N__45788),
            .in1(_gnd_net_),
            .in2(N__34698),
            .in3(N__39171),
            .lcout(n22120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20166_3_lut_LC_10_15_7.C_ON=1'b0;
    defparam i20166_3_lut_LC_10_15_7.SEQ_MODE=4'b0000;
    defparam i20166_3_lut_LC_10_15_7.LUT_INIT=16'b0111011111111111;
    LogicCell40 i20166_3_lut_LC_10_15_7 (
            .in0(N__31747),
            .in1(N__34678),
            .in2(_gnd_net_),
            .in3(N__45789),
            .lcout(n12369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i21_LC_10_16_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i21_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i21_LC_10_16_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i21_LC_10_16_0  (
            .in0(N__39772),
            .in1(N__39398),
            .in2(N__32122),
            .in3(N__38606),
            .lcout(buf_adcdata_iac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61914),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i3_LC_10_16_1.C_ON=1'b0;
    defparam buf_dds1_i3_LC_10_16_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i3_LC_10_16_1.LUT_INIT=16'b1011111110110000;
    LogicCell40 buf_dds1_i3_LC_10_16_1 (
            .in0(N__48943),
            .in1(N__63778),
            .in2(N__55400),
            .in3(N__36860),
            .lcout(buf_dds1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61914),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_10_16_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_10_16_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i30_LC_10_16_2  (
            .in0(N__39773),
            .in1(N__31778),
            .in2(N__32121),
            .in3(N__37836),
            .lcout(cmd_rdadctmp_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61914),
            .ce(),
            .sr(_gnd_net_));
    defparam i19796_2_lut_3_lut_LC_10_16_4.C_ON=1'b0;
    defparam i19796_2_lut_3_lut_LC_10_16_4.SEQ_MODE=4'b0000;
    defparam i19796_2_lut_3_lut_LC_10_16_4.LUT_INIT=16'b0011111100000000;
    LogicCell40 i19796_2_lut_3_lut_LC_10_16_4 (
            .in0(_gnd_net_),
            .in1(N__32146),
            .in2(N__31918),
            .in3(N__34672),
            .lcout(n22312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_265_LC_10_16_5.C_ON=1'b0;
    defparam i24_4_lut_adj_265_LC_10_16_5.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_265_LC_10_16_5.LUT_INIT=16'b1111110010101100;
    LogicCell40 i24_4_lut_adj_265_LC_10_16_5 (
            .in0(N__43843),
            .in1(N__31761),
            .in2(N__34791),
            .in3(N__38872),
            .lcout(n11_adj_1592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_10_16_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_10_16_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i7_LC_10_16_6  (
            .in0(N__39774),
            .in1(N__32161),
            .in2(N__38160),
            .in3(N__37837),
            .lcout(cmd_rdadctmp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61914),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_206_LC_10_16_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_206_LC_10_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_206_LC_10_16_7.LUT_INIT=16'b0100000001000000;
    LogicCell40 i1_2_lut_3_lut_adj_206_LC_10_16_7 (
            .in0(N__34671),
            .in1(N__31914),
            .in2(N__32149),
            .in3(_gnd_net_),
            .lcout(n17633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_adj_49_LC_10_17_2 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_adj_49_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_adj_49_LC_10_17_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VAC.i1_2_lut_adj_49_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__31912),
            .in2(_gnd_net_),
            .in3(N__32142),
            .lcout(iac_raw_buf_N_823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i7_LC_10_17_3.C_ON=1'b0;
    defparam buf_dds0_i7_LC_10_17_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i7_LC_10_17_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_dds0_i7_LC_10_17_3 (
            .in0(N__47521),
            .in1(N__50754),
            .in2(_gnd_net_),
            .in3(N__32312),
            .lcout(buf_dds0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61934),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_10_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_10_17_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i29_LC_10_17_4  (
            .in0(N__32114),
            .in1(N__37188),
            .in2(N__39808),
            .in3(N__37795),
            .lcout(cmd_rdadctmp_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61934),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.DTRIG_39_LC_10_17_5 .C_ON=1'b0;
    defparam \ADC_VAC.DTRIG_39_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.DTRIG_39_LC_10_17_5 .LUT_INIT=16'b1010101011101000;
    LogicCell40 \ADC_VAC.DTRIG_39_LC_10_17_5  (
            .in0(N__31913),
            .in1(N__32101),
            .in2(N__32011),
            .in3(N__36002),
            .lcout(acadc_dtrig_v),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61934),
            .ce(),
            .sr(_gnd_net_));
    defparam n23534_bdd_4_lut_LC_10_17_6.C_ON=1'b0;
    defparam n23534_bdd_4_lut_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam n23534_bdd_4_lut_LC_10_17_6.LUT_INIT=16'b1100110010111000;
    LogicCell40 n23534_bdd_4_lut_LC_10_17_6 (
            .in0(N__31890),
            .in1(N__31861),
            .in2(N__50644),
            .in3(N__60564),
            .lcout(n22177),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i10_LC_10_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i10_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i10_LC_10_18_0 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \SIG_DDS.tmp_buf_i10_LC_10_18_0  (
            .in0(N__50549),
            .in1(N__31855),
            .in2(N__32332),
            .in3(N__50415),
            .lcout(\SIG_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61950),
            .ce(N__42208),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i6_LC_10_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i6_LC_10_18_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i6_LC_10_18_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i6_LC_10_18_2  (
            .in0(N__50552),
            .in1(N__50414),
            .in2(N__32341),
            .in3(N__31840),
            .lcout(\SIG_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61950),
            .ce(N__42208),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i4_LC_10_18_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i4_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i4_LC_10_18_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i4_LC_10_18_4  (
            .in0(N__50550),
            .in1(N__50413),
            .in2(N__37438),
            .in3(N__47269),
            .lcout(\SIG_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61950),
            .ce(N__42208),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i5_LC_10_18_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i5_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i5_LC_10_18_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \SIG_DDS.tmp_buf_i5_LC_10_18_5  (
            .in0(N__50411),
            .in1(N__50551),
            .in2(N__32380),
            .in3(N__32347),
            .lcout(\SIG_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61950),
            .ce(N__42208),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i9_LC_10_18_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i9_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i9_LC_10_18_6 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \SIG_DDS.tmp_buf_i9_LC_10_18_6  (
            .in0(N__50640),
            .in1(N__50554),
            .in2(N__32170),
            .in3(N__50416),
            .lcout(\SIG_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61950),
            .ce(N__42208),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i7_LC_10_18_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i7_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i7_LC_10_18_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i7_LC_10_18_7  (
            .in0(N__50412),
            .in1(N__50553),
            .in2(N__32323),
            .in3(N__32313),
            .lcout(\SIG_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61950),
            .ce(N__42208),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i12_LC_10_19_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i12_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i12_LC_10_19_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \SIG_DDS.tmp_buf_i12_LC_10_19_0  (
            .in0(N__50544),
            .in1(N__50407),
            .in2(N__32293),
            .in3(N__32887),
            .lcout(\SIG_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61968),
            .ce(N__42206),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i13_LC_10_19_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i13_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i13_LC_10_19_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i13_LC_10_19_2  (
            .in0(N__50545),
            .in1(N__50408),
            .in2(N__32260),
            .in3(N__55549),
            .lcout(\SIG_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61968),
            .ce(N__42206),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i14_LC_10_19_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i14_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i14_LC_10_19_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i14_LC_10_19_4  (
            .in0(N__50546),
            .in1(N__50409),
            .in2(N__32251),
            .in3(N__32242),
            .lcout(\SIG_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61968),
            .ce(N__42206),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i15_LC_10_19_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i15_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i15_LC_10_19_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i15_LC_10_19_6  (
            .in0(N__50547),
            .in1(N__50410),
            .in2(N__32212),
            .in3(N__32196),
            .lcout(tmp_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61968),
            .ce(N__42206),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i8_LC_10_19_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i8_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i8_LC_10_19_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \SIG_DDS.tmp_buf_i8_LC_10_19_7  (
            .in0(N__50406),
            .in1(N__50548),
            .in2(N__40236),
            .in3(N__32176),
            .lcout(\SIG_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61968),
            .ce(N__42206),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i11_LC_10_20_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i11_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i11_LC_10_20_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i11_LC_10_20_0  (
            .in0(N__50543),
            .in1(N__50403),
            .in2(N__32923),
            .in3(N__32911),
            .lcout(\SIG_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61982),
            .ce(N__42207),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19141_2_lut_LC_11_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.i19141_2_lut_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19141_2_lut_LC_11_4_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ADC_VDC.i19141_2_lut_LC_11_4_0  (
            .in0(N__32854),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33577),
            .lcout(\ADC_VDC.n22067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19137_2_lut_LC_11_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.i19137_2_lut_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19137_2_lut_LC_11_4_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i19137_2_lut_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__33010),
            .in2(_gnd_net_),
            .in3(N__33043),
            .lcout(\ADC_VDC.n22063 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_LC_11_4_5 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_LC_11_4_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \RTD.i2_3_lut_LC_11_4_5  (
            .in0(N__35096),
            .in1(N__35061),
            .in2(_gnd_net_),
            .in3(N__35080),
            .lcout(\RTD.n20050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_7_LC_11_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_7_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_7_LC_11_5_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_7_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__33579),
            .in2(_gnd_net_),
            .in3(N__32851),
            .lcout(),
            .ltout(\ADC_VDC.n35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i14816_4_lut_LC_11_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.i14816_4_lut_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i14816_4_lut_LC_11_5_3 .LUT_INIT=16'b1011101101010000;
    LogicCell40 \ADC_VDC.i14816_4_lut_LC_11_5_3  (
            .in0(N__32702),
            .in1(N__32749),
            .in2(N__32752),
            .in3(N__33379),
            .lcout(\ADC_VDC.n17542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_8_LC_11_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_8_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_8_LC_11_5_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_8_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(N__33578),
            .in2(_gnd_net_),
            .in3(N__32459),
            .lcout(\ADC_VDC.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i24_4_lut_LC_11_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i24_4_lut_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i24_4_lut_LC_11_5_6 .LUT_INIT=16'b1010101001110010;
    LogicCell40 \ADC_VDC.i24_4_lut_LC_11_5_6  (
            .in0(N__33378),
            .in1(N__32460),
            .in2(N__32743),
            .in3(N__32703),
            .lcout(\ADC_VDC.n17565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7 .LUT_INIT=16'b0100101001101010;
    LogicCell40 \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7  (
            .in0(N__32458),
            .in1(N__33580),
            .in2(N__33431),
            .in3(N__33163),
            .lcout(\ADC_VDC.n23528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.bit_cnt_3791__i0_LC_11_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3791__i0_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i0_LC_11_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i0_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__33150),
            .in2(_gnd_net_),
            .in3(N__33121),
            .lcout(\ADC_VDC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\ADC_VDC.n20812 ),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \ADC_VDC.bit_cnt_3791__i1_LC_11_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3791__i1_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i1_LC_11_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i1_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__33118),
            .in2(_gnd_net_),
            .in3(N__33091),
            .lcout(\ADC_VDC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n20812 ),
            .carryout(\ADC_VDC.n20813 ),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \ADC_VDC.bit_cnt_3791__i2_LC_11_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3791__i2_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i2_LC_11_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i2_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__33076),
            .in2(_gnd_net_),
            .in3(N__33046),
            .lcout(\ADC_VDC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n20813 ),
            .carryout(\ADC_VDC.n20814 ),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \ADC_VDC.bit_cnt_3791__i3_LC_11_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3791__i3_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i3_LC_11_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i3_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__33042),
            .in2(_gnd_net_),
            .in3(N__33013),
            .lcout(\ADC_VDC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n20814 ),
            .carryout(\ADC_VDC.n20815 ),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \ADC_VDC.bit_cnt_3791__i4_LC_11_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3791__i4_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i4_LC_11_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i4_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__33009),
            .in2(_gnd_net_),
            .in3(N__32980),
            .lcout(\ADC_VDC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n20815 ),
            .carryout(\ADC_VDC.n20816 ),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \ADC_VDC.bit_cnt_3791__i5_LC_11_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3791__i5_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i5_LC_11_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i5_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__32977),
            .in2(_gnd_net_),
            .in3(N__32965),
            .lcout(\ADC_VDC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n20816 ),
            .carryout(\ADC_VDC.n20817 ),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \ADC_VDC.bit_cnt_3791__i6_LC_11_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3791__i6_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i6_LC_11_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i6_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__32962),
            .in2(_gnd_net_),
            .in3(N__32950),
            .lcout(\ADC_VDC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n20817 ),
            .carryout(\ADC_VDC.n20818 ),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \ADC_VDC.bit_cnt_3791__i7_LC_11_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.bit_cnt_3791__i7_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3791__i7_LC_11_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3791__i7_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__32944),
            .in2(_gnd_net_),
            .in3(N__32947),
            .lcout(\ADC_VDC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42690),
            .ce(N__32932),
            .sr(N__33781));
    defparam \comm_spi.data_tx_i4_12632_12633_reset_LC_11_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12632_12633_reset_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i4_12632_12633_reset_LC_11_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_12632_12633_reset_LC_11_7_0  (
            .in0(N__34035),
            .in1(N__36231),
            .in2(_gnd_net_),
            .in3(N__51045),
            .lcout(\comm_spi.n15361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53602),
            .ce(),
            .sr(N__36274));
    defparam mux_127_Mux_3_i19_3_lut_LC_11_8_0.C_ON=1'b0;
    defparam mux_127_Mux_3_i19_3_lut_LC_11_8_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_3_i19_3_lut_LC_11_8_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_3_i19_3_lut_LC_11_8_0 (
            .in0(N__33748),
            .in1(N__33644),
            .in2(_gnd_net_),
            .in3(N__59398),
            .lcout(),
            .ltout(n19_adj_1703_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_3_i22_3_lut_LC_11_8_1.C_ON=1'b0;
    defparam mux_127_Mux_3_i22_3_lut_LC_11_8_1.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_3_i22_3_lut_LC_11_8_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_127_Mux_3_i22_3_lut_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(N__33689),
            .in2(N__33724),
            .in3(N__60008),
            .lcout(),
            .ltout(n22_adj_1704_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_3_i30_3_lut_LC_11_8_2.C_ON=1'b0;
    defparam mux_127_Mux_3_i30_3_lut_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_3_i30_3_lut_LC_11_8_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_127_Mux_3_i30_3_lut_LC_11_8_2 (
            .in0(_gnd_net_),
            .in1(N__33721),
            .in2(N__33703),
            .in3(N__61013),
            .lcout(n30_adj_1705),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i1_LC_11_8_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i1_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i1_LC_11_8_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i1_LC_11_8_3  (
            .in0(N__35625),
            .in1(N__35927),
            .in2(N__33805),
            .in3(N__33606),
            .lcout(buf_adcdata_vac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61830),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_8_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_8_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i3_LC_11_8_4  (
            .in0(N__33690),
            .in1(N__39404),
            .in2(N__35388),
            .in3(N__39817),
            .lcout(buf_adcdata_iac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61830),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_8_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_8_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i3_LC_11_8_5  (
            .in0(N__33645),
            .in1(N__35928),
            .in2(N__35629),
            .in3(N__33676),
            .lcout(buf_adcdata_vac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61830),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_3_lut_4_lut_LC_11_8_6.C_ON=1'b0;
    defparam i3_3_lut_4_lut_LC_11_8_6.SEQ_MODE=4'b0000;
    defparam i3_3_lut_4_lut_LC_11_8_6.LUT_INIT=16'b0000000000001000;
    LogicCell40 i3_3_lut_4_lut_LC_11_8_6 (
            .in0(N__54609),
            .in1(N__64079),
            .in2(N__54424),
            .in3(N__63076),
            .lcout(n8_adj_1755),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_1_i19_3_lut_LC_11_9_0.C_ON=1'b0;
    defparam mux_127_Mux_1_i19_3_lut_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_1_i19_3_lut_LC_11_9_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_1_i19_3_lut_LC_11_9_0 (
            .in0(N__33631),
            .in1(N__33602),
            .in2(_gnd_net_),
            .in3(N__59250),
            .lcout(),
            .ltout(n19_adj_1710_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_1_i22_3_lut_LC_11_9_1.C_ON=1'b0;
    defparam mux_127_Mux_1_i22_3_lut_LC_11_9_1.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_1_i22_3_lut_LC_11_9_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_127_Mux_1_i22_3_lut_LC_11_9_1 (
            .in0(_gnd_net_),
            .in1(N__36086),
            .in2(N__34066),
            .in3(N__60040),
            .lcout(),
            .ltout(n22_adj_1711_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_1_i30_3_lut_LC_11_9_2.C_ON=1'b0;
    defparam mux_127_Mux_1_i30_3_lut_LC_11_9_2.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_1_i30_3_lut_LC_11_9_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_127_Mux_1_i30_3_lut_LC_11_9_2 (
            .in0(_gnd_net_),
            .in1(N__34063),
            .in2(N__34051),
            .in3(N__61056),
            .lcout(),
            .ltout(n30_adj_1712_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_1_i127_3_lut_LC_11_9_3.C_ON=1'b0;
    defparam mux_127_Mux_1_i127_3_lut_LC_11_9_3.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_1_i127_3_lut_LC_11_9_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_127_Mux_1_i127_3_lut_LC_11_9_3 (
            .in0(_gnd_net_),
            .in1(N__41867),
            .in2(N__34048),
            .in3(N__61398),
            .lcout(comm_buf_2_7_N_575_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20233_4_lut_3_lut_LC_11_9_4 .C_ON=1'b0;
    defparam \comm_spi.i20233_4_lut_3_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20233_4_lut_3_lut_LC_11_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.i20233_4_lut_3_lut_LC_11_9_4  (
            .in0(N__34023),
            .in1(N__57177),
            .in2(_gnd_net_),
            .in3(N__46078),
            .lcout(\comm_spi.n24031 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_3_i127_3_lut_LC_11_9_5.C_ON=1'b0;
    defparam mux_127_Mux_3_i127_3_lut_LC_11_9_5.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_3_i127_3_lut_LC_11_9_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_3_i127_3_lut_LC_11_9_5 (
            .in0(N__34186),
            .in1(N__34012),
            .in2(_gnd_net_),
            .in3(N__61399),
            .lcout(comm_buf_2_7_N_575_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_11_9_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_11_9_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i9_LC_11_9_6  (
            .in0(N__35990),
            .in1(N__33797),
            .in2(N__36126),
            .in3(N__33993),
            .lcout(cmd_rdadctmp_9_adj_1539),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61834),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_11_9_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_11_9_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i10_LC_11_9_7  (
            .in0(N__33992),
            .in1(N__36029),
            .in2(N__33804),
            .in3(N__35991),
            .lcout(cmd_rdadctmp_10_adj_1538),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61834),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_6_i2_3_lut_LC_11_10_0.C_ON=1'b0;
    defparam mux_134_Mux_6_i2_3_lut_LC_11_10_0.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_6_i2_3_lut_LC_11_10_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_134_Mux_6_i2_3_lut_LC_11_10_0 (
            .in0(N__36342),
            .in1(N__40753),
            .in2(_gnd_net_),
            .in3(N__54422),
            .lcout(),
            .ltout(n2_adj_1666_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i6_LC_11_10_1.C_ON=1'b0;
    defparam comm_tx_buf_i6_LC_11_10_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i6_LC_11_10_1.LUT_INIT=16'b1111101001000100;
    LogicCell40 comm_tx_buf_i6_LC_11_10_1 (
            .in0(N__54611),
            .in1(N__34123),
            .in2(N__33784),
            .in3(N__34204),
            .lcout(comm_tx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61840),
            .ce(N__46426),
            .sr(N__46348));
    defparam i20030_2_lut_LC_11_10_2.C_ON=1'b0;
    defparam i20030_2_lut_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam i20030_2_lut_LC_11_10_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i20030_2_lut_LC_11_10_2 (
            .in0(_gnd_net_),
            .in1(N__37990),
            .in2(_gnd_net_),
            .in3(N__54420),
            .lcout(n22295),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_6_i4_3_lut_LC_11_10_3.C_ON=1'b0;
    defparam mux_134_Mux_6_i4_3_lut_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_6_i4_3_lut_LC_11_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_134_Mux_6_i4_3_lut_LC_11_10_3 (
            .in0(N__54421),
            .in1(N__43126),
            .in2(_gnd_net_),
            .in3(N__53800),
            .lcout(n4_adj_1667),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_6_i1_3_lut_LC_11_10_5.C_ON=1'b0;
    defparam mux_134_Mux_6_i1_3_lut_LC_11_10_5.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_6_i1_3_lut_LC_11_10_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_134_Mux_6_i1_3_lut_LC_11_10_5 (
            .in0(N__49239),
            .in1(N__40503),
            .in2(_gnd_net_),
            .in3(N__54423),
            .lcout(n1_adj_1665),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10505_3_lut_LC_11_10_6.C_ON=1'b0;
    defparam i10505_3_lut_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam i10505_3_lut_LC_11_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i10505_3_lut_LC_11_10_6 (
            .in0(N__36341),
            .in1(N__40517),
            .in2(_gnd_net_),
            .in3(N__46204),
            .lcout(n13231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_11_10_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_11_10_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.RESET_I_0_101_2_lut_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__57178),
            .in2(_gnd_net_),
            .in3(N__36200),
            .lcout(\comm_spi.data_tx_7__N_865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i1_LC_11_11_0.C_ON=1'b0;
    defparam comm_test_buf_24_i1_LC_11_11_0.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i1_LC_11_11_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_test_buf_24_i1_LC_11_11_0 (
            .in0(N__36693),
            .in1(N__52144),
            .in2(_gnd_net_),
            .in3(N__38278),
            .lcout(comm_test_buf_24_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam comm_test_buf_24_i2_LC_11_11_1.C_ON=1'b0;
    defparam comm_test_buf_24_i2_LC_11_11_1.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i2_LC_11_11_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_test_buf_24_i2_LC_11_11_1 (
            .in0(N__52936),
            .in1(N__36697),
            .in2(_gnd_net_),
            .in3(N__40867),
            .lcout(comm_test_buf_24_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam comm_test_buf_24_i4_LC_11_11_2.C_ON=1'b0;
    defparam comm_test_buf_24_i4_LC_11_11_2.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i4_LC_11_11_2.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_test_buf_24_i4_LC_11_11_2 (
            .in0(N__36695),
            .in1(_gnd_net_),
            .in2(N__56109),
            .in3(N__36301),
            .lcout(comm_test_buf_24_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam comm_test_buf_24_i6_LC_11_11_3.C_ON=1'b0;
    defparam comm_test_buf_24_i6_LC_11_11_3.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i6_LC_11_11_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_test_buf_24_i6_LC_11_11_3 (
            .in0(N__49230),
            .in1(N__36699),
            .in2(_gnd_net_),
            .in3(N__34072),
            .lcout(comm_test_buf_24_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam comm_test_buf_24_i7_LC_11_11_4.C_ON=1'b0;
    defparam comm_test_buf_24_i7_LC_11_11_4.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i7_LC_11_11_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_test_buf_24_i7_LC_11_11_4 (
            .in0(N__36696),
            .in1(N__55848),
            .in2(_gnd_net_),
            .in3(N__34237),
            .lcout(comm_test_buf_24_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam comm_test_buf_24_i0_LC_11_11_5.C_ON=1'b0;
    defparam comm_test_buf_24_i0_LC_11_11_5.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i0_LC_11_11_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_test_buf_24_i0_LC_11_11_5 (
            .in0(N__43198),
            .in1(_gnd_net_),
            .in2(N__49141),
            .in3(N__36700),
            .lcout(comm_test_buf_24_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam comm_test_buf_24_i3_LC_11_11_6.C_ON=1'b0;
    defparam comm_test_buf_24_i3_LC_11_11_6.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i3_LC_11_11_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_test_buf_24_i3_LC_11_11_6 (
            .in0(N__36694),
            .in1(N__49326),
            .in2(_gnd_net_),
            .in3(N__46093),
            .lcout(comm_test_buf_24_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam comm_test_buf_24_i5_LC_11_11_7.C_ON=1'b0;
    defparam comm_test_buf_24_i5_LC_11_11_7.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i5_LC_11_11_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_test_buf_24_i5_LC_11_11_7 (
            .in0(N__56587),
            .in1(N__36698),
            .in2(_gnd_net_),
            .in3(N__37969),
            .lcout(comm_test_buf_24_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61846),
            .ce(N__41188),
            .sr(N__34156));
    defparam n23324_bdd_4_lut_LC_11_12_0.C_ON=1'b0;
    defparam n23324_bdd_4_lut_LC_11_12_0.SEQ_MODE=4'b0000;
    defparam n23324_bdd_4_lut_LC_11_12_0.LUT_INIT=16'b1100110010111000;
    LogicCell40 n23324_bdd_4_lut_LC_11_12_0 (
            .in0(N__34136),
            .in1(N__34354),
            .in2(N__40240),
            .in3(N__60462),
            .lcout(n23327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_20419_LC_11_12_1.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_20419_LC_11_12_1.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_20419_LC_11_12_1.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_index_1__bdd_4_lut_20419_LC_11_12_1 (
            .in0(N__54610),
            .in1(N__34228),
            .in2(N__34216),
            .in3(N__51837),
            .lcout(n23294),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_0_i127_3_lut_LC_11_12_2.C_ON=1'b0;
    defparam mux_127_Mux_0_i127_3_lut_LC_11_12_2.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_0_i127_3_lut_LC_11_12_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_0_i127_3_lut_LC_11_12_2 (
            .in0(N__48986),
            .in1(N__34195),
            .in2(_gnd_net_),
            .in3(N__61400),
            .lcout(comm_buf_2_7_N_575_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i112_3_lut_LC_11_12_3.C_ON=1'b0;
    defparam mux_125_Mux_3_i112_3_lut_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i112_3_lut_LC_11_12_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_125_Mux_3_i112_3_lut_LC_11_12_3 (
            .in0(N__60461),
            .in1(N__34179),
            .in2(_gnd_net_),
            .in3(N__34162),
            .lcout(n112_adj_1795),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12822_2_lut_3_lut_LC_11_12_4.C_ON=1'b0;
    defparam i12822_2_lut_3_lut_LC_11_12_4.SEQ_MODE=4'b0000;
    defparam i12822_2_lut_3_lut_LC_11_12_4.LUT_INIT=16'b1100110010001000;
    LogicCell40 i12822_2_lut_3_lut_LC_11_12_4 (
            .in0(N__64097),
            .in1(N__41187),
            .in2(_gnd_net_),
            .in3(N__62607),
            .lcout(n15545),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i8_LC_11_12_6.C_ON=1'b0;
    defparam buf_dds1_i8_LC_11_12_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i8_LC_11_12_6.LUT_INIT=16'b1101100000000000;
    LogicCell40 buf_dds1_i8_LC_11_12_6 (
            .in0(N__55430),
            .in1(N__43955),
            .in2(N__34143),
            .in3(N__49537),
            .lcout(buf_dds1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61854),
            .ce(),
            .sr(_gnd_net_));
    defparam i12815_2_lut_3_lut_LC_11_12_7.C_ON=1'b0;
    defparam i12815_2_lut_3_lut_LC_11_12_7.SEQ_MODE=4'b0000;
    defparam i12815_2_lut_3_lut_LC_11_12_7.LUT_INIT=16'b1010101010001000;
    LogicCell40 i12815_2_lut_3_lut_LC_11_12_7 (
            .in0(N__36777),
            .in1(N__62603),
            .in2(_gnd_net_),
            .in3(N__64096),
            .lcout(n15538),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i8_LC_11_13_0.C_ON=1'b0;
    defparam comm_test_buf_24_i8_LC_11_13_0.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i8_LC_11_13_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_test_buf_24_i8_LC_11_13_0 (
            .in0(N__43939),
            .in1(N__49106),
            .in2(_gnd_net_),
            .in3(N__36671),
            .lcout(comm_test_buf_24_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_test_buf_24_i11_LC_11_13_1.C_ON=1'b0;
    defparam comm_test_buf_24_i11_LC_11_13_1.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i11_LC_11_13_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_test_buf_24_i11_LC_11_13_1 (
            .in0(N__36665),
            .in1(N__62086),
            .in2(_gnd_net_),
            .in3(N__49318),
            .lcout(comm_test_buf_24_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_test_buf_24_i13_LC_11_13_2.C_ON=1'b0;
    defparam comm_test_buf_24_i13_LC_11_13_2.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i13_LC_11_13_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_test_buf_24_i13_LC_11_13_2 (
            .in0(N__45335),
            .in1(N__56583),
            .in2(_gnd_net_),
            .in3(N__36669),
            .lcout(comm_test_buf_24_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_test_buf_24_i9_LC_11_13_3.C_ON=1'b0;
    defparam comm_test_buf_24_i9_LC_11_13_3.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i9_LC_11_13_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_test_buf_24_i9_LC_11_13_3 (
            .in0(N__52138),
            .in1(_gnd_net_),
            .in2(N__44630),
            .in3(N__36692),
            .lcout(comm_test_buf_24_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_test_buf_24_i10_LC_11_13_4.C_ON=1'b0;
    defparam comm_test_buf_24_i10_LC_11_13_4.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i10_LC_11_13_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_test_buf_24_i10_LC_11_13_4 (
            .in0(N__52934),
            .in1(N__40935),
            .in2(_gnd_net_),
            .in3(N__36668),
            .lcout(comm_test_buf_24_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_test_buf_24_i12_LC_11_13_5.C_ON=1'b0;
    defparam comm_test_buf_24_i12_LC_11_13_5.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i12_LC_11_13_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_test_buf_24_i12_LC_11_13_5 (
            .in0(N__36666),
            .in1(N__44703),
            .in2(_gnd_net_),
            .in3(N__56110),
            .lcout(comm_test_buf_24_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_test_buf_24_i14_LC_11_13_6.C_ON=1'b0;
    defparam comm_test_buf_24_i14_LC_11_13_6.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i14_LC_11_13_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_test_buf_24_i14_LC_11_13_6 (
            .in0(N__49231),
            .in1(N__40539),
            .in2(_gnd_net_),
            .in3(N__36670),
            .lcout(comm_test_buf_24_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_test_buf_24_i15_LC_11_13_7.C_ON=1'b0;
    defparam comm_test_buf_24_i15_LC_11_13_7.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i15_LC_11_13_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_test_buf_24_i15_LC_11_13_7 (
            .in0(N__36667),
            .in1(_gnd_net_),
            .in2(N__46629),
            .in3(N__55823),
            .lcout(comm_test_buf_24_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61862),
            .ce(N__44044),
            .sr(N__41338));
    defparam comm_cmd_0__bdd_4_lut_20562_LC_11_14_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20562_LC_11_14_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20562_LC_11_14_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_20562_LC_11_14_0 (
            .in0(N__34343),
            .in1(N__60589),
            .in2(N__43842),
            .in3(N__59113),
            .lcout(n23522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_20409_LC_11_14_1.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20409_LC_11_14_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20409_LC_11_14_1.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_20409_LC_11_14_1 (
            .in0(N__59114),
            .in1(N__34386),
            .in2(N__37083),
            .in3(N__60627),
            .lcout(n23324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i8_LC_11_14_2.C_ON=1'b0;
    defparam req_data_cnt_i8_LC_11_14_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i8_LC_11_14_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i8_LC_11_14_2 (
            .in0(N__34344),
            .in1(N__48870),
            .in2(_gnd_net_),
            .in3(N__51361),
            .lcout(req_data_cnt_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61873),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_256_LC_11_14_3.C_ON=1'b0;
    defparam i3_4_lut_adj_256_LC_11_14_3.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_256_LC_11_14_3.LUT_INIT=16'b0111101111011110;
    LogicCell40 i3_4_lut_adj_256_LC_11_14_3 (
            .in0(N__49756),
            .in1(N__50065),
            .in2(N__34345),
            .in3(N__60689),
            .lcout(),
            .ltout(n19_adj_1727_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_11_14_4.C_ON=1'b0;
    defparam i13_4_lut_LC_11_14_4.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_11_14_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_LC_11_14_4 (
            .in0(N__44056),
            .in1(N__44128),
            .in2(N__34327),
            .in3(N__38452),
            .lcout(),
            .ltout(n29_adj_1770_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_11_14_5.C_ON=1'b0;
    defparam i1_3_lut_LC_11_14_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_11_14_5.LUT_INIT=16'b1100110011001111;
    LogicCell40 i1_3_lut_LC_11_14_5 (
            .in0(_gnd_net_),
            .in1(N__38867),
            .in2(N__34324),
            .in3(N__41464),
            .lcout(n16_adj_1683),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i13_LC_11_14_6.C_ON=1'b0;
    defparam req_data_cnt_i13_LC_11_14_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i13_LC_11_14_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i13_LC_11_14_6 (
            .in0(N__60690),
            .in1(N__55276),
            .in2(_gnd_net_),
            .in3(N__51360),
            .lcout(req_data_cnt_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61873),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_6_i111_3_lut_LC_11_14_7.C_ON=1'b0;
    defparam mux_126_Mux_6_i111_3_lut_LC_11_14_7.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_6_i111_3_lut_LC_11_14_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_126_Mux_6_i111_3_lut_LC_11_14_7 (
            .in0(N__59115),
            .in1(_gnd_net_),
            .in2(N__34320),
            .in3(N__34293),
            .lcout(n111_adj_1726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14917_4_lut_LC_11_15_0.C_ON=1'b0;
    defparam i14917_4_lut_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam i14917_4_lut_LC_11_15_0.LUT_INIT=16'b1100010111001111;
    LogicCell40 i14917_4_lut_LC_11_15_0 (
            .in0(N__43835),
            .in1(N__34276),
            .in2(N__34695),
            .in3(N__41551),
            .lcout(),
            .ltout(n17642_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i0_LC_11_15_1.C_ON=1'b0;
    defparam eis_state_i0_LC_11_15_1.SEQ_MODE=4'b1010;
    defparam eis_state_i0_LC_11_15_1.LUT_INIT=16'b1111101000010001;
    LogicCell40 eis_state_i0_LC_11_15_1 (
            .in0(N__34774),
            .in1(N__34670),
            .in2(N__34261),
            .in3(N__34555),
            .lcout(eis_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__34419),
            .sr(N__39172));
    defparam eis_state_1__bdd_4_lut_4_lut_LC_11_15_2.C_ON=1'b0;
    defparam eis_state_1__bdd_4_lut_4_lut_LC_11_15_2.SEQ_MODE=4'b0000;
    defparam eis_state_1__bdd_4_lut_4_lut_LC_11_15_2.LUT_INIT=16'b0100101011101010;
    LogicCell40 eis_state_1__bdd_4_lut_4_lut_LC_11_15_2 (
            .in0(N__45797),
            .in1(N__34561),
            .in2(N__34786),
            .in3(N__34548),
            .lcout(n23330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3823_3_lut_3_lut_4_lut_LC_11_15_4.C_ON=1'b0;
    defparam i3823_3_lut_3_lut_4_lut_LC_11_15_4.SEQ_MODE=4'b0000;
    defparam i3823_3_lut_3_lut_4_lut_LC_11_15_4.LUT_INIT=16'b0010000000000000;
    LogicCell40 i3823_3_lut_3_lut_4_lut_LC_11_15_4 (
            .in0(N__45798),
            .in1(N__39132),
            .in2(N__34787),
            .in3(N__34549),
            .lcout(iac_raw_buf_N_821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_4_lut_LC_11_15_6.C_ON=1'b0;
    defparam i2_4_lut_4_lut_4_lut_LC_11_15_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_4_lut_LC_11_15_6.LUT_INIT=16'b0000000001010001;
    LogicCell40 i2_4_lut_4_lut_4_lut_LC_11_15_6 (
            .in0(N__34666),
            .in1(N__45783),
            .in2(N__34785),
            .in3(N__39131),
            .lcout(n12394),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i1_LC_11_15_7.C_ON=1'b0;
    defparam eis_state_i1_LC_11_15_7.SEQ_MODE=4'b1010;
    defparam eis_state_i1_LC_11_15_7.LUT_INIT=16'b1010101010101110;
    LogicCell40 eis_state_i1_LC_11_15_7 (
            .in0(N__34429),
            .in1(N__45799),
            .in2(N__34795),
            .in3(N__41371),
            .lcout(eis_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__34419),
            .sr(N__39172));
    defparam buf_device_acadc_i2_LC_11_16_1.C_ON=1'b0;
    defparam buf_device_acadc_i2_LC_11_16_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i2_LC_11_16_1.LUT_INIT=16'b1111111011101110;
    LogicCell40 buf_device_acadc_i2_LC_11_16_1 (
            .in0(N__37018),
            .in1(N__34804),
            .in2(N__44647),
            .in3(N__43617),
            .lcout(IAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61901),
            .ce(N__36790),
            .sr(N__37134));
    defparam buf_device_acadc_i6_LC_11_16_2.C_ON=1'b0;
    defparam buf_device_acadc_i6_LC_11_16_2.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i6_LC_11_16_2.LUT_INIT=16'b1111111111111000;
    LogicCell40 buf_device_acadc_i6_LC_11_16_2 (
            .in0(N__43616),
            .in1(N__45326),
            .in2(N__34402),
            .in3(N__37012),
            .lcout(VAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61901),
            .ce(N__36790),
            .sr(N__37134));
    defparam i16467_2_lut_3_lut_LC_11_16_4.C_ON=1'b0;
    defparam i16467_2_lut_3_lut_LC_11_16_4.SEQ_MODE=4'b0000;
    defparam i16467_2_lut_3_lut_LC_11_16_4.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16467_2_lut_3_lut_LC_11_16_4 (
            .in0(N__64109),
            .in1(N__52107),
            .in2(_gnd_net_),
            .in3(N__62604),
            .lcout(n14_adj_1613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16445_2_lut_3_lut_LC_11_16_6.C_ON=1'b0;
    defparam i16445_2_lut_3_lut_LC_11_16_6.SEQ_MODE=4'b0000;
    defparam i16445_2_lut_3_lut_LC_11_16_6.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16445_2_lut_3_lut_LC_11_16_6 (
            .in0(N__64111),
            .in1(N__56570),
            .in2(_gnd_net_),
            .in3(N__62605),
            .lcout(n14_adj_1661),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_77_LC_11_16_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_77_LC_11_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_77_LC_11_16_7.LUT_INIT=16'b0000000000100010;
    LogicCell40 i1_2_lut_3_lut_adj_77_LC_11_16_7 (
            .in0(N__45325),
            .in1(N__62606),
            .in2(_gnd_net_),
            .in3(N__64110),
            .lcout(n14_adj_1660),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_335_LC_11_17_0.C_ON=1'b0;
    defparam i1_4_lut_adj_335_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_335_LC_11_17_0.LUT_INIT=16'b1100100000001000;
    LogicCell40 i1_4_lut_adj_335_LC_11_17_0 (
            .in0(N__52143),
            .in1(N__37382),
            .in2(N__59514),
            .in3(N__38311),
            .lcout(n11980),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i9_LC_11_17_1.C_ON=1'b0;
    defparam data_index_i9_LC_11_17_1.SEQ_MODE=4'b1000;
    defparam data_index_i9_LC_11_17_1.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i9_LC_11_17_1 (
            .in0(N__63526),
            .in1(N__44515),
            .in2(N__57747),
            .in3(N__44497),
            .lcout(data_index_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61915),
            .ce(),
            .sr(_gnd_net_));
    defparam i20191_3_lut_4_lut_LC_11_17_2.C_ON=1'b0;
    defparam i20191_3_lut_4_lut_LC_11_17_2.SEQ_MODE=4'b0000;
    defparam i20191_3_lut_4_lut_LC_11_17_2.LUT_INIT=16'b0000000000010101;
    LogicCell40 i20191_3_lut_4_lut_LC_11_17_2 (
            .in0(N__45800),
            .in1(N__34696),
            .in2(N__34797),
            .in3(N__39130),
            .lcout(n12450),
            .ltout(n12450_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20174_2_lut_LC_11_17_3.C_ON=1'b0;
    defparam i20174_2_lut_LC_11_17_3.SEQ_MODE=4'b0000;
    defparam i20174_2_lut_LC_11_17_3.LUT_INIT=16'b0101000001010000;
    LogicCell40 i20174_2_lut_LC_11_17_3 (
            .in0(N__34697),
            .in1(_gnd_net_),
            .in2(N__34618),
            .in3(_gnd_net_),
            .lcout(n15439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i12_LC_11_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i12_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i12_LC_11_17_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i12_LC_11_17_4  (
            .in0(N__39762),
            .in1(N__39370),
            .in2(N__37254),
            .in3(N__36977),
            .lcout(buf_adcdata_iac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61915),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i21_LC_11_17_5.C_ON=1'b0;
    defparam comm_test_buf_24_i21_LC_11_17_5.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i21_LC_11_17_5.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_test_buf_24_i21_LC_11_17_5 (
            .in0(N__57661),
            .in1(N__45327),
            .in2(N__36955),
            .in3(N__45426),
            .lcout(comm_test_buf_24_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61915),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i8_LC_11_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i8_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i8_LC_11_17_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i8_LC_11_17_6  (
            .in0(N__39763),
            .in1(N__39371),
            .in2(N__34615),
            .in3(N__46946),
            .lcout(buf_adcdata_iac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61915),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i0_LC_11_18_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i0_LC_11_18_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i0_LC_11_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i0_LC_11_18_0 (
            .in0(_gnd_net_),
            .in1(N__49412),
            .in2(N__39982),
            .in3(_gnd_net_),
            .lcout(acadc_skipcnt_0),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(n20637),
            .clk(INVacadc_skipcnt_i0_i0C_net),
            .ce(N__35171),
            .sr(N__34573));
    defparam add_70_2_THRU_CRY_0_LC_11_18_1.C_ON=1'b1;
    defparam add_70_2_THRU_CRY_0_LC_11_18_1.SEQ_MODE=4'b0000;
    defparam add_70_2_THRU_CRY_0_LC_11_18_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_70_2_THRU_CRY_0_LC_11_18_1 (
            .in0(_gnd_net_),
            .in1(N__64807),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n20637),
            .carryout(n20637_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_70_2_THRU_CRY_1_LC_11_18_2.C_ON=1'b1;
    defparam add_70_2_THRU_CRY_1_LC_11_18_2.SEQ_MODE=4'b0000;
    defparam add_70_2_THRU_CRY_1_LC_11_18_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_70_2_THRU_CRY_1_LC_11_18_2 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__64852),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n20637_THRU_CRY_0_THRU_CO),
            .carryout(n20637_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_70_2_THRU_CRY_2_LC_11_18_3.C_ON=1'b1;
    defparam add_70_2_THRU_CRY_2_LC_11_18_3.SEQ_MODE=4'b0000;
    defparam add_70_2_THRU_CRY_2_LC_11_18_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_70_2_THRU_CRY_2_LC_11_18_3 (
            .in0(_gnd_net_),
            .in1(N__64811),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n20637_THRU_CRY_1_THRU_CO),
            .carryout(n20637_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_70_2_THRU_CRY_3_LC_11_18_4.C_ON=1'b1;
    defparam add_70_2_THRU_CRY_3_LC_11_18_4.SEQ_MODE=4'b0000;
    defparam add_70_2_THRU_CRY_3_LC_11_18_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_70_2_THRU_CRY_3_LC_11_18_4 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__64853),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n20637_THRU_CRY_2_THRU_CO),
            .carryout(n20637_THRU_CRY_3_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_70_2_THRU_CRY_4_LC_11_18_5.C_ON=1'b1;
    defparam add_70_2_THRU_CRY_4_LC_11_18_5.SEQ_MODE=4'b0000;
    defparam add_70_2_THRU_CRY_4_LC_11_18_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_70_2_THRU_CRY_4_LC_11_18_5 (
            .in0(_gnd_net_),
            .in1(N__64815),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n20637_THRU_CRY_3_THRU_CO),
            .carryout(n20637_THRU_CRY_4_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_70_2_THRU_CRY_5_LC_11_18_6.C_ON=1'b1;
    defparam add_70_2_THRU_CRY_5_LC_11_18_6.SEQ_MODE=4'b0000;
    defparam add_70_2_THRU_CRY_5_LC_11_18_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_70_2_THRU_CRY_5_LC_11_18_6 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__64854),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n20637_THRU_CRY_4_THRU_CO),
            .carryout(n20637_THRU_CRY_5_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_70_2_THRU_CRY_6_LC_11_18_7.C_ON=1'b1;
    defparam add_70_2_THRU_CRY_6_LC_11_18_7.SEQ_MODE=4'b0000;
    defparam add_70_2_THRU_CRY_6_LC_11_18_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_70_2_THRU_CRY_6_LC_11_18_7 (
            .in0(_gnd_net_),
            .in1(N__64819),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n20637_THRU_CRY_5_THRU_CO),
            .carryout(n20637_THRU_CRY_6_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i1_LC_11_19_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i1_LC_11_19_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i1_LC_11_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i1_LC_11_19_0 (
            .in0(_gnd_net_),
            .in1(N__44010),
            .in2(_gnd_net_),
            .in3(N__34813),
            .lcout(acadc_skipcnt_1),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(n20638),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i2_LC_11_19_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i2_LC_11_19_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i2_LC_11_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i2_LC_11_19_1 (
            .in0(_gnd_net_),
            .in1(N__38961),
            .in2(_gnd_net_),
            .in3(N__34810),
            .lcout(acadc_skipcnt_2),
            .ltout(),
            .carryin(n20638),
            .carryout(n20639),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i3_LC_11_19_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i3_LC_11_19_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i3_LC_11_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i3_LC_11_19_2 (
            .in0(_gnd_net_),
            .in1(N__41526),
            .in2(_gnd_net_),
            .in3(N__34807),
            .lcout(acadc_skipcnt_3),
            .ltout(),
            .carryin(n20639),
            .carryout(n20640),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i4_LC_11_19_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i4_LC_11_19_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i4_LC_11_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i4_LC_11_19_3 (
            .in0(_gnd_net_),
            .in1(N__43986),
            .in2(_gnd_net_),
            .in3(N__34840),
            .lcout(acadc_skipcnt_4),
            .ltout(),
            .carryin(n20640),
            .carryout(n20641),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i5_LC_11_19_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i5_LC_11_19_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i5_LC_11_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i5_LC_11_19_4 (
            .in0(_gnd_net_),
            .in1(N__41157),
            .in2(_gnd_net_),
            .in3(N__34837),
            .lcout(acadc_skipcnt_5),
            .ltout(),
            .carryin(n20641),
            .carryout(n20642),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i6_LC_11_19_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i6_LC_11_19_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i6_LC_11_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i6_LC_11_19_5 (
            .in0(_gnd_net_),
            .in1(N__39957),
            .in2(_gnd_net_),
            .in3(N__34834),
            .lcout(acadc_skipcnt_6),
            .ltout(),
            .carryin(n20642),
            .carryout(n20643),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i7_LC_11_19_6.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i7_LC_11_19_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i7_LC_11_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i7_LC_11_19_6 (
            .in0(_gnd_net_),
            .in1(N__38979),
            .in2(_gnd_net_),
            .in3(N__34831),
            .lcout(acadc_skipcnt_7),
            .ltout(),
            .carryin(n20643),
            .carryout(n20644),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i8_LC_11_19_7.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i8_LC_11_19_7.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i8_LC_11_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i8_LC_11_19_7 (
            .in0(_gnd_net_),
            .in1(N__41601),
            .in2(_gnd_net_),
            .in3(N__34828),
            .lcout(acadc_skipcnt_8),
            .ltout(),
            .carryin(n20644),
            .carryout(n20645),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__35188),
            .sr(N__35154));
    defparam acadc_skipcnt_i0_i9_LC_11_20_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i9_LC_11_20_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i9_LC_11_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i9_LC_11_20_0 (
            .in0(_gnd_net_),
            .in1(N__37329),
            .in2(_gnd_net_),
            .in3(N__34825),
            .lcout(acadc_skipcnt_9),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(n20646),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__35187),
            .sr(N__35155));
    defparam acadc_skipcnt_i0_i10_LC_11_20_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i10_LC_11_20_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i10_LC_11_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i10_LC_11_20_1 (
            .in0(_gnd_net_),
            .in1(N__38925),
            .in2(_gnd_net_),
            .in3(N__34822),
            .lcout(acadc_skipcnt_10),
            .ltout(),
            .carryin(n20646),
            .carryout(n20647),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__35187),
            .sr(N__35155));
    defparam acadc_skipcnt_i0_i11_LC_11_20_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i11_LC_11_20_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i11_LC_11_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i11_LC_11_20_2 (
            .in0(_gnd_net_),
            .in1(N__37299),
            .in2(_gnd_net_),
            .in3(N__34819),
            .lcout(acadc_skipcnt_11),
            .ltout(),
            .carryin(n20647),
            .carryout(n20648),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__35187),
            .sr(N__35155));
    defparam acadc_skipcnt_i0_i12_LC_11_20_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i12_LC_11_20_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i12_LC_11_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i12_LC_11_20_3 (
            .in0(_gnd_net_),
            .in1(N__38943),
            .in2(_gnd_net_),
            .in3(N__34816),
            .lcout(acadc_skipcnt_12),
            .ltout(),
            .carryin(n20648),
            .carryout(n20649),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__35187),
            .sr(N__35155));
    defparam acadc_skipcnt_i0_i13_LC_11_20_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i13_LC_11_20_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i13_LC_11_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i13_LC_11_20_4 (
            .in0(_gnd_net_),
            .in1(N__38835),
            .in2(_gnd_net_),
            .in3(N__35197),
            .lcout(acadc_skipcnt_13),
            .ltout(),
            .carryin(n20649),
            .carryout(n20650),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__35187),
            .sr(N__35155));
    defparam acadc_skipcnt_i0_i14_LC_11_20_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i14_LC_11_20_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i14_LC_11_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i14_LC_11_20_5 (
            .in0(_gnd_net_),
            .in1(N__37314),
            .in2(_gnd_net_),
            .in3(N__35194),
            .lcout(acadc_skipcnt_14),
            .ltout(),
            .carryin(n20650),
            .carryout(n20651),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__35187),
            .sr(N__35155));
    defparam acadc_skipcnt_i0_i15_LC_11_20_6.C_ON=1'b0;
    defparam acadc_skipcnt_i0_i15_LC_11_20_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i15_LC_11_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i15_LC_11_20_6 (
            .in0(_gnd_net_),
            .in1(N__37347),
            .in2(_gnd_net_),
            .in3(N__35191),
            .lcout(acadc_skipcnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__35187),
            .sr(N__35155));
    defparam clk_RTD_290_LC_12_3_0.C_ON=1'b0;
    defparam clk_RTD_290_LC_12_3_0.SEQ_MODE=4'b1000;
    defparam clk_RTD_290_LC_12_3_0.LUT_INIT=16'b0110011010101010;
    LogicCell40 clk_RTD_290_LC_12_3_0 (
            .in0(N__34885),
            .in1(N__36465),
            .in2(_gnd_net_),
            .in3(N__36439),
            .lcout(clk_RTD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48395),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.bit_cnt_3789__i3_LC_12_4_0 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3789__i3_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3789__i3_LC_12_4_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \RTD.bit_cnt_3789__i3_LC_12_4_0  (
            .in0(N__35065),
            .in1(N__35117),
            .in2(N__35101),
            .in3(N__35083),
            .lcout(\RTD.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34886),
            .ce(N__34864),
            .sr(N__34852));
    defparam \RTD.bit_cnt_3789__i2_LC_12_4_1 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3789__i2_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3789__i2_LC_12_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RTD.bit_cnt_3789__i2_LC_12_4_1  (
            .in0(N__35082),
            .in1(N__35097),
            .in2(_gnd_net_),
            .in3(N__35064),
            .lcout(\RTD.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34886),
            .ce(N__34864),
            .sr(N__34852));
    defparam \RTD.bit_cnt_3789__i1_LC_12_4_2 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3789__i1_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3789__i1_LC_12_4_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \RTD.bit_cnt_3789__i1_LC_12_4_2  (
            .in0(N__35063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35081),
            .lcout(\RTD.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34886),
            .ce(N__34864),
            .sr(N__34852));
    defparam \RTD.bit_cnt_3789__i0_LC_12_4_7 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3789__i0_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3789__i0_LC_12_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \RTD.bit_cnt_3789__i0_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35062),
            .lcout(\RTD.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34886),
            .ce(N__34864),
            .sr(N__34852));
    defparam clk_cnt_3781_3782__i2_LC_12_5_0.C_ON=1'b0;
    defparam clk_cnt_3781_3782__i2_LC_12_5_0.SEQ_MODE=4'b1000;
    defparam clk_cnt_3781_3782__i2_LC_12_5_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 clk_cnt_3781_3782__i2_LC_12_5_0 (
            .in0(N__36437),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36458),
            .lcout(clk_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48396),
            .ce(),
            .sr(N__36415));
    defparam clk_cnt_3781_3782__i1_LC_12_5_1.C_ON=1'b0;
    defparam clk_cnt_3781_3782__i1_LC_12_5_1.SEQ_MODE=4'b1000;
    defparam clk_cnt_3781_3782__i1_LC_12_5_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 clk_cnt_3781_3782__i1_LC_12_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36436),
            .lcout(clk_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48396),
            .ce(),
            .sr(N__36415));
    defparam comm_cmd_0__bdd_4_lut_20518_LC_12_6_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20518_LC_12_6_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20518_LC_12_6_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_20518_LC_12_6_0 (
            .in0(N__35344),
            .in1(N__60590),
            .in2(N__35311),
            .in3(N__59397),
            .lcout(n23432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_257_LC_12_6_1.C_ON=1'b0;
    defparam i1_4_lut_adj_257_LC_12_6_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_257_LC_12_6_1.LUT_INIT=16'b1010101100000000;
    LogicCell40 i1_4_lut_adj_257_LC_12_6_1 (
            .in0(N__57740),
            .in1(N__51396),
            .in2(N__42781),
            .in3(N__63649),
            .lcout(n12610),
            .ltout(n12610_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i5_LC_12_6_2.C_ON=1'b0;
    defparam buf_control_i5_LC_12_6_2.SEQ_MODE=4'b1000;
    defparam buf_control_i5_LC_12_6_2.LUT_INIT=16'b0010111100100000;
    LogicCell40 buf_control_i5_LC_12_6_2 (
            .in0(N__45312),
            .in1(N__57741),
            .in2(N__35275),
            .in3(N__36500),
            .lcout(AMPV_POW),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61826),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_2_lut_LC_12_6_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_2_lut_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_2_lut_LC_12_6_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_2_lut_LC_12_6_3  (
            .in0(N__57137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43277),
            .lcout(\comm_spi.data_tx_7__N_883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12608_3_lut_LC_12_6_6 .C_ON=1'b0;
    defparam \comm_spi.i12608_3_lut_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12608_3_lut_LC_12_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.i12608_3_lut_LC_12_6_6  (
            .in0(N__41981),
            .in1(N__37492),
            .in2(_gnd_net_),
            .in3(N__41935),
            .lcout(ICE_SPI_MISO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_308_LC_12_7_4.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_308_LC_12_7_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_308_LC_12_7_4.LUT_INIT=16'b1100100011001100;
    LogicCell40 i1_3_lut_4_lut_adj_308_LC_12_7_4 (
            .in0(N__64065),
            .in1(N__63648),
            .in2(N__62677),
            .in3(N__63047),
            .lcout(n13117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_12_7_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_12_7_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_102_2_lut_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__45653),
            .in2(_gnd_net_),
            .in3(N__57109),
            .lcout(\comm_spi.data_tx_7__N_868 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_2_i19_3_lut_LC_12_8_0.C_ON=1'b0;
    defparam mux_127_Mux_2_i19_3_lut_LC_12_8_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_2_i19_3_lut_LC_12_8_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_2_i19_3_lut_LC_12_8_0 (
            .in0(N__35221),
            .in1(N__35447),
            .in2(_gnd_net_),
            .in3(N__59181),
            .lcout(),
            .ltout(n19_adj_1706_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_2_i22_3_lut_LC_12_8_1.C_ON=1'b0;
    defparam mux_127_Mux_2_i22_3_lut_LC_12_8_1.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_2_i22_3_lut_LC_12_8_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_127_Mux_2_i22_3_lut_LC_12_8_1 (
            .in0(_gnd_net_),
            .in1(N__36056),
            .in2(N__36130),
            .in3(N__60007),
            .lcout(n22_adj_1707),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i0_LC_12_8_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i0_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i0_LC_12_8_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i0_LC_12_8_2  (
            .in0(N__35623),
            .in1(N__35929),
            .in2(N__36127),
            .in3(N__37878),
            .lcout(buf_adcdata_vac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61828),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i1_LC_12_8_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i1_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i1_LC_12_8_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i1_LC_12_8_3  (
            .in0(N__39419),
            .in1(N__39812),
            .in2(N__36093),
            .in3(N__35433),
            .lcout(buf_adcdata_iac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61828),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i2_LC_12_8_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i2_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i2_LC_12_8_4 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i2_LC_12_8_4  (
            .in0(N__36057),
            .in1(N__35409),
            .in2(N__39820),
            .in3(N__39420),
            .lcout(buf_adcdata_iac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61828),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i2_LC_12_8_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i2_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i2_LC_12_8_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i2_LC_12_8_5  (
            .in0(N__35448),
            .in1(N__36033),
            .in2(N__35989),
            .in3(N__35624),
            .lcout(buf_adcdata_vac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61828),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_12_8_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_12_8_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i10_LC_12_8_6  (
            .in0(N__39811),
            .in1(N__35405),
            .in2(N__35434),
            .in3(N__37839),
            .lcout(cmd_rdadctmp_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61828),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_12_8_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_12_8_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i11_LC_12_8_7  (
            .in0(N__37838),
            .in1(N__35378),
            .in2(N__35410),
            .in3(N__39816),
            .lcout(cmd_rdadctmp_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61828),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_9_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_9_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_96_2_lut_LC_12_9_0  (
            .in0(N__57172),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46071),
            .lcout(\comm_spi.data_tx_7__N_858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20228_4_lut_3_lut_LC_12_9_1 .C_ON=1'b0;
    defparam \comm_spi.i20228_4_lut_3_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20228_4_lut_3_lut_LC_12_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i20228_4_lut_3_lut_LC_12_9_1  (
            .in0(N__51114),
            .in1(N__40855),
            .in2(_gnd_net_),
            .in3(N__57174),
            .lcout(\comm_spi.n24034 ),
            .ltout(\comm_spi.n24034_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_12628_12629_set_LC_12_9_2 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12628_12629_set_LC_12_9_2 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i3_12628_12629_set_LC_12_9_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.data_tx_i3_12628_12629_set_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__51093),
            .in2(N__36241),
            .in3(N__51075),
            .lcout(\comm_spi.n15356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53627),
            .ce(),
            .sr(N__36214));
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_12_9_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_12_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_97_2_lut_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__40854),
            .in2(_gnd_net_),
            .in3(N__57173),
            .lcout(\comm_spi.data_tx_7__N_859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_12_9_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_12_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_93_2_lut_LC_12_9_5  (
            .in0(N__36201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57170),
            .lcout(\comm_spi.data_tx_7__N_855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20248_4_lut_3_lut_LC_12_9_6 .C_ON=1'b0;
    defparam \comm_spi.i20248_4_lut_3_lut_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20248_4_lut_3_lut_LC_12_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i20248_4_lut_3_lut_LC_12_9_6  (
            .in0(N__57175),
            .in1(N__36202),
            .in2(_gnd_net_),
            .in3(N__36168),
            .lcout(\comm_spi.n24013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_12_9_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_12_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_94_2_lut_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__45658),
            .in2(_gnd_net_),
            .in3(N__57171),
            .lcout(\comm_spi.data_tx_7__N_856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_4_i2_3_lut_LC_12_10_0.C_ON=1'b0;
    defparam mux_134_Mux_4_i2_3_lut_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_4_i2_3_lut_LC_12_10_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_134_Mux_4_i2_3_lut_LC_12_10_0 (
            .in0(N__36834),
            .in1(N__40699),
            .in2(_gnd_net_),
            .in3(N__54416),
            .lcout(),
            .ltout(n2_adj_1669_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i4_LC_12_10_1.C_ON=1'b0;
    defparam comm_tx_buf_i4_LC_12_10_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i4_LC_12_10_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 comm_tx_buf_i4_LC_12_10_1 (
            .in0(N__36310),
            .in1(N__36136),
            .in2(N__36142),
            .in3(N__54613),
            .lcout(comm_tx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61833),
            .ce(N__46427),
            .sr(N__46350));
    defparam mux_134_Mux_4_i4_3_lut_LC_12_10_2.C_ON=1'b0;
    defparam mux_134_Mux_4_i4_3_lut_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_4_i4_3_lut_LC_12_10_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_134_Mux_4_i4_3_lut_LC_12_10_2 (
            .in0(N__43084),
            .in1(N__54979),
            .in2(_gnd_net_),
            .in3(N__54415),
            .lcout(),
            .ltout(n4_adj_1670_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_20463_LC_12_10_3.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_20463_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_20463_LC_12_10_3.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_index_1__bdd_4_lut_20463_LC_12_10_3 (
            .in0(N__36316),
            .in1(N__54612),
            .in2(N__36139),
            .in3(N__51838),
            .lcout(n23402),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20124_2_lut_LC_12_10_4.C_ON=1'b0;
    defparam i20124_2_lut_LC_12_10_4.SEQ_MODE=4'b0000;
    defparam i20124_2_lut_LC_12_10_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 i20124_2_lut_LC_12_10_4 (
            .in0(_gnd_net_),
            .in1(N__38139),
            .in2(_gnd_net_),
            .in3(N__54413),
            .lcout(n22669),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_4_i1_3_lut_LC_12_10_5.C_ON=1'b0;
    defparam mux_134_Mux_4_i1_3_lut_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_4_i1_3_lut_LC_12_10_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_134_Mux_4_i1_3_lut_LC_12_10_5 (
            .in0(N__54414),
            .in1(_gnd_net_),
            .in2(N__44693),
            .in3(N__56096),
            .lcout(n1_adj_1668),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10493_3_lut_LC_12_10_6.C_ON=1'b0;
    defparam i10493_3_lut_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam i10493_3_lut_LC_12_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i10493_3_lut_LC_12_10_6 (
            .in0(N__36833),
            .in1(N__44677),
            .in2(_gnd_net_),
            .in3(N__46164),
            .lcout(n13219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_12_10_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_12_10_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_103_2_lut_LC_12_10_7  (
            .in0(N__57176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36285),
            .lcout(\comm_spi.data_tx_7__N_871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i0_LC_12_11_0.C_ON=1'b0;
    defparam comm_buf_0__i0_LC_12_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i0_LC_12_11_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_0__i0_LC_12_11_0 (
            .in0(N__62657),
            .in1(N__54024),
            .in2(_gnd_net_),
            .in3(N__38377),
            .lcout(comm_buf_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61839),
            .ce(N__61438),
            .sr(N__64417));
    defparam comm_buf_0__i1_LC_12_11_1.C_ON=1'b0;
    defparam comm_buf_0__i1_LC_12_11_1.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i1_LC_12_11_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i1_LC_12_11_1 (
            .in0(N__54809),
            .in1(N__62660),
            .in2(_gnd_net_),
            .in3(N__43555),
            .lcout(comm_buf_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61839),
            .ce(N__61438),
            .sr(N__64417));
    defparam comm_buf_0__i2_LC_12_11_2.C_ON=1'b0;
    defparam comm_buf_0__i2_LC_12_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i2_LC_12_11_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_0__i2_LC_12_11_2 (
            .in0(N__54939),
            .in1(_gnd_net_),
            .in2(N__38488),
            .in3(N__62663),
            .lcout(comm_buf_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61839),
            .ce(N__61438),
            .sr(N__64417));
    defparam comm_buf_0__i4_LC_12_11_3.C_ON=1'b0;
    defparam comm_buf_0__i4_LC_12_11_3.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i4_LC_12_11_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i4_LC_12_11_3 (
            .in0(N__55071),
            .in1(N__62661),
            .in2(_gnd_net_),
            .in3(N__36262),
            .lcout(comm_buf_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61839),
            .ce(N__61438),
            .sr(N__64417));
    defparam comm_buf_0__i5_LC_12_11_4.C_ON=1'b0;
    defparam comm_buf_0__i5_LC_12_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i5_LC_12_11_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_0__i5_LC_12_11_4 (
            .in0(N__62658),
            .in1(N__55206),
            .in2(_gnd_net_),
            .in3(N__57919),
            .lcout(comm_buf_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61839),
            .ce(N__61438),
            .sr(N__64417));
    defparam comm_buf_0__i6_LC_12_11_5.C_ON=1'b0;
    defparam comm_buf_0__i6_LC_12_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i6_LC_12_11_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i6_LC_12_11_5 (
            .in0(N__53895),
            .in1(N__62662),
            .in2(_gnd_net_),
            .in3(N__36253),
            .lcout(comm_buf_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61839),
            .ce(N__61438),
            .sr(N__64417));
    defparam comm_buf_0__i7_LC_12_11_6.C_ON=1'b0;
    defparam comm_buf_0__i7_LC_12_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i7_LC_12_11_6.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_0__i7_LC_12_11_6 (
            .in0(N__62659),
            .in1(N__55937),
            .in2(N__36481),
            .in3(_gnd_net_),
            .lcout(comm_buf_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61839),
            .ce(N__61438),
            .sr(N__64417));
    defparam i16298_2_lut_LC_12_11_7.C_ON=1'b0;
    defparam i16298_2_lut_LC_12_11_7.SEQ_MODE=4'b0000;
    defparam i16298_2_lut_LC_12_11_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i16298_2_lut_LC_12_11_7 (
            .in0(N__36466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36438),
            .lcout(n18996),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i0_LC_12_12_0.C_ON=1'b0;
    defparam comm_buf_2__i0_LC_12_12_0.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i0_LC_12_12_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_2__i0_LC_12_12_0 (
            .in0(N__36400),
            .in1(N__62620),
            .in2(_gnd_net_),
            .in3(N__54025),
            .lcout(comm_buf_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam comm_buf_2__i1_LC_12_12_1.C_ON=1'b0;
    defparam comm_buf_2__i1_LC_12_12_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i1_LC_12_12_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_2__i1_LC_12_12_1 (
            .in0(N__62616),
            .in1(_gnd_net_),
            .in2(N__36394),
            .in3(N__54800),
            .lcout(comm_buf_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam comm_buf_2__i2_LC_12_12_2.C_ON=1'b0;
    defparam comm_buf_2__i2_LC_12_12_2.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i2_LC_12_12_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_2__i2_LC_12_12_2 (
            .in0(N__41047),
            .in1(N__54940),
            .in2(_gnd_net_),
            .in3(N__62621),
            .lcout(comm_buf_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam comm_buf_2__i3_LC_12_12_3.C_ON=1'b0;
    defparam comm_buf_2__i3_LC_12_12_3.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i3_LC_12_12_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i3_LC_12_12_3 (
            .in0(N__62617),
            .in1(N__62789),
            .in2(_gnd_net_),
            .in3(N__36382),
            .lcout(comm_buf_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam comm_buf_2__i4_LC_12_12_4.C_ON=1'b0;
    defparam comm_buf_2__i4_LC_12_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i4_LC_12_12_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i4_LC_12_12_4 (
            .in0(N__55072),
            .in1(N__36373),
            .in2(_gnd_net_),
            .in3(N__62622),
            .lcout(comm_buf_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam comm_buf_2__i5_LC_12_12_5.C_ON=1'b0;
    defparam comm_buf_2__i5_LC_12_12_5.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i5_LC_12_12_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i5_LC_12_12_5 (
            .in0(N__62618),
            .in1(N__55207),
            .in2(_gnd_net_),
            .in3(N__36364),
            .lcout(comm_buf_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam comm_buf_2__i6_LC_12_12_6.C_ON=1'b0;
    defparam comm_buf_2__i6_LC_12_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i6_LC_12_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i6_LC_12_12_6 (
            .in0(N__53896),
            .in1(N__36355),
            .in2(_gnd_net_),
            .in3(N__62623),
            .lcout(comm_buf_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam comm_buf_2__i7_LC_12_12_7.C_ON=1'b0;
    defparam comm_buf_2__i7_LC_12_12_7.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i7_LC_12_12_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_2__i7_LC_12_12_7 (
            .in0(N__62619),
            .in1(_gnd_net_),
            .in2(N__55945),
            .in3(N__36727),
            .lcout(comm_buf_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61844),
            .ce(N__43462),
            .sr(N__38425));
    defparam \comm_spi.data_tx_i2_12624_12625_set_LC_12_13_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12624_12625_set_LC_12_13_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i2_12624_12625_set_LC_12_13_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \comm_spi.data_tx_i2_12624_12625_set_LC_12_13_0  (
            .in0(N__37519),
            .in1(_gnd_net_),
            .in2(N__37573),
            .in3(N__37540),
            .lcout(\comm_spi.n15352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53697),
            .ce(),
            .sr(N__36715));
    defparam i4032_2_lut_3_lut_LC_12_13_3.C_ON=1'b0;
    defparam i4032_2_lut_3_lut_LC_12_13_3.SEQ_MODE=4'b0000;
    defparam i4032_2_lut_3_lut_LC_12_13_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 i4032_2_lut_3_lut_LC_12_13_3 (
            .in0(N__41019),
            .in1(N__38583),
            .in2(_gnd_net_),
            .in3(N__59367),
            .lcout(n6774),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i45_3_lut_LC_12_13_4.C_ON=1'b0;
    defparam i45_3_lut_LC_12_13_4.SEQ_MODE=4'b0000;
    defparam i45_3_lut_LC_12_13_4.LUT_INIT=16'b0011001111101110;
    LogicCell40 i45_3_lut_LC_12_13_4 (
            .in0(N__59364),
            .in1(N__61382),
            .in2(_gnd_net_),
            .in3(N__58652),
            .lcout(n40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_2_i111_3_lut_LC_12_13_5.C_ON=1'b0;
    defparam mux_125_Mux_2_i111_3_lut_LC_12_13_5.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_2_i111_3_lut_LC_12_13_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_2_i111_3_lut_LC_12_13_5 (
            .in0(N__38371),
            .in1(N__36630),
            .in2(_gnd_net_),
            .in3(N__59365),
            .lcout(),
            .ltout(n111_adj_1796_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_2_i112_3_lut_LC_12_13_6.C_ON=1'b0;
    defparam mux_125_Mux_2_i112_3_lut_LC_12_13_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_2_i112_3_lut_LC_12_13_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_125_Mux_2_i112_3_lut_LC_12_13_6 (
            .in0(_gnd_net_),
            .in1(N__41066),
            .in2(N__36634),
            .in3(N__60597),
            .lcout(n112_adj_1797),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_2_i111_3_lut_LC_12_13_7.C_ON=1'b0;
    defparam mux_126_Mux_2_i111_3_lut_LC_12_13_7.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_2_i111_3_lut_LC_12_13_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_126_Mux_2_i111_3_lut_LC_12_13_7 (
            .in0(N__41067),
            .in1(N__36631),
            .in2(_gnd_net_),
            .in3(N__59366),
            .lcout(n111_adj_1750),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_12640_12641_set_LC_12_14_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12640_12641_set_LC_12_14_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i6_12640_12641_set_LC_12_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.data_tx_i6_12640_12641_set_LC_12_14_0  (
            .in0(N__36622),
            .in1(N__36598),
            .in2(_gnd_net_),
            .in3(N__36574),
            .lcout(\comm_spi.n15368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53698),
            .ce(),
            .sr(N__36529));
    defparam mux_125_Mux_5_i23_3_lut_LC_12_14_1.C_ON=1'b0;
    defparam mux_125_Mux_5_i23_3_lut_LC_12_14_1.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_5_i23_3_lut_LC_12_14_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_125_Mux_5_i23_3_lut_LC_12_14_1 (
            .in0(N__36501),
            .in1(N__59351),
            .in2(_gnd_net_),
            .in3(N__38821),
            .lcout(n23_adj_1773),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_7_i111_3_lut_LC_12_14_2.C_ON=1'b0;
    defparam mux_125_Mux_7_i111_3_lut_LC_12_14_2.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_7_i111_3_lut_LC_12_14_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_125_Mux_7_i111_3_lut_LC_12_14_2 (
            .in0(N__59353),
            .in1(N__42376),
            .in2(_gnd_net_),
            .in3(N__38322),
            .lcout(n111_adj_1761),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_1_i111_3_lut_LC_12_14_5.C_ON=1'b0;
    defparam mux_126_Mux_1_i111_3_lut_LC_12_14_5.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_1_i111_3_lut_LC_12_14_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_126_Mux_1_i111_3_lut_LC_12_14_5 (
            .in0(N__41871),
            .in1(N__38391),
            .in2(_gnd_net_),
            .in3(N__59355),
            .lcout(n111_adj_1754),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_3_i16_3_lut_LC_12_14_6.C_ON=1'b0;
    defparam mux_126_Mux_3_i16_3_lut_LC_12_14_6.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_3_i16_3_lut_LC_12_14_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_126_Mux_3_i16_3_lut_LC_12_14_6 (
            .in0(N__59352),
            .in1(N__36867),
            .in2(_gnd_net_),
            .in3(N__40069),
            .lcout(n16_adj_1738),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_4_i16_3_lut_LC_12_14_7.C_ON=1'b0;
    defparam mux_126_Mux_4_i16_3_lut_LC_12_14_7.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_4_i16_3_lut_LC_12_14_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_4_i16_3_lut_LC_12_14_7 (
            .in0(N__49458),
            .in1(N__47268),
            .in2(_gnd_net_),
            .in3(N__59354),
            .lcout(n16_adj_1733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_51_LC_12_15_0.C_ON=1'b0;
    defparam i1_4_lut_adj_51_LC_12_15_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_51_LC_12_15_0.LUT_INIT=16'b1010100000100000;
    LogicCell40 i1_4_lut_adj_51_LC_12_15_0 (
            .in0(N__37393),
            .in1(N__59446),
            .in2(N__56078),
            .in3(N__36841),
            .lcout(),
            .ltout(n11987_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i5_LC_12_15_1.C_ON=1'b0;
    defparam buf_device_acadc_i5_LC_12_15_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i5_LC_12_15_1.LUT_INIT=16'b1111111011111100;
    LogicCell40 buf_device_acadc_i5_LC_12_15_1 (
            .in0(N__44714),
            .in1(N__38707),
            .in2(N__36817),
            .in3(N__43612),
            .lcout(VAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61870),
            .ce(N__36794),
            .sr(N__37130));
    defparam mux_125_Mux_4_i17_3_lut_LC_12_15_2.C_ON=1'b0;
    defparam mux_125_Mux_4_i17_3_lut_LC_12_15_2.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i17_3_lut_LC_12_15_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_4_i17_3_lut_LC_12_15_2 (
            .in0(N__37164),
            .in1(N__38792),
            .in2(_gnd_net_),
            .in3(N__59444),
            .lcout(n17_adj_1779),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_258_LC_12_15_3.C_ON=1'b0;
    defparam i1_4_lut_adj_258_LC_12_15_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_258_LC_12_15_3.LUT_INIT=16'b1110010000000000;
    LogicCell40 i1_4_lut_adj_258_LC_12_15_3 (
            .in0(N__59445),
            .in1(N__49146),
            .in2(N__43228),
            .in3(N__37392),
            .lcout(),
            .ltout(n11985_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i1_LC_12_15_4.C_ON=1'b0;
    defparam buf_device_acadc_i1_LC_12_15_4.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i1_LC_12_15_4.LUT_INIT=16'b1111111011111100;
    LogicCell40 buf_device_acadc_i1_LC_12_15_4 (
            .in0(N__43933),
            .in1(N__37060),
            .in2(N__36802),
            .in3(N__43415),
            .lcout(IAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61870),
            .ce(N__36794),
            .sr(N__37130));
    defparam i1_2_lut_4_lut_adj_268_LC_12_15_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_268_LC_12_15_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_268_LC_12_15_5.LUT_INIT=16'b1111101100000000;
    LogicCell40 i1_2_lut_4_lut_adj_268_LC_12_15_5 (
            .in0(N__50890),
            .in1(N__55650),
            .in2(N__38758),
            .in3(N__37079),
            .lcout(n24_adj_1575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_269_LC_12_15_7.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_269_LC_12_15_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_269_LC_12_15_7.LUT_INIT=16'b1111101100000000;
    LogicCell40 i1_2_lut_4_lut_adj_269_LC_12_15_7 (
            .in0(N__50889),
            .in1(N__55649),
            .in2(N__38759),
            .in3(N__37037),
            .lcout(n24_adj_1601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_54_LC_12_16_0.C_ON=1'b0;
    defparam i1_4_lut_adj_54_LC_12_16_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_54_LC_12_16_0.LUT_INIT=16'b1101100000000000;
    LogicCell40 i1_4_lut_adj_54_LC_12_16_0 (
            .in0(N__59363),
            .in1(N__45699),
            .in2(N__56582),
            .in3(N__37381),
            .lcout(n11984),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i9_LC_12_16_1.C_ON=1'b0;
    defparam acadc_skipCount_i9_LC_12_16_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i9_LC_12_16_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 acadc_skipCount_i9_LC_12_16_1 (
            .in0(N__46842),
            .in1(N__50814),
            .in2(_gnd_net_),
            .in3(N__49848),
            .lcout(acadc_skipCount_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61883),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i1_LC_12_16_2.C_ON=1'b0;
    defparam buf_cfgRTD_i1_LC_12_16_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i1_LC_12_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i1_LC_12_16_2 (
            .in0(N__50815),
            .in1(N__48799),
            .in2(_gnd_net_),
            .in3(N__38215),
            .lcout(buf_cfgRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61883),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_330_LC_12_16_3.C_ON=1'b0;
    defparam acadc_rst_330_LC_12_16_3.SEQ_MODE=4'b1000;
    defparam acadc_rst_330_LC_12_16_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_rst_330_LC_12_16_3 (
            .in0(N__40948),
            .in1(N__43872),
            .in2(_gnd_net_),
            .in3(N__39148),
            .lcout(acadc_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61883),
            .ce(),
            .sr(_gnd_net_));
    defparam n23438_bdd_4_lut_LC_12_16_4.C_ON=1'b0;
    defparam n23438_bdd_4_lut_LC_12_16_4.SEQ_MODE=4'b0000;
    defparam n23438_bdd_4_lut_LC_12_16_4.LUT_INIT=16'b1100110011100010;
    LogicCell40 n23438_bdd_4_lut_LC_12_16_4 (
            .in0(N__37006),
            .in1(N__36997),
            .in2(N__36978),
            .in3(N__60072),
            .lcout(n23441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_5_i111_3_lut_LC_12_16_5.C_ON=1'b0;
    defparam mux_125_Mux_5_i111_3_lut_LC_12_16_5.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_5_i111_3_lut_LC_12_16_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_5_i111_3_lut_LC_12_16_5 (
            .in0(N__36951),
            .in1(N__36933),
            .in2(_gnd_net_),
            .in3(N__59362),
            .lcout(),
            .ltout(n111_adj_1776_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_5_i112_3_lut_LC_12_16_6.C_ON=1'b0;
    defparam mux_125_Mux_5_i112_3_lut_LC_12_16_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_5_i112_3_lut_LC_12_16_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_125_Mux_5_i112_3_lut_LC_12_16_6 (
            .in0(_gnd_net_),
            .in1(N__36914),
            .in2(N__36883),
            .in3(N__60635),
            .lcout(n112_adj_1777),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_59_LC_12_16_7.C_ON=1'b0;
    defparam i2_3_lut_adj_59_LC_12_16_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_59_LC_12_16_7.LUT_INIT=16'b0000101000000000;
    LogicCell40 i2_3_lut_adj_59_LC_12_16_7 (
            .in0(N__60636),
            .in1(_gnd_net_),
            .in2(N__60097),
            .in3(N__41020),
            .lcout(n11979),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i11_LC_12_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i11_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i11_LC_12_17_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i11_LC_12_17_0  (
            .in0(N__39400),
            .in1(N__39799),
            .in2(N__44228),
            .in3(N__37284),
            .lcout(buf_adcdata_iac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61895),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_12_17_1.C_ON=1'b0;
    defparam i8_4_lut_LC_12_17_1.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_12_17_1.LUT_INIT=16'b0111101111011110;
    LogicCell40 i8_4_lut_LC_12_17_1 (
            .in0(N__37351),
            .in1(N__37333),
            .in2(N__41511),
            .in3(N__49844),
            .lcout(n24_adj_1513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_233_LC_12_17_2.C_ON=1'b0;
    defparam i7_4_lut_adj_233_LC_12_17_2.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_233_LC_12_17_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i7_4_lut_adj_233_LC_12_17_2 (
            .in0(N__37315),
            .in1(N__37300),
            .in2(N__52743),
            .in3(N__37475),
            .lcout(n23_adj_1514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_12_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_12_17_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i20_LC_12_17_3  (
            .in0(N__39798),
            .in1(N__37244),
            .in2(N__37285),
            .in3(N__37796),
            .lcout(cmd_rdadctmp_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61895),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i14_LC_12_17_4.C_ON=1'b0;
    defparam acadc_skipCount_i14_LC_12_17_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i14_LC_12_17_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i14_LC_12_17_4 (
            .in0(N__57848),
            .in1(N__46852),
            .in2(N__40569),
            .in3(N__37476),
            .lcout(acadc_skipCount_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61895),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_0_i16_3_lut_LC_12_17_5.C_ON=1'b0;
    defparam mux_126_Mux_0_i16_3_lut_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_0_i16_3_lut_LC_12_17_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 mux_126_Mux_0_i16_3_lut_LC_12_17_5 (
            .in0(N__37227),
            .in1(_gnd_net_),
            .in2(N__59513),
            .in3(N__47232),
            .lcout(n16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i20_LC_12_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i20_LC_12_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i20_LC_12_17_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i20_LC_12_17_7  (
            .in0(N__39797),
            .in1(N__39401),
            .in2(N__37198),
            .in3(N__37163),
            .lcout(buf_adcdata_iac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61895),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i10_LC_12_18_1.C_ON=1'b0;
    defparam acadc_skipCount_i10_LC_12_18_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i10_LC_12_18_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_skipCount_i10_LC_12_18_1 (
            .in0(N__47454),
            .in1(N__46846),
            .in2(_gnd_net_),
            .in3(N__39910),
            .lcout(acadc_skipCount_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61910),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i15_LC_12_18_2.C_ON=1'b0;
    defparam acadc_skipCount_i15_LC_12_18_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i15_LC_12_18_2.LUT_INIT=16'b0111001001010000;
    LogicCell40 acadc_skipCount_i15_LC_12_18_2 (
            .in0(N__46845),
            .in1(N__57850),
            .in2(N__41510),
            .in3(N__46646),
            .lcout(acadc_skipCount_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61910),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i6_LC_12_18_3.C_ON=1'b0;
    defparam buf_control_i6_LC_12_18_3.SEQ_MODE=4'b1000;
    defparam buf_control_i6_LC_12_18_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i6_LC_12_18_3 (
            .in0(N__57849),
            .in1(N__46738),
            .in2(N__40568),
            .in3(N__37486),
            .lcout(buf_control_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61910),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i2_LC_12_18_4.C_ON=1'b0;
    defparam buf_control_i2_LC_12_18_4.SEQ_MODE=4'b1000;
    defparam buf_control_i2_LC_12_18_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 buf_control_i2_LC_12_18_4 (
            .in0(N__46736),
            .in1(N__47455),
            .in2(_gnd_net_),
            .in3(N__39927),
            .lcout(SELIRNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61910),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_6_i23_3_lut_LC_12_18_6.C_ON=1'b0;
    defparam mux_125_Mux_6_i23_3_lut_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_6_i23_3_lut_LC_12_18_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_125_Mux_6_i23_3_lut_LC_12_18_6 (
            .in0(N__37485),
            .in1(N__59479),
            .in2(_gnd_net_),
            .in3(N__37477),
            .lcout(n23_adj_1767),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i4_LC_12_18_7.C_ON=1'b0;
    defparam buf_control_i4_LC_12_18_7.SEQ_MODE=4'b1000;
    defparam buf_control_i4_LC_12_18_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_control_i4_LC_12_18_7 (
            .in0(N__47356),
            .in1(N__46737),
            .in2(_gnd_net_),
            .in3(N__39875),
            .lcout(VDC_RNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61910),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i1_LC_12_19_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i1_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i1_LC_12_19_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i1_LC_12_19_0  (
            .in0(N__50540),
            .in1(N__50374),
            .in2(N__37447),
            .in3(N__42153),
            .lcout(\SIG_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61929),
            .ce(N__42205),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i0_LC_12_19_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i0_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i0_LC_12_19_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i0_LC_12_19_2  (
            .in0(N__50539),
            .in1(N__50373),
            .in2(N__40044),
            .in3(N__47233),
            .lcout(\SIG_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61929),
            .ce(N__42205),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i3_LC_12_19_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i3_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i3_LC_12_19_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i3_LC_12_19_3  (
            .in0(N__50372),
            .in1(N__50542),
            .in2(N__37414),
            .in3(N__40065),
            .lcout(\SIG_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61929),
            .ce(N__42205),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i2_LC_12_19_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i2_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i2_LC_12_19_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i2_LC_12_19_6  (
            .in0(N__50541),
            .in1(N__50375),
            .in2(N__37423),
            .in3(N__42358),
            .lcout(\SIG_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61929),
            .ce(N__42205),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i1_12620_12621_reset_LC_13_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12620_12621_reset_LC_13_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i1_12620_12621_reset_LC_13_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12620_12621_reset_LC_13_3_0  (
            .in0(N__37603),
            .in1(N__40288),
            .in2(_gnd_net_),
            .in3(N__37626),
            .lcout(\comm_spi.n15349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53568),
            .ce(),
            .sr(N__37582));
    defparam \comm_spi.data_tx_i1_12620_12621_set_LC_13_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12620_12621_set_LC_13_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i1_12620_12621_set_LC_13_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12620_12621_set_LC_13_4_0  (
            .in0(N__37599),
            .in1(N__40287),
            .in2(_gnd_net_),
            .in3(N__37633),
            .lcout(\comm_spi.n15348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53588),
            .ce(),
            .sr(N__37612));
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_13_4_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_13_4_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_98_2_lut_LC_13_4_2  (
            .in0(N__57115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37941),
            .lcout(\comm_spi.data_tx_7__N_860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_13_4_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_13_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_99_2_lut_LC_13_4_3  (
            .in0(_gnd_net_),
            .in1(N__43285),
            .in2(_gnd_net_),
            .in3(N__57116),
            .lcout(\comm_spi.data_tx_7__N_861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20218_4_lut_3_lut_LC_13_4_4 .C_ON=1'b0;
    defparam \comm_spi.i20218_4_lut_3_lut_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20218_4_lut_3_lut_LC_13_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i20218_4_lut_3_lut_LC_13_4_4  (
            .in0(N__57117),
            .in1(N__37942),
            .in2(_gnd_net_),
            .in3(N__37556),
            .lcout(\comm_spi.n24037 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_20449_LC_13_5_1.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_20449_LC_13_5_1.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_20449_LC_13_5_1.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_1__bdd_4_lut_20449_LC_13_5_1 (
            .in0(N__42520),
            .in1(N__54608),
            .in2(N__37921),
            .in3(N__51823),
            .lcout(n23390),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20253_4_lut_3_lut_LC_13_5_3 .C_ON=1'b0;
    defparam \comm_spi.i20253_4_lut_3_lut_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20253_4_lut_3_lut_LC_13_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i20253_4_lut_3_lut_LC_13_5_3  (
            .in0(N__57114),
            .in1(N__43284),
            .in2(_gnd_net_),
            .in3(N__37598),
            .lcout(\comm_spi.n24040 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_13_5_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_13_5_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \comm_spi.RESET_I_0_106_2_lut_LC_13_5_4  (
            .in0(N__37940),
            .in1(N__57113),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i2_12624_12625_reset_LC_13_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12624_12625_reset_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i2_12624_12625_reset_LC_13_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12624_12625_reset_LC_13_6_0  (
            .in0(N__37563),
            .in1(N__37533),
            .in2(_gnd_net_),
            .in3(N__37509),
            .lcout(\comm_spi.n15353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53601),
            .ce(),
            .sr(N__40834));
    defparam \comm_spi.MISO_48_12606_12607_reset_LC_13_7_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12606_12607_reset_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.MISO_48_12606_12607_reset_LC_13_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.MISO_48_12606_12607_reset_LC_13_7_0  (
            .in0(N__41970),
            .in1(N__42021),
            .in2(_gnd_net_),
            .in3(N__42003),
            .lcout(\comm_spi.n15335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12606_12607_resetC_net ),
            .ce(),
            .sr(N__40619));
    defparam mux_134_Mux_1_i1_3_lut_LC_13_8_0.C_ON=1'b0;
    defparam mux_134_Mux_1_i1_3_lut_LC_13_8_0.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_1_i1_3_lut_LC_13_8_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_134_Mux_1_i1_3_lut_LC_13_8_0 (
            .in0(N__52121),
            .in1(N__44592),
            .in2(_gnd_net_),
            .in3(N__54372),
            .lcout(),
            .ltout(n1_adj_1674_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i1_LC_13_8_1.C_ON=1'b0;
    defparam comm_tx_buf_i1_LC_13_8_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i1_LC_13_8_1.LUT_INIT=16'b1100110010111000;
    LogicCell40 comm_tx_buf_i1_LC_13_8_1 (
            .in0(N__37909),
            .in1(N__37957),
            .in2(N__37945),
            .in3(N__54584),
            .lcout(comm_tx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61831),
            .ce(N__46402),
            .sr(N__46354));
    defparam i19782_2_lut_LC_13_8_2.C_ON=1'b0;
    defparam i19782_2_lut_LC_13_8_2.SEQ_MODE=4'b0000;
    defparam i19782_2_lut_LC_13_8_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19782_2_lut_LC_13_8_2 (
            .in0(_gnd_net_),
            .in1(N__40461),
            .in2(_gnd_net_),
            .in3(N__54370),
            .lcout(n22341),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_1_i2_3_lut_LC_13_8_4.C_ON=1'b0;
    defparam mux_134_Mux_1_i2_3_lut_LC_13_8_4.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_1_i2_3_lut_LC_13_8_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_134_Mux_1_i2_3_lut_LC_13_8_4 (
            .in0(N__41107),
            .in1(N__38307),
            .in2(_gnd_net_),
            .in3(N__54371),
            .lcout(n2_adj_1675),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_0_i19_3_lut_LC_13_9_2.C_ON=1'b0;
    defparam mux_127_Mux_0_i19_3_lut_LC_13_9_2.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_0_i19_3_lut_LC_13_9_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_0_i19_3_lut_LC_13_9_2 (
            .in0(N__37903),
            .in1(N__37874),
            .in2(_gnd_net_),
            .in3(N__59436),
            .lcout(),
            .ltout(n19_adj_1590_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_0_i22_3_lut_LC_13_9_3.C_ON=1'b0;
    defparam mux_127_Mux_0_i22_3_lut_LC_13_9_3.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_0_i22_3_lut_LC_13_9_3.LUT_INIT=16'b1110001011100010;
    LogicCell40 mux_127_Mux_0_i22_3_lut_LC_13_9_3 (
            .in0(N__38087),
            .in1(N__59993),
            .in2(N__37858),
            .in3(_gnd_net_),
            .lcout(n22_adj_1589),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_13_9_4.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_13_9_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_13_9_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_4_lut_LC_13_9_4 (
            .in0(N__59994),
            .in1(N__60467),
            .in2(N__46534),
            .in3(N__59437),
            .lcout(n21965),
            .ltout(n21965_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_295_LC_13_9_5.C_ON=1'b0;
    defparam i1_3_lut_adj_295_LC_13_9_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_295_LC_13_9_5.LUT_INIT=16'b1100111100000000;
    LogicCell40 i1_3_lut_adj_295_LC_13_9_5 (
            .in0(_gnd_net_),
            .in1(N__57665),
            .in2(N__37843),
            .in3(N__63610),
            .lcout(n13093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_13_9_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_13_9_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i8_LC_13_9_6  (
            .in0(N__37800),
            .in1(N__38117),
            .in2(N__38170),
            .in3(N__39810),
            .lcout(cmd_rdadctmp_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61835),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i4_LC_13_9_7.C_ON=1'b0;
    defparam comm_buf_6__i4_LC_13_9_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i4_LC_13_9_7.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i4_LC_13_9_7 (
            .in0(N__38140),
            .in1(N__63611),
            .in2(N__55076),
            .in3(N__45562),
            .lcout(comm_buf_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61835),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i0_LC_13_10_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i0_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i0_LC_13_10_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i0_LC_13_10_0  (
            .in0(N__39405),
            .in1(N__39758),
            .in2(N__38097),
            .in3(N__38118),
            .lcout(buf_adcdata_iac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61841),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_5_i19_3_lut_LC_13_10_1.C_ON=1'b0;
    defparam mux_126_Mux_5_i19_3_lut_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_5_i19_3_lut_LC_13_10_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_5_i19_3_lut_LC_13_10_1 (
            .in0(N__38071),
            .in1(N__38043),
            .in2(_gnd_net_),
            .in3(N__59435),
            .lcout(),
            .ltout(n19_adj_1729_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20424_LC_13_10_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20424_LC_13_10_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20424_LC_13_10_2.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20424_LC_13_10_2 (
            .in0(N__38017),
            .in1(N__59991),
            .in2(N__37993),
            .in3(N__60668),
            .lcout(n23354),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i6_LC_13_10_3.C_ON=1'b0;
    defparam comm_buf_6__i6_LC_13_10_3.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i6_LC_13_10_3.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i6_LC_13_10_3 (
            .in0(N__37989),
            .in1(N__63612),
            .in2(N__53894),
            .in3(N__45569),
            .lcout(comm_buf_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61841),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_3_lut_LC_13_10_4.C_ON=1'b0;
    defparam i3_2_lut_3_lut_LC_13_10_4.SEQ_MODE=4'b0000;
    defparam i3_2_lut_3_lut_LC_13_10_4.LUT_INIT=16'b0011001100100010;
    LogicCell40 i3_2_lut_3_lut_LC_13_10_4 (
            .in0(N__59432),
            .in1(N__59992),
            .in2(_gnd_net_),
            .in3(N__60666),
            .lcout(n9_adj_1600),
            .ltout(n9_adj_1600_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4034_2_lut_3_lut_4_lut_LC_13_10_5.C_ON=1'b0;
    defparam i4034_2_lut_3_lut_4_lut_LC_13_10_5.SEQ_MODE=4'b0000;
    defparam i4034_2_lut_3_lut_4_lut_LC_13_10_5.LUT_INIT=16'b1000000011000000;
    LogicCell40 i4034_2_lut_3_lut_4_lut_LC_13_10_5 (
            .in0(N__60667),
            .in1(N__41005),
            .in2(N__37975),
            .in3(N__59433),
            .lcout(n6776),
            .ltout(n6776_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16190_3_lut_LC_13_10_6.C_ON=1'b0;
    defparam i16190_3_lut_LC_13_10_6.SEQ_MODE=4'b0000;
    defparam i16190_3_lut_LC_13_10_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 i16190_3_lut_LC_13_10_6 (
            .in0(N__45695),
            .in1(_gnd_net_),
            .in2(N__37972),
            .in3(N__45283),
            .lcout(n18890),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_1_i111_3_lut_LC_13_10_7.C_ON=1'b0;
    defparam mux_125_Mux_1_i111_3_lut_LC_13_10_7.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_1_i111_3_lut_LC_13_10_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_1_i111_3_lut_LC_13_10_7 (
            .in0(N__43060),
            .in1(N__38395),
            .in2(_gnd_net_),
            .in3(N__59434),
            .lcout(n111_adj_1798),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_0_i127_3_lut_LC_13_11_0.C_ON=1'b0;
    defparam mux_125_Mux_0_i127_3_lut_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_0_i127_3_lut_LC_13_11_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_125_Mux_0_i127_3_lut_LC_13_11_0 (
            .in0(N__38521),
            .in1(N__61254),
            .in2(_gnd_net_),
            .in3(N__38530),
            .lcout(comm_buf_0_7_N_543_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i16_LC_13_11_1.C_ON=1'b0;
    defparam comm_test_buf_24_i16_LC_13_11_1.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i16_LC_13_11_1.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_test_buf_24_i16_LC_13_11_1 (
            .in0(N__57878),
            .in1(N__38472),
            .in2(N__43940),
            .in3(N__45401),
            .lcout(comm_test_buf_24_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61847),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i18_LC_13_11_2.C_ON=1'b0;
    defparam comm_test_buf_24_i18_LC_13_11_2.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i18_LC_13_11_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_test_buf_24_i18_LC_13_11_2 (
            .in0(N__45400),
            .in1(N__57879),
            .in2(N__40924),
            .in3(N__38367),
            .lcout(comm_test_buf_24_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61847),
            .ce(),
            .sr(_gnd_net_));
    defparam i16302_2_lut_LC_13_11_3.C_ON=1'b0;
    defparam i16302_2_lut_LC_13_11_3.SEQ_MODE=4'b0000;
    defparam i16302_2_lut_LC_13_11_3.LUT_INIT=16'b1111111100110011;
    LogicCell40 i16302_2_lut_LC_13_11_3 (
            .in0(_gnd_net_),
            .in1(N__60269),
            .in2(_gnd_net_),
            .in3(N__58855),
            .lcout(n112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_7_i111_3_lut_LC_13_11_4.C_ON=1'b0;
    defparam mux_126_Mux_7_i111_3_lut_LC_13_11_4.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_7_i111_3_lut_LC_13_11_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_126_Mux_7_i111_3_lut_LC_13_11_4 (
            .in0(N__58857),
            .in1(N__38353),
            .in2(_gnd_net_),
            .in3(N__38329),
            .lcout(n111_adj_1719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10475_3_lut_LC_13_11_5.C_ON=1'b0;
    defparam i10475_3_lut_LC_13_11_5.SEQ_MODE=4'b0000;
    defparam i10475_3_lut_LC_13_11_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i10475_3_lut_LC_13_11_5 (
            .in0(N__38297),
            .in1(N__44565),
            .in2(_gnd_net_),
            .in3(N__46195),
            .lcout(n13201),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_20538_LC_13_11_6.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20538_LC_13_11_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20538_LC_13_11_6.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_0__bdd_4_lut_20538_LC_13_11_6 (
            .in0(N__58856),
            .in1(N__38266),
            .in2(N__60397),
            .in3(N__38233),
            .lcout(n23486),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19795_2_lut_3_lut_LC_13_11_7.C_ON=1'b0;
    defparam i19795_2_lut_3_lut_LC_13_11_7.SEQ_MODE=4'b0000;
    defparam i19795_2_lut_3_lut_LC_13_11_7.LUT_INIT=16'b0010001000000000;
    LogicCell40 i19795_2_lut_3_lut_LC_13_11_7 (
            .in0(N__38582),
            .in1(N__60980),
            .in2(_gnd_net_),
            .in3(N__58648),
            .lcout(n22354),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imiso_83_12612_12613_set_LC_13_12_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12612_12613_set_LC_13_12_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imiso_83_12612_12613_set_LC_13_12_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.imiso_83_12612_12613_set_LC_13_12_0  (
            .in0(N__38191),
            .in1(N__41980),
            .in2(_gnd_net_),
            .in3(N__38443),
            .lcout(\comm_spi.n15340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12612_12613_setC_net ),
            .ce(),
            .sr(N__41914));
    defparam i16457_2_lut_3_lut_LC_13_12_1.C_ON=1'b0;
    defparam i16457_2_lut_3_lut_LC_13_12_1.SEQ_MODE=4'b0000;
    defparam i16457_2_lut_3_lut_LC_13_12_1.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16457_2_lut_3_lut_LC_13_12_1 (
            .in0(N__62610),
            .in1(N__40890),
            .in2(_gnd_net_),
            .in3(N__63990),
            .lcout(n14_adj_1655),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16462_2_lut_3_lut_LC_13_12_2.C_ON=1'b0;
    defparam i16462_2_lut_3_lut_LC_13_12_2.SEQ_MODE=4'b0000;
    defparam i16462_2_lut_3_lut_LC_13_12_2.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16462_2_lut_3_lut_LC_13_12_2 (
            .in0(N__63991),
            .in1(N__43914),
            .in2(_gnd_net_),
            .in3(N__62611),
            .lcout(n14_adj_1608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_13_12_3.C_ON=1'b0;
    defparam i2_3_lut_LC_13_12_3.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_13_12_3.LUT_INIT=16'b1111111110111011;
    LogicCell40 i2_3_lut_LC_13_12_3 (
            .in0(N__62609),
            .in1(N__63988),
            .in2(_gnd_net_),
            .in3(N__51614),
            .lcout(n11254),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_193_LC_13_12_4.C_ON=1'b0;
    defparam i1_2_lut_adj_193_LC_13_12_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_193_LC_13_12_4.LUT_INIT=16'b1111111101010101;
    LogicCell40 i1_2_lut_adj_193_LC_13_12_4 (
            .in0(N__63989),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63603),
            .lcout(n21968),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12520_2_lut_LC_13_12_5.C_ON=1'b0;
    defparam i12520_2_lut_LC_13_12_5.SEQ_MODE=4'b0000;
    defparam i12520_2_lut_LC_13_12_5.LUT_INIT=16'b0101000001010000;
    LogicCell40 i12520_2_lut_LC_13_12_5 (
            .in0(N__63604),
            .in1(_gnd_net_),
            .in2(N__62676),
            .in3(_gnd_net_),
            .lcout(n15238),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12773_2_lut_LC_13_12_6.C_ON=1'b0;
    defparam i12773_2_lut_LC_13_12_6.SEQ_MODE=4'b0000;
    defparam i12773_2_lut_LC_13_12_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12773_2_lut_LC_13_12_6 (
            .in0(_gnd_net_),
            .in1(N__63606),
            .in2(_gnd_net_),
            .in3(N__43458),
            .lcout(n15496),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12780_2_lut_LC_13_12_7.C_ON=1'b0;
    defparam i12780_2_lut_LC_13_12_7.SEQ_MODE=4'b0000;
    defparam i12780_2_lut_LC_13_12_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12780_2_lut_LC_13_12_7 (
            .in0(N__63605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41031),
            .lcout(n15503),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19343_4_lut_LC_13_13_0.C_ON=1'b0;
    defparam i19343_4_lut_LC_13_13_0.SEQ_MODE=4'b0000;
    defparam i19343_4_lut_LC_13_13_0.LUT_INIT=16'b1111110110101000;
    LogicCell40 i19343_4_lut_LC_13_13_0 (
            .in0(N__60595),
            .in1(N__59321),
            .in2(N__38416),
            .in3(N__46864),
            .lcout(),
            .ltout(n22270_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_20503_LC_13_13_1.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_20503_LC_13_13_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_20503_LC_13_13_1.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_2__bdd_4_lut_20503_LC_13_13_1 (
            .in0(N__59995),
            .in1(N__38500),
            .in2(N__38398),
            .in3(N__60992),
            .lcout(),
            .ltout(n23450_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23450_bdd_4_lut_LC_13_13_2.C_ON=1'b0;
    defparam n23450_bdd_4_lut_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam n23450_bdd_4_lut_LC_13_13_2.LUT_INIT=16'b1110010111100000;
    LogicCell40 n23450_bdd_4_lut_LC_13_13_2 (
            .in0(N__60993),
            .in1(N__43474),
            .in2(N__38545),
            .in3(N__38542),
            .lcout(n23453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_0_i112_3_lut_LC_13_13_3.C_ON=1'b0;
    defparam mux_125_Mux_0_i112_3_lut_LC_13_13_3.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_0_i112_3_lut_LC_13_13_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_125_Mux_0_i112_3_lut_LC_13_13_3 (
            .in0(N__48993),
            .in1(N__38458),
            .in2(_gnd_net_),
            .in3(N__60596),
            .lcout(n112_adj_1583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23522_bdd_4_lut_LC_13_13_5.C_ON=1'b0;
    defparam n23522_bdd_4_lut_LC_13_13_5.SEQ_MODE=4'b0000;
    defparam n23522_bdd_4_lut_LC_13_13_5.LUT_INIT=16'b1011101010011000;
    LogicCell40 n23522_bdd_4_lut_LC_13_13_5 (
            .in0(N__38512),
            .in1(N__60594),
            .in2(N__52642),
            .in3(N__44116),
            .lcout(n22267),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_2_i127_3_lut_LC_13_13_6.C_ON=1'b0;
    defparam mux_125_Mux_2_i127_3_lut_LC_13_13_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_2_i127_3_lut_LC_13_13_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_125_Mux_2_i127_3_lut_LC_13_13_6 (
            .in0(N__38494),
            .in1(N__61253),
            .in2(_gnd_net_),
            .in3(N__41413),
            .lcout(comm_buf_0_7_N_543_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_0_i111_3_lut_LC_13_13_7.C_ON=1'b0;
    defparam mux_125_Mux_0_i111_3_lut_LC_13_13_7.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_0_i111_3_lut_LC_13_13_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_125_Mux_0_i111_3_lut_LC_13_13_7 (
            .in0(N__59320),
            .in1(N__38476),
            .in2(_gnd_net_),
            .in3(N__48957),
            .lcout(n111_adj_1584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_254_LC_13_14_0.C_ON=1'b0;
    defparam i4_4_lut_adj_254_LC_13_14_0.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_254_LC_13_14_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_adj_254_LC_13_14_0 (
            .in0(N__44336),
            .in1(N__51985),
            .in2(N__51948),
            .in3(N__49819),
            .lcout(n20_adj_1804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i5_LC_13_14_1.C_ON=1'b0;
    defparam req_data_cnt_i5_LC_13_14_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i5_LC_13_14_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 req_data_cnt_i5_LC_13_14_1 (
            .in0(N__51352),
            .in1(N__51944),
            .in2(_gnd_net_),
            .in3(N__47112),
            .lcout(req_data_cnt_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61874),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i10_LC_13_14_2.C_ON=1'b0;
    defparam req_data_cnt_i10_LC_13_14_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i10_LC_13_14_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i10_LC_13_14_2 (
            .in0(N__39192),
            .in1(N__47424),
            .in2(_gnd_net_),
            .in3(N__51353),
            .lcout(req_data_cnt_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61874),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_253_LC_13_14_3.C_ON=1'b0;
    defparam i5_4_lut_adj_253_LC_13_14_3.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_253_LC_13_14_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_adj_253_LC_13_14_3 (
            .in0(N__50128),
            .in1(N__50086),
            .in2(N__38690),
            .in3(N__39191),
            .lcout(n21_adj_1803),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i12_LC_13_14_4.C_ON=1'b0;
    defparam req_data_cnt_i12_LC_13_14_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i12_LC_13_14_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i12_LC_13_14_4 (
            .in0(N__38694),
            .in1(N__47363),
            .in2(_gnd_net_),
            .in3(N__51354),
            .lcout(req_data_cnt_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61874),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_20478_LC_13_14_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20478_LC_13_14_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20478_LC_13_14_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_20478_LC_13_14_5 (
            .in0(N__38661),
            .in1(N__60631),
            .in2(N__38619),
            .in3(N__59305),
            .lcout(n23348),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19165_3_lut_1_lut_2_lut_LC_13_14_6.C_ON=1'b0;
    defparam i19165_3_lut_1_lut_2_lut_LC_13_14_6.SEQ_MODE=4'b0000;
    defparam i19165_3_lut_1_lut_2_lut_LC_13_14_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 i19165_3_lut_1_lut_2_lut_LC_13_14_6 (
            .in0(_gnd_net_),
            .in1(N__41015),
            .in2(_gnd_net_),
            .in3(N__38584),
            .lcout(n22092),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_stop_331_LC_13_14_7.C_ON=1'b0;
    defparam eis_stop_331_LC_13_14_7.SEQ_MODE=4'b1000;
    defparam eis_stop_331_LC_13_14_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_stop_331_LC_13_14_7 (
            .in0(N__44613),
            .in1(N__43865),
            .in2(_gnd_net_),
            .in3(N__38866),
            .lcout(eis_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61874),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_2_lut_LC_13_15_0.C_ON=1'b1;
    defparam add_122_2_lut_LC_13_15_0.SEQ_MODE=4'b0000;
    defparam add_122_2_lut_LC_13_15_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_2_lut_LC_13_15_0 (
            .in0(N__47815),
            .in1(N__47814),
            .in2(N__47769),
            .in3(N__38560),
            .lcout(n7),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(n20652),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_3_lut_LC_13_15_1.C_ON=1'b1;
    defparam add_122_3_lut_LC_13_15_1.SEQ_MODE=4'b0000;
    defparam add_122_3_lut_LC_13_15_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_3_lut_LC_13_15_1 (
            .in0(N__40204),
            .in1(N__40203),
            .in2(N__47773),
            .in3(N__38557),
            .lcout(n7_adj_1629),
            .ltout(),
            .carryin(n20652),
            .carryout(n20653),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_4_lut_LC_13_15_2.C_ON=1'b1;
    defparam add_122_4_lut_LC_13_15_2.SEQ_MODE=4'b0000;
    defparam add_122_4_lut_LC_13_15_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_4_lut_LC_13_15_2 (
            .in0(N__41790),
            .in1(N__41789),
            .in2(N__47770),
            .in3(N__38554),
            .lcout(n7_adj_1627),
            .ltout(),
            .carryin(n20653),
            .carryout(n20654),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_5_lut_LC_13_15_3.C_ON=1'b1;
    defparam add_122_5_lut_LC_13_15_3.SEQ_MODE=4'b0000;
    defparam add_122_5_lut_LC_13_15_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_5_lut_LC_13_15_3 (
            .in0(N__41625),
            .in1(N__41624),
            .in2(N__47774),
            .in3(N__38551),
            .lcout(n7_adj_1626),
            .ltout(),
            .carryin(n20654),
            .carryout(n20655),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_6_lut_LC_13_15_4.C_ON=1'b1;
    defparam add_122_6_lut_LC_13_15_4.SEQ_MODE=4'b0000;
    defparam add_122_6_lut_LC_13_15_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_6_lut_LC_13_15_4 (
            .in0(N__44164),
            .in1(N__44163),
            .in2(N__47771),
            .in3(N__38548),
            .lcout(n7_adj_1624),
            .ltout(),
            .carryin(n20655),
            .carryout(n20656),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_7_lut_LC_13_15_5.C_ON=1'b1;
    defparam add_122_7_lut_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam add_122_7_lut_LC_13_15_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_7_lut_LC_13_15_5 (
            .in0(N__56503),
            .in1(N__56502),
            .in2(N__47776),
            .in3(N__38887),
            .lcout(n7_adj_1622),
            .ltout(),
            .carryin(n20656),
            .carryout(n20657),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_8_lut_LC_13_15_6.C_ON=1'b1;
    defparam add_122_8_lut_LC_13_15_6.SEQ_MODE=4'b0000;
    defparam add_122_8_lut_LC_13_15_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_8_lut_LC_13_15_6 (
            .in0(N__45148),
            .in1(N__45147),
            .in2(N__47772),
            .in3(N__38884),
            .lcout(n7_adj_1620),
            .ltout(),
            .carryin(n20657),
            .carryout(n20658),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_9_lut_LC_13_15_7.C_ON=1'b1;
    defparam add_122_9_lut_LC_13_15_7.SEQ_MODE=4'b0000;
    defparam add_122_9_lut_LC_13_15_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_9_lut_LC_13_15_7 (
            .in0(N__45007),
            .in1(N__45006),
            .in2(N__47775),
            .in3(N__38881),
            .lcout(n7_adj_1618),
            .ltout(),
            .carryin(n20658),
            .carryout(n20659),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_10_lut_LC_13_16_0.C_ON=1'b1;
    defparam add_122_10_lut_LC_13_16_0.SEQ_MODE=4'b0000;
    defparam add_122_10_lut_LC_13_16_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_10_lut_LC_13_16_0 (
            .in0(N__44953),
            .in1(N__44952),
            .in2(N__47784),
            .in3(N__38878),
            .lcout(n7_adj_1616),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(n20660),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_122_11_lut_LC_13_16_1.C_ON=1'b0;
    defparam add_122_11_lut_LC_13_16_1.SEQ_MODE=4'b0000;
    defparam add_122_11_lut_LC_13_16_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_122_11_lut_LC_13_16_1 (
            .in0(N__42332),
            .in1(N__42333),
            .in2(N__47783),
            .in3(N__38875),
            .lcout(n7_adj_1614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_20523_LC_13_16_2.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20523_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20523_LC_13_16_2.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_0__bdd_4_lut_20523_LC_13_16_2 (
            .in0(N__59438),
            .in1(N__38871),
            .in2(N__60663),
            .in3(N__44080),
            .lcout(n23480),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_58_i14_2_lut_LC_13_16_3.C_ON=1'b0;
    defparam equal_58_i14_2_lut_LC_13_16_3.SEQ_MODE=4'b0000;
    defparam equal_58_i14_2_lut_LC_13_16_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 equal_58_i14_2_lut_LC_13_16_3 (
            .in0(_gnd_net_),
            .in1(N__38839),
            .in2(_gnd_net_),
            .in3(N__38816),
            .lcout(n14_adj_1599),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i13_LC_13_16_4.C_ON=1'b0;
    defparam acadc_skipCount_i13_LC_13_16_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i13_LC_13_16_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 acadc_skipCount_i13_LC_13_16_4 (
            .in0(N__38817),
            .in1(_gnd_net_),
            .in2(N__55283),
            .in3(N__46819),
            .lcout(acadc_skipCount_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61902),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_121_LC_13_16_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_121_LC_13_16_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_121_LC_13_16_5.LUT_INIT=16'b1010101010100010;
    LogicCell40 i1_2_lut_4_lut_adj_121_LC_13_16_5 (
            .in0(N__38793),
            .in1(N__55640),
            .in2(N__38773),
            .in3(N__50891),
            .lcout(n24_adj_1505),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16164_3_lut_LC_13_16_6.C_ON=1'b0;
    defparam i16164_3_lut_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam i16164_3_lut_LC_13_16_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 i16164_3_lut_LC_13_16_6 (
            .in0(N__49293),
            .in1(N__41626),
            .in2(_gnd_net_),
            .in3(N__56469),
            .lcout(n18865),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19240_3_lut_LC_13_16_7.C_ON=1'b0;
    defparam i19240_3_lut_LC_13_16_7.SEQ_MODE=4'b0000;
    defparam i19240_3_lut_LC_13_16_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 i19240_3_lut_LC_13_16_7 (
            .in0(N__39196),
            .in1(N__39133),
            .in2(_gnd_net_),
            .in3(N__59439),
            .lcout(n22167),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_3_i15_4_lut_LC_13_17_0.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_3_i15_4_lut_LC_13_17_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_3_i15_4_lut_LC_13_17_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 comm_state_3__I_0_358_Mux_3_i15_4_lut_LC_13_17_0 (
            .in0(N__41652),
            .in1(N__63607),
            .in2(N__57746),
            .in3(N__41641),
            .lcout(data_index_9_N_236_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_232_LC_13_17_1.C_ON=1'b0;
    defparam i6_4_lut_adj_232_LC_13_17_1.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_232_LC_13_17_1.LUT_INIT=16'b0111110110111110;
    LogicCell40 i6_4_lut_adj_232_LC_13_17_1 (
            .in0(N__38983),
            .in1(N__38965),
            .in2(N__52811),
            .in3(N__55469),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i7_LC_13_17_2.C_ON=1'b0;
    defparam acadc_skipCount_i7_LC_13_17_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i7_LC_13_17_2.LUT_INIT=16'b1100101011001010;
    LogicCell40 acadc_skipCount_i7_LC_13_17_2 (
            .in0(N__55470),
            .in1(N__47517),
            .in2(N__46844),
            .in3(_gnd_net_),
            .lcout(acadc_skipCount_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61916),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i11_LC_13_17_4.C_ON=1'b0;
    defparam acadc_skipCount_i11_LC_13_17_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i11_LC_13_17_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 acadc_skipCount_i11_LC_13_17_4 (
            .in0(N__56839),
            .in1(_gnd_net_),
            .in2(N__46843),
            .in3(N__52742),
            .lcout(acadc_skipCount_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61916),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_234_LC_13_17_5.C_ON=1'b0;
    defparam i5_4_lut_adj_234_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_234_LC_13_17_5.LUT_INIT=16'b0111101111011110;
    LogicCell40 i5_4_lut_adj_234_LC_13_17_5 (
            .in0(N__38947),
            .in1(N__38929),
            .in2(N__39855),
            .in3(N__39908),
            .lcout(),
            .ltout(n21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_238_LC_13_17_6.C_ON=1'b0;
    defparam i14_4_lut_adj_238_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_238_LC_13_17_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_238_LC_13_17_6 (
            .in0(N__38911),
            .in1(N__38902),
            .in2(N__38896),
            .in3(N__38893),
            .lcout(n30_adj_1743),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i12_LC_13_17_7.C_ON=1'b0;
    defparam acadc_skipCount_i12_LC_13_17_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i12_LC_13_17_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 acadc_skipCount_i12_LC_13_17_7 (
            .in0(_gnd_net_),
            .in1(N__47367),
            .in2(N__39856),
            .in3(N__46810),
            .lcout(acadc_skipCount_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61916),
            .ce(),
            .sr(_gnd_net_));
    defparam i16464_2_lut_3_lut_LC_13_18_0.C_ON=1'b0;
    defparam i16464_2_lut_3_lut_LC_13_18_0.SEQ_MODE=4'b0000;
    defparam i16464_2_lut_3_lut_LC_13_18_0.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16464_2_lut_3_lut_LC_13_18_0 (
            .in0(N__63992),
            .in1(N__49232),
            .in2(_gnd_net_),
            .in3(N__62692),
            .lcout(n14_adj_1610),
            .ltout(n14_adj_1610_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i6_LC_13_18_1.C_ON=1'b0;
    defparam acadc_skipCount_i6_LC_13_18_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i6_LC_13_18_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 acadc_skipCount_i6_LC_13_18_1 (
            .in0(N__49683),
            .in1(_gnd_net_),
            .in2(N__39985),
            .in3(N__46847),
            .lcout(acadc_skipCount_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61936),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_240_LC_13_18_2.C_ON=1'b0;
    defparam i1_4_lut_adj_240_LC_13_18_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_240_LC_13_18_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_240_LC_13_18_2 (
            .in0(N__39981),
            .in1(N__49682),
            .in2(N__39964),
            .in3(N__47030),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19239_3_lut_LC_13_18_3.C_ON=1'b0;
    defparam i19239_3_lut_LC_13_18_3.SEQ_MODE=4'b0000;
    defparam i19239_3_lut_LC_13_18_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 i19239_3_lut_LC_13_18_3 (
            .in0(N__39926),
            .in1(N__59441),
            .in2(_gnd_net_),
            .in3(N__39909),
            .lcout(n22166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_4_i23_3_lut_LC_13_18_4.C_ON=1'b0;
    defparam mux_125_Mux_4_i23_3_lut_LC_13_18_4.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_4_i23_3_lut_LC_13_18_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_125_Mux_4_i23_3_lut_LC_13_18_4 (
            .in0(N__59440),
            .in1(_gnd_net_),
            .in2(N__39879),
            .in3(N__39854),
            .lcout(n23_adj_1783),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i0_LC_13_18_5.C_ON=1'b0;
    defparam acadc_skipCount_i0_LC_13_18_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i0_LC_13_18_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i0_LC_13_18_5 (
            .in0(N__47031),
            .in1(N__57856),
            .in2(N__49142),
            .in3(N__46848),
            .lcout(acadc_skipCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61936),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i9_LC_13_18_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i9_LC_13_18_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i9_LC_13_18_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i9_LC_13_18_7  (
            .in0(N__39806),
            .in1(N__39385),
            .in2(N__39223),
            .in3(N__52704),
            .lcout(buf_adcdata_iac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61936),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i1_LC_13_19_0.C_ON=1'b0;
    defparam buf_dds0_i1_LC_13_19_0.SEQ_MODE=4'b1000;
    defparam buf_dds0_i1_LC_13_19_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_dds0_i1_LC_13_19_0 (
            .in0(N__50737),
            .in1(N__52091),
            .in2(N__57880),
            .in3(N__42152),
            .lcout(buf_dds0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61952),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i1_LC_13_19_1.C_ON=1'b0;
    defparam data_index_i1_LC_13_19_1.SEQ_MODE=4'b1000;
    defparam data_index_i1_LC_13_19_1.LUT_INIT=16'b0000110010101010;
    LogicCell40 data_index_i1_LC_13_19_1 (
            .in0(N__40171),
            .in1(N__40180),
            .in2(N__57871),
            .in3(N__63609),
            .lcout(data_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61952),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i8_LC_13_19_2.C_ON=1'b0;
    defparam buf_dds0_i8_LC_13_19_2.SEQ_MODE=4'b1000;
    defparam buf_dds0_i8_LC_13_19_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 buf_dds0_i8_LC_13_19_2 (
            .in0(N__50736),
            .in1(N__48857),
            .in2(_gnd_net_),
            .in3(N__40226),
            .lcout(buf_dds0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61952),
            .ce(),
            .sr(_gnd_net_));
    defparam i6651_3_lut_LC_13_19_3.C_ON=1'b0;
    defparam i6651_3_lut_LC_13_19_3.SEQ_MODE=4'b0000;
    defparam i6651_3_lut_LC_13_19_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6651_3_lut_LC_13_19_3 (
            .in0(N__52090),
            .in1(N__40196),
            .in2(_gnd_net_),
            .in3(N__56474),
            .lcout(n8_adj_1630),
            .ltout(n8_adj_1630_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_1_i15_4_lut_LC_13_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_1_i15_4_lut_LC_13_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_1_i15_4_lut_LC_13_19_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_state_3__I_0_358_Mux_1_i15_4_lut_LC_13_19_4 (
            .in0(N__63608),
            .in1(N__57833),
            .in2(N__40174),
            .in3(N__40170),
            .lcout(data_index_9_N_236_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i3_LC_13_19_5.C_ON=1'b0;
    defparam buf_dds0_i3_LC_13_19_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i3_LC_13_19_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_dds0_i3_LC_13_19_5 (
            .in0(N__57834),
            .in1(N__50738),
            .in2(N__49311),
            .in3(N__40064),
            .lcout(buf_dds0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61952),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i3_LC_13_19_6.C_ON=1'b0;
    defparam buf_control_i3_LC_13_19_6.SEQ_MODE=4'b1000;
    defparam buf_control_i3_LC_13_19_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_control_i3_LC_13_19_6 (
            .in0(N__56849),
            .in1(N__46750),
            .in2(_gnd_net_),
            .in3(N__52763),
            .lcout(SELIRNG1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61952),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.MOSI_31_LC_13_20_4 .C_ON=1'b0;
    defparam \SIG_DDS.MOSI_31_LC_13_20_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.MOSI_31_LC_13_20_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \SIG_DDS.MOSI_31_LC_13_20_4  (
            .in0(N__40045),
            .in1(N__40011),
            .in2(_gnd_net_),
            .in3(N__50368),
            .lcout(DDS_MOSI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61970),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_12598_12599_set_LC_14_2_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12598_12599_set_LC_14_2_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.iclk_40_12598_12599_set_LC_14_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12598_12599_set_LC_14_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42498),
            .lcout(\comm_spi.n15326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61824),
            .ce(),
            .sr(N__42166));
    defparam \comm_spi.i20203_4_lut_3_lut_LC_14_3_2 .C_ON=1'b0;
    defparam \comm_spi.i20203_4_lut_3_lut_LC_14_3_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20203_4_lut_3_lut_LC_14_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i20203_4_lut_3_lut_LC_14_3_2  (
            .in0(N__42499),
            .in1(N__40000),
            .in2(_gnd_net_),
            .in3(N__57130),
            .lcout(\comm_spi.n24016 ),
            .ltout(\comm_spi.n24016_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12600_3_lut_LC_14_3_3 .C_ON=1'b0;
    defparam \comm_spi.i12600_3_lut_LC_14_3_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12600_3_lut_LC_14_3_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.i12600_3_lut_LC_14_3_3  (
            .in0(N__39994),
            .in1(_gnd_net_),
            .in2(N__39988),
            .in3(N__42766),
            .lcout(\comm_spi.iclk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12594_12595_set_LC_14_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12594_12595_set_LC_14_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i0_12594_12595_set_LC_14_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_12594_12595_set_LC_14_4_0  (
            .in0(N__64676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n15322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53617),
            .ce(),
            .sr(N__40276));
    defparam secclk_cnt_3785_3786__i1_LC_14_5_0.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i1_LC_14_5_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i1_LC_14_5_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i1_LC_14_5_0 (
            .in0(_gnd_net_),
            .in1(N__45223),
            .in2(_gnd_net_),
            .in3(N__40264),
            .lcout(secclk_cnt_0),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(n20790),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i2_LC_14_5_1.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i2_LC_14_5_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i2_LC_14_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i2_LC_14_5_1 (
            .in0(_gnd_net_),
            .in1(N__42405),
            .in2(_gnd_net_),
            .in3(N__40261),
            .lcout(secclk_cnt_1),
            .ltout(),
            .carryin(n20790),
            .carryout(n20791),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i3_LC_14_5_2.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i3_LC_14_5_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i3_LC_14_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i3_LC_14_5_2 (
            .in0(_gnd_net_),
            .in1(N__42865),
            .in2(_gnd_net_),
            .in3(N__40258),
            .lcout(secclk_cnt_2),
            .ltout(),
            .carryin(n20791),
            .carryout(n20792),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i4_LC_14_5_3.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i4_LC_14_5_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i4_LC_14_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i4_LC_14_5_3 (
            .in0(_gnd_net_),
            .in1(N__42922),
            .in2(_gnd_net_),
            .in3(N__40255),
            .lcout(secclk_cnt_3),
            .ltout(),
            .carryin(n20792),
            .carryout(n20793),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i5_LC_14_5_4.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i5_LC_14_5_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i5_LC_14_5_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i5_LC_14_5_4 (
            .in0(_gnd_net_),
            .in1(N__45168),
            .in2(_gnd_net_),
            .in3(N__40252),
            .lcout(secclk_cnt_4),
            .ltout(),
            .carryin(n20793),
            .carryout(n20794),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i6_LC_14_5_5.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i6_LC_14_5_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i6_LC_14_5_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i6_LC_14_5_5 (
            .in0(_gnd_net_),
            .in1(N__42391),
            .in2(_gnd_net_),
            .in3(N__40249),
            .lcout(secclk_cnt_5),
            .ltout(),
            .carryin(n20794),
            .carryout(n20795),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i7_LC_14_5_6.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i7_LC_14_5_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i7_LC_14_5_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i7_LC_14_5_6 (
            .in0(_gnd_net_),
            .in1(N__42961),
            .in2(_gnd_net_),
            .in3(N__40246),
            .lcout(secclk_cnt_6),
            .ltout(),
            .carryin(n20795),
            .carryout(n20796),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i8_LC_14_5_7.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i8_LC_14_5_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i8_LC_14_5_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i8_LC_14_5_7 (
            .in0(_gnd_net_),
            .in1(N__42892),
            .in2(_gnd_net_),
            .in3(N__40243),
            .lcout(secclk_cnt_7),
            .ltout(),
            .carryin(n20796),
            .carryout(n20797),
            .clk(N__48400),
            .ce(),
            .sr(N__42846));
    defparam secclk_cnt_3785_3786__i9_LC_14_6_0.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i9_LC_14_6_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i9_LC_14_6_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i9_LC_14_6_0 (
            .in0(_gnd_net_),
            .in1(N__42418),
            .in2(_gnd_net_),
            .in3(N__40315),
            .lcout(secclk_cnt_8),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(n20798),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i10_LC_14_6_1.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i10_LC_14_6_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i10_LC_14_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i10_LC_14_6_1 (
            .in0(_gnd_net_),
            .in1(N__42994),
            .in2(_gnd_net_),
            .in3(N__40312),
            .lcout(secclk_cnt_9),
            .ltout(),
            .carryin(n20798),
            .carryout(n20799),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i11_LC_14_6_2.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i11_LC_14_6_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i11_LC_14_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i11_LC_14_6_2 (
            .in0(_gnd_net_),
            .in1(N__42936),
            .in2(_gnd_net_),
            .in3(N__40309),
            .lcout(secclk_cnt_10),
            .ltout(),
            .carryin(n20799),
            .carryout(n20800),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i12_LC_14_6_3.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i12_LC_14_6_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i12_LC_14_6_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i12_LC_14_6_3 (
            .in0(_gnd_net_),
            .in1(N__45183),
            .in2(_gnd_net_),
            .in3(N__40306),
            .lcout(secclk_cnt_11),
            .ltout(),
            .carryin(n20800),
            .carryout(n20801),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i13_LC_14_6_4.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i13_LC_14_6_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i13_LC_14_6_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i13_LC_14_6_4 (
            .in0(_gnd_net_),
            .in1(N__40341),
            .in2(_gnd_net_),
            .in3(N__40303),
            .lcout(secclk_cnt_12),
            .ltout(),
            .carryin(n20801),
            .carryout(n20802),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i14_LC_14_6_5.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i14_LC_14_6_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i14_LC_14_6_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i14_LC_14_6_5 (
            .in0(_gnd_net_),
            .in1(N__42879),
            .in2(_gnd_net_),
            .in3(N__40300),
            .lcout(secclk_cnt_13),
            .ltout(),
            .carryin(n20802),
            .carryout(n20803),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i15_LC_14_6_6.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i15_LC_14_6_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i15_LC_14_6_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i15_LC_14_6_6 (
            .in0(_gnd_net_),
            .in1(N__42949),
            .in2(_gnd_net_),
            .in3(N__40297),
            .lcout(secclk_cnt_14),
            .ltout(),
            .carryin(n20803),
            .carryout(n20804),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i16_LC_14_6_7.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i16_LC_14_6_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i16_LC_14_6_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i16_LC_14_6_7 (
            .in0(_gnd_net_),
            .in1(N__42430),
            .in2(_gnd_net_),
            .in3(N__40294),
            .lcout(secclk_cnt_15),
            .ltout(),
            .carryin(n20804),
            .carryout(n20805),
            .clk(N__48401),
            .ce(),
            .sr(N__42845));
    defparam secclk_cnt_3785_3786__i17_LC_14_7_0.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i17_LC_14_7_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i17_LC_14_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i17_LC_14_7_0 (
            .in0(_gnd_net_),
            .in1(N__42904),
            .in2(_gnd_net_),
            .in3(N__40291),
            .lcout(secclk_cnt_16),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(n20806),
            .clk(N__48403),
            .ce(),
            .sr(N__42847));
    defparam secclk_cnt_3785_3786__i18_LC_14_7_1.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i18_LC_14_7_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i18_LC_14_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i18_LC_14_7_1 (
            .in0(_gnd_net_),
            .in1(N__42981),
            .in2(_gnd_net_),
            .in3(N__40387),
            .lcout(secclk_cnt_17),
            .ltout(),
            .carryin(n20806),
            .carryout(n20807),
            .clk(N__48403),
            .ce(),
            .sr(N__42847));
    defparam secclk_cnt_3785_3786__i19_LC_14_7_2.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i19_LC_14_7_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i19_LC_14_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i19_LC_14_7_2 (
            .in0(_gnd_net_),
            .in1(N__45207),
            .in2(_gnd_net_),
            .in3(N__40384),
            .lcout(secclk_cnt_18),
            .ltout(),
            .carryin(n20807),
            .carryout(n20808),
            .clk(N__48403),
            .ce(),
            .sr(N__42847));
    defparam secclk_cnt_3785_3786__i20_LC_14_7_3.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i20_LC_14_7_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i20_LC_14_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i20_LC_14_7_3 (
            .in0(_gnd_net_),
            .in1(N__40369),
            .in2(_gnd_net_),
            .in3(N__40381),
            .lcout(secclk_cnt_19),
            .ltout(),
            .carryin(n20808),
            .carryout(n20809),
            .clk(N__48403),
            .ce(),
            .sr(N__42847));
    defparam secclk_cnt_3785_3786__i21_LC_14_7_4.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i21_LC_14_7_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i21_LC_14_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i21_LC_14_7_4 (
            .in0(_gnd_net_),
            .in1(N__43018),
            .in2(_gnd_net_),
            .in3(N__40378),
            .lcout(secclk_cnt_20),
            .ltout(),
            .carryin(n20809),
            .carryout(n20810),
            .clk(N__48403),
            .ce(),
            .sr(N__42847));
    defparam secclk_cnt_3785_3786__i22_LC_14_7_5.C_ON=1'b1;
    defparam secclk_cnt_3785_3786__i22_LC_14_7_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i22_LC_14_7_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i22_LC_14_7_5 (
            .in0(_gnd_net_),
            .in1(N__40357),
            .in2(_gnd_net_),
            .in3(N__40375),
            .lcout(secclk_cnt_21),
            .ltout(),
            .carryin(n20810),
            .carryout(n20811),
            .clk(N__48403),
            .ce(),
            .sr(N__42847));
    defparam secclk_cnt_3785_3786__i23_LC_14_7_6.C_ON=1'b0;
    defparam secclk_cnt_3785_3786__i23_LC_14_7_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3785_3786__i23_LC_14_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3785_3786__i23_LC_14_7_6 (
            .in0(_gnd_net_),
            .in1(N__40327),
            .in2(_gnd_net_),
            .in3(N__40372),
            .lcout(secclk_cnt_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48403),
            .ce(),
            .sr(N__42847));
    defparam i6_4_lut_adj_204_LC_14_8_0.C_ON=1'b0;
    defparam i6_4_lut_adj_204_LC_14_8_0.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_204_LC_14_8_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_adj_204_LC_14_8_0 (
            .in0(N__40368),
            .in1(N__40356),
            .in2(N__40345),
            .in3(N__40326),
            .lcout(n14_adj_1678),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_287_LC_14_8_1.C_ON=1'b0;
    defparam i1_4_lut_adj_287_LC_14_8_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_287_LC_14_8_1.LUT_INIT=16'b1000110010001000;
    LogicCell40 i1_4_lut_adj_287_LC_14_8_1 (
            .in0(N__63483),
            .in1(N__63163),
            .in2(N__64101),
            .in3(N__51542),
            .lcout(n15378),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_333_LC_14_8_2.C_ON=1'b0;
    defparam i1_4_lut_adj_333_LC_14_8_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_333_LC_14_8_2.LUT_INIT=16'b1010101010000000;
    LogicCell40 i1_4_lut_adj_333_LC_14_8_2 (
            .in0(N__63162),
            .in1(N__64090),
            .in2(N__51546),
            .in3(N__63482),
            .lcout(n13076),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16454_2_lut_3_lut_LC_14_8_3.C_ON=1'b0;
    defparam i16454_2_lut_3_lut_LC_14_8_3.SEQ_MODE=4'b0000;
    defparam i16454_2_lut_3_lut_LC_14_8_3.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16454_2_lut_3_lut_LC_14_8_3 (
            .in0(N__64091),
            .in1(N__40563),
            .in2(_gnd_net_),
            .in3(N__62624),
            .lcout(n14_adj_1652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i1_LC_14_8_4.C_ON=1'b0;
    defparam comm_buf_6__i1_LC_14_8_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i1_LC_14_8_4.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i1_LC_14_8_4 (
            .in0(N__40465),
            .in1(N__63484),
            .in2(N__54823),
            .in3(N__45570),
            .lcout(comm_buf_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61836),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_127_Mux_2_i30_3_lut_LC_14_8_5.C_ON=1'b0;
    defparam mux_127_Mux_2_i30_3_lut_LC_14_8_5.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_2_i30_3_lut_LC_14_8_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_127_Mux_2_i30_3_lut_LC_14_8_5 (
            .in0(N__40450),
            .in1(N__40438),
            .in2(_gnd_net_),
            .in3(N__60991),
            .lcout(n30_adj_1708),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_215_LC_14_8_6.C_ON=1'b0;
    defparam i1_4_lut_adj_215_LC_14_8_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_215_LC_14_8_6.LUT_INIT=16'b1011000010100000;
    LogicCell40 i1_4_lut_adj_215_LC_14_8_6 (
            .in0(N__63485),
            .in1(N__64095),
            .in2(N__63189),
            .in3(N__56884),
            .lcout(n12585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i13_LC_14_8_7.C_ON=1'b0;
    defparam buf_dds0_i13_LC_14_8_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i13_LC_14_8_7.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i13_LC_14_8_7 (
            .in0(N__57764),
            .in1(N__55529),
            .in2(N__45339),
            .in3(N__50688),
            .lcout(buf_dds0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61836),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_7_i2_3_lut_LC_14_9_0.C_ON=1'b0;
    defparam mux_134_Mux_7_i2_3_lut_LC_14_9_0.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_7_i2_3_lut_LC_14_9_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_134_Mux_7_i2_3_lut_LC_14_9_0 (
            .in0(N__40424),
            .in1(N__40783),
            .in2(_gnd_net_),
            .in3(N__54407),
            .lcout(n2_adj_1663),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19758_2_lut_LC_14_9_1.C_ON=1'b0;
    defparam i19758_2_lut_LC_14_9_1.SEQ_MODE=4'b0000;
    defparam i19758_2_lut_LC_14_9_1.LUT_INIT=16'b0100010001000100;
    LogicCell40 i19758_2_lut_LC_14_9_1 (
            .in0(N__54408),
            .in1(N__43071),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n22331_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_20429_LC_14_9_2.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_20429_LC_14_9_2.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_20429_LC_14_9_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_1__bdd_4_lut_20429_LC_14_9_2 (
            .in0(N__40669),
            .in1(N__54599),
            .in2(N__40399),
            .in3(N__51822),
            .lcout(),
            .ltout(n23360_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i7_LC_14_9_3.C_ON=1'b0;
    defparam comm_tx_buf_i7_LC_14_9_3.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i7_LC_14_9_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 comm_tx_buf_i7_LC_14_9_3 (
            .in0(N__54600),
            .in1(N__40663),
            .in2(N__40396),
            .in3(N__40393),
            .lcout(comm_tx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61842),
            .ce(N__46403),
            .sr(N__46351));
    defparam mux_134_Mux_7_i4_3_lut_LC_14_9_4.C_ON=1'b0;
    defparam mux_134_Mux_7_i4_3_lut_LC_14_9_4.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_7_i4_3_lut_LC_14_9_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_134_Mux_7_i4_3_lut_LC_14_9_4 (
            .in0(N__53908),
            .in1(N__43147),
            .in2(_gnd_net_),
            .in3(N__54405),
            .lcout(n4_adj_1664),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_7_i1_3_lut_LC_14_9_5.C_ON=1'b0;
    defparam mux_134_Mux_7_i1_3_lut_LC_14_9_5.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_7_i1_3_lut_LC_14_9_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_134_Mux_7_i1_3_lut_LC_14_9_5 (
            .in0(N__54406),
            .in1(N__46622),
            .in2(_gnd_net_),
            .in3(N__55841),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20213_4_lut_3_lut_LC_14_9_6 .C_ON=1'b0;
    defparam \comm_spi.i20213_4_lut_3_lut_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20213_4_lut_3_lut_LC_14_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i20213_4_lut_3_lut_LC_14_9_6  (
            .in0(N__41963),
            .in1(N__40643),
            .in2(_gnd_net_),
            .in3(N__57111),
            .lcout(\comm_spi.n15333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_9_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_9_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \comm_spi.RESET_I_0_100_2_lut_LC_14_9_7  (
            .in0(N__57112),
            .in1(_gnd_net_),
            .in2(N__40650),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_862 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_2_i4_3_lut_LC_14_10_0.C_ON=1'b0;
    defparam mux_134_Mux_2_i4_3_lut_LC_14_10_0.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_2_i4_3_lut_LC_14_10_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_134_Mux_2_i4_3_lut_LC_14_10_0 (
            .in0(N__43354),
            .in1(N__54838),
            .in2(_gnd_net_),
            .in3(N__54398),
            .lcout(n4_adj_1673),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19747_2_lut_LC_14_10_1.C_ON=1'b0;
    defparam i19747_2_lut_LC_14_10_1.SEQ_MODE=4'b0000;
    defparam i19747_2_lut_LC_14_10_1.LUT_INIT=16'b0101000001010000;
    LogicCell40 i19747_2_lut_LC_14_10_1 (
            .in0(N__54399),
            .in1(_gnd_net_),
            .in2(N__45517),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n22342_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_20454_LC_14_10_2.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_20454_LC_14_10_2.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_20454_LC_14_10_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_1__bdd_4_lut_20454_LC_14_10_2 (
            .in0(N__40597),
            .in1(N__54601),
            .in2(N__40591),
            .in3(N__51830),
            .lcout(n23396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_2_i1_3_lut_LC_14_10_3.C_ON=1'b0;
    defparam mux_134_Mux_2_i1_3_lut_LC_14_10_3.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_2_i1_3_lut_LC_14_10_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_134_Mux_2_i1_3_lut_LC_14_10_3 (
            .in0(N__54401),
            .in1(_gnd_net_),
            .in2(N__40939),
            .in3(N__52926),
            .lcout(),
            .ltout(n1_adj_1671_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i2_LC_14_10_4.C_ON=1'b0;
    defparam comm_tx_buf_i2_LC_14_10_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i2_LC_14_10_4.LUT_INIT=16'b1011101010011000;
    LogicCell40 comm_tx_buf_i2_LC_14_10_4 (
            .in0(N__40588),
            .in1(N__54602),
            .in2(N__40582),
            .in3(N__40579),
            .lcout(comm_tx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61848),
            .ce(N__46431),
            .sr(N__46349));
    defparam mux_134_Mux_2_i2_3_lut_LC_14_10_5.C_ON=1'b0;
    defparam mux_134_Mux_2_i2_3_lut_LC_14_10_5.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_2_i2_3_lut_LC_14_10_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_134_Mux_2_i2_3_lut_LC_14_10_5 (
            .in0(N__54400),
            .in1(N__41128),
            .in2(_gnd_net_),
            .in3(N__40973),
            .lcout(n2_adj_1672),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10481_3_lut_LC_14_10_6.C_ON=1'b0;
    defparam i10481_3_lut_LC_14_10_6.SEQ_MODE=4'b0000;
    defparam i10481_3_lut_LC_14_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i10481_3_lut_LC_14_10_6 (
            .in0(N__40974),
            .in1(N__40925),
            .in2(_gnd_net_),
            .in3(N__46163),
            .lcout(n13207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_14_10_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_14_10_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_105_2_lut_LC_14_10_7  (
            .in0(N__57110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40845),
            .lcout(\comm_spi.data_tx_7__N_877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i0_LC_14_11_0.C_ON=1'b0;
    defparam comm_buf_3__i0_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i0_LC_14_11_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i0_LC_14_11_0 (
            .in0(N__54016),
            .in1(N__40816),
            .in2(_gnd_net_),
            .in3(N__62653),
            .lcout(comm_buf_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam comm_buf_3__i7_LC_14_11_1.C_ON=1'b0;
    defparam comm_buf_3__i7_LC_14_11_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i7_LC_14_11_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_3__i7_LC_14_11_1 (
            .in0(N__62652),
            .in1(_gnd_net_),
            .in2(N__55936),
            .in3(N__40801),
            .lcout(comm_buf_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam comm_buf_3__i6_LC_14_11_2.C_ON=1'b0;
    defparam comm_buf_3__i6_LC_14_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i6_LC_14_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i6_LC_14_11_2 (
            .in0(N__53879),
            .in1(N__40774),
            .in2(_gnd_net_),
            .in3(N__62656),
            .lcout(comm_buf_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam comm_buf_3__i5_LC_14_11_3.C_ON=1'b0;
    defparam comm_buf_3__i5_LC_14_11_3.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i5_LC_14_11_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_3__i5_LC_14_11_3 (
            .in0(N__62648),
            .in1(_gnd_net_),
            .in2(N__55194),
            .in3(N__40738),
            .lcout(comm_buf_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam comm_buf_3__i4_LC_14_11_4.C_ON=1'b0;
    defparam comm_buf_3__i4_LC_14_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i4_LC_14_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i4_LC_14_11_4 (
            .in0(N__55077),
            .in1(N__40717),
            .in2(_gnd_net_),
            .in3(N__62655),
            .lcout(comm_buf_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam comm_buf_3__i3_LC_14_11_5.C_ON=1'b0;
    defparam comm_buf_3__i3_LC_14_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i3_LC_14_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i3_LC_14_11_5 (
            .in0(N__62647),
            .in1(N__62790),
            .in2(_gnd_net_),
            .in3(N__40687),
            .lcout(comm_buf_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam comm_buf_3__i2_LC_14_11_6.C_ON=1'b0;
    defparam comm_buf_3__i2_LC_14_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i2_LC_14_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i2_LC_14_11_6 (
            .in0(N__54938),
            .in1(N__41143),
            .in2(_gnd_net_),
            .in3(N__62654),
            .lcout(comm_buf_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam comm_buf_3__i1_LC_14_11_7.C_ON=1'b0;
    defparam comm_buf_3__i1_LC_14_11_7.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i1_LC_14_11_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 comm_buf_3__i1_LC_14_11_7 (
            .in0(N__54816),
            .in1(_gnd_net_),
            .in2(N__62685),
            .in3(N__41122),
            .lcout(comm_buf_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61855),
            .ce(N__41038),
            .sr(N__41095));
    defparam mux_127_Mux_2_i127_3_lut_LC_14_12_0.C_ON=1'b0;
    defparam mux_127_Mux_2_i127_3_lut_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam mux_127_Mux_2_i127_3_lut_LC_14_12_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_127_Mux_2_i127_3_lut_LC_14_12_0 (
            .in0(N__41080),
            .in1(N__41071),
            .in2(_gnd_net_),
            .in3(N__61182),
            .lcout(comm_buf_2_7_N_575_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_316_LC_14_12_1.C_ON=1'b0;
    defparam i1_3_lut_adj_316_LC_14_12_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_316_LC_14_12_1.LUT_INIT=16'b1100110010001000;
    LogicCell40 i1_3_lut_adj_316_LC_14_12_1 (
            .in0(N__54136),
            .in1(N__54085),
            .in2(_gnd_net_),
            .in3(N__48889),
            .lcout(n12880),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i6_LC_14_12_2.C_ON=1'b0;
    defparam comm_cmd_i6_LC_14_12_2.SEQ_MODE=4'b1000;
    defparam comm_cmd_i6_LC_14_12_2.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i6_LC_14_12_2 (
            .in0(N__45933),
            .in1(N__45995),
            .in2(N__53893),
            .in3(N__61183),
            .lcout(comm_cmd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61863),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_14_12_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_14_12_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_14_12_3.LUT_INIT=16'b0000000010000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_14_12_3 (
            .in0(N__58585),
            .in1(N__58469),
            .in2(N__61260),
            .in3(N__60793),
            .lcout(n21886),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_310_LC_14_12_4.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_310_LC_14_12_4.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_310_LC_14_12_4.LUT_INIT=16'b1111111111011111;
    LogicCell40 i2_3_lut_4_lut_adj_310_LC_14_12_4 (
            .in0(N__60792),
            .in1(N__61178),
            .in2(N__58491),
            .in3(N__58584),
            .lcout(n12),
            .ltout(n12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_14_12_5.C_ON=1'b0;
    defparam i1_2_lut_LC_14_12_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_14_12_5.LUT_INIT=16'b1111001111110011;
    LogicCell40 i1_2_lut_LC_14_12_5 (
            .in0(_gnd_net_),
            .in1(N__58836),
            .in2(N__40981),
            .in3(_gnd_net_),
            .lcout(n12015),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_338_LC_14_12_6.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_338_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_338_LC_14_12_6.LUT_INIT=16'b1111111111111101;
    LogicCell40 i1_2_lut_4_lut_adj_338_LC_14_12_6 (
            .in0(N__59672),
            .in1(N__41349),
            .in2(N__63075),
            .in3(N__41400),
            .lcout(n11258),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12830_2_lut_3_lut_LC_14_12_7.C_ON=1'b0;
    defparam i12830_2_lut_3_lut_LC_14_12_7.SEQ_MODE=4'b0000;
    defparam i12830_2_lut_3_lut_LC_14_12_7.LUT_INIT=16'b1111000011000000;
    LogicCell40 i12830_2_lut_3_lut_LC_14_12_7 (
            .in0(_gnd_net_),
            .in1(N__64089),
            .in2(N__44040),
            .in3(N__62615),
            .lcout(n15553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16466_2_lut_3_lut_LC_14_13_0.C_ON=1'b0;
    defparam i16466_2_lut_3_lut_LC_14_13_0.SEQ_MODE=4'b0000;
    defparam i16466_2_lut_3_lut_LC_14_13_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 i16466_2_lut_3_lut_LC_14_13_0 (
            .in0(N__52909),
            .in1(N__62689),
            .in2(_gnd_net_),
            .in3(N__64088),
            .lcout(n14_adj_1612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23288_bdd_4_lut_LC_14_13_1.C_ON=1'b0;
    defparam n23288_bdd_4_lut_LC_14_13_1.SEQ_MODE=4'b0000;
    defparam n23288_bdd_4_lut_LC_14_13_1.LUT_INIT=16'b1010101011100100;
    LogicCell40 n23288_bdd_4_lut_LC_14_13_1 (
            .in0(N__43660),
            .in1(N__41326),
            .in2(N__41311),
            .in3(N__59999),
            .lcout(n23291),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_14_13_2.C_ON=1'b0;
    defparam i3_4_lut_LC_14_13_2.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_14_13_2.LUT_INIT=16'b1111111111111101;
    LogicCell40 i3_4_lut_LC_14_13_2 (
            .in0(N__60000),
            .in1(N__63078),
            .in2(N__41266),
            .in3(N__60468),
            .lcout(n9324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i3_LC_14_13_4.C_ON=1'b0;
    defparam req_data_cnt_i3_LC_14_13_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i3_LC_14_13_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 req_data_cnt_i3_LC_14_13_4 (
            .in0(N__51348),
            .in1(_gnd_net_),
            .in2(N__48941),
            .in3(N__44340),
            .lcout(req_data_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61875),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_372_i8_2_lut_LC_14_13_5.C_ON=1'b0;
    defparam comm_cmd_6__I_0_372_i8_2_lut_LC_14_13_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_372_i8_2_lut_LC_14_13_5.LUT_INIT=16'b1111111101010101;
    LogicCell40 comm_cmd_6__I_0_372_i8_2_lut_LC_14_13_5 (
            .in0(N__60469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60001),
            .lcout(),
            .ltout(n8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_210_LC_14_13_6.C_ON=1'b0;
    defparam i2_4_lut_adj_210_LC_14_13_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_210_LC_14_13_6.LUT_INIT=16'b0000000000000100;
    LogicCell40 i2_4_lut_adj_210_LC_14_13_6 (
            .in0(N__41265),
            .in1(N__63726),
            .in2(N__41254),
            .in3(N__63079),
            .lcout(n11172),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_3_i19_3_lut_LC_14_13_7.C_ON=1'b0;
    defparam mux_126_Mux_3_i19_3_lut_LC_14_13_7.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_3_i19_3_lut_LC_14_13_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_3_i19_3_lut_LC_14_13_7 (
            .in0(N__41251),
            .in1(N__41220),
            .in2(_gnd_net_),
            .in3(N__59306),
            .lcout(n19_adj_1739),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_73_LC_14_14_1.C_ON=1'b0;
    defparam i1_4_lut_adj_73_LC_14_14_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_73_LC_14_14_1.LUT_INIT=16'b1111010000000000;
    LogicCell40 i1_4_lut_adj_73_LC_14_14_1 (
            .in0(N__63081),
            .in1(N__41194),
            .in2(N__57844),
            .in3(N__63725),
            .lcout(n13211),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_14_14_2.C_ON=1'b0;
    defparam i4_4_lut_LC_14_14_2.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_14_14_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_LC_14_14_2 (
            .in0(N__41164),
            .in1(N__41533),
            .in2(N__44296),
            .in3(N__51917),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_7_i23_3_lut_LC_14_14_3.C_ON=1'b0;
    defparam mux_125_Mux_7_i23_3_lut_LC_14_14_3.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_7_i23_3_lut_LC_14_14_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_125_Mux_7_i23_3_lut_LC_14_14_3 (
            .in0(N__46024),
            .in1(N__59307),
            .in2(_gnd_net_),
            .in3(N__41512),
            .lcout(n23_adj_1756),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_313_LC_14_14_4.C_ON=1'b0;
    defparam i14_4_lut_adj_313_LC_14_14_4.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_313_LC_14_14_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_313_LC_14_14_4 (
            .in0(N__51685),
            .in1(N__41470),
            .in2(N__44092),
            .in3(N__43573),
            .lcout(n30_adj_1769),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23546_bdd_4_lut_LC_14_14_5.C_ON=1'b0;
    defparam n23546_bdd_4_lut_LC_14_14_5.SEQ_MODE=4'b0000;
    defparam n23546_bdd_4_lut_LC_14_14_5.LUT_INIT=16'b1110111000110000;
    LogicCell40 n23546_bdd_4_lut_LC_14_14_5 (
            .in0(N__41455),
            .in1(N__60002),
            .in2(N__41446),
            .in3(N__44140),
            .lcout(),
            .ltout(n23549_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19247_3_lut_LC_14_14_6.C_ON=1'b0;
    defparam i19247_3_lut_LC_14_14_6.SEQ_MODE=4'b0000;
    defparam i19247_3_lut_LC_14_14_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 i19247_3_lut_LC_14_14_6 (
            .in0(_gnd_net_),
            .in1(N__41431),
            .in2(N__41416),
            .in3(N__60994),
            .lcout(n22174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i0_LC_14_15_0.C_ON=1'b0;
    defparam comm_length_i0_LC_14_15_0.SEQ_MODE=4'b1000;
    defparam comm_length_i0_LC_14_15_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_length_i0_LC_14_15_0 (
            .in0(N__44134),
            .in1(N__61348),
            .in2(_gnd_net_),
            .in3(N__41407),
            .lcout(comm_length_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61903),
            .ce(N__46678),
            .sr(N__48291));
    defparam comm_length_i1_LC_14_15_1.C_ON=1'b0;
    defparam comm_length_i1_LC_14_15_1.SEQ_MODE=4'b1000;
    defparam comm_length_i1_LC_14_15_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_length_i1_LC_14_15_1 (
            .in0(N__61347),
            .in1(N__41389),
            .in2(_gnd_net_),
            .in3(N__60664),
            .lcout(comm_length_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61903),
            .ce(N__46678),
            .sr(N__48291));
    defparam i1_2_lut_adj_244_LC_14_15_2.C_ON=1'b0;
    defparam i1_2_lut_adj_244_LC_14_15_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_244_LC_14_15_2.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_244_LC_14_15_2 (
            .in0(_gnd_net_),
            .in1(N__43818),
            .in2(_gnd_net_),
            .in3(N__41544),
            .lcout(n17650),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_331_LC_14_15_3.C_ON=1'b0;
    defparam i1_2_lut_adj_331_LC_14_15_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_331_LC_14_15_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_331_LC_14_15_3 (
            .in0(_gnd_net_),
            .in1(N__63080),
            .in2(_gnd_net_),
            .in3(N__41353),
            .lcout(n21983),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20055_2_lut_LC_14_15_5.C_ON=1'b0;
    defparam i20055_2_lut_LC_14_15_5.SEQ_MODE=4'b0000;
    defparam i20055_2_lut_LC_14_15_5.LUT_INIT=16'b0000000011001100;
    LogicCell40 i20055_2_lut_LC_14_15_5 (
            .in0(_gnd_net_),
            .in1(N__41806),
            .in2(_gnd_net_),
            .in3(N__59322),
            .lcout(n22301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i2_LC_14_16_0.C_ON=1'b0;
    defparam data_index_i2_LC_14_16_0.SEQ_MODE=4'b1000;
    defparam data_index_i2_LC_14_16_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i2_LC_14_16_0 (
            .in0(N__63735),
            .in1(N__41773),
            .in2(N__57778),
            .in3(N__41764),
            .lcout(data_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61917),
            .ce(),
            .sr(_gnd_net_));
    defparam i6641_3_lut_LC_14_16_1.C_ON=1'b0;
    defparam i6641_3_lut_LC_14_16_1.SEQ_MODE=4'b0000;
    defparam i6641_3_lut_LC_14_16_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6641_3_lut_LC_14_16_1 (
            .in0(N__52888),
            .in1(N__41791),
            .in2(_gnd_net_),
            .in3(N__56462),
            .lcout(n8_adj_1628),
            .ltout(n8_adj_1628_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_2_i15_4_lut_LC_14_16_2.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_2_i15_4_lut_LC_14_16_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_2_i15_4_lut_LC_14_16_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_358_Mux_2_i15_4_lut_LC_14_16_2 (
            .in0(N__57692),
            .in1(N__63618),
            .in2(N__41767),
            .in3(N__41763),
            .lcout(data_index_9_N_236_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i2_LC_14_16_3.C_ON=1'b0;
    defparam acadc_skipCount_i2_LC_14_16_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i2_LC_14_16_3.LUT_INIT=16'b0011000010111000;
    LogicCell40 acadc_skipCount_i2_LC_14_16_3 (
            .in0(N__52889),
            .in1(N__46818),
            .in2(N__52816),
            .in3(N__57700),
            .lcout(acadc_skipCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61917),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i3_LC_14_16_4.C_ON=1'b0;
    defparam data_index_i3_LC_14_16_4.SEQ_MODE=4'b1000;
    defparam data_index_i3_LC_14_16_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i3_LC_14_16_4 (
            .in0(N__63736),
            .in1(N__41653),
            .in2(N__57779),
            .in3(N__41640),
            .lcout(data_index_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61917),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_236_LC_14_16_5.C_ON=1'b0;
    defparam i10_4_lut_adj_236_LC_14_16_5.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_236_LC_14_16_5.LUT_INIT=16'b1111111111110110;
    LogicCell40 i10_4_lut_adj_236_LC_14_16_5 (
            .in0(N__41608),
            .in1(N__44105),
            .in2(N__41587),
            .in3(N__41575),
            .lcout(),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_241_LC_14_16_6.C_ON=1'b0;
    defparam i15_4_lut_adj_241_LC_14_16_6.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_241_LC_14_16_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_241_LC_14_16_6 (
            .in0(N__43972),
            .in1(N__41569),
            .in2(N__41560),
            .in3(N__41557),
            .lcout(n31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_321_LC_14_16_7.C_ON=1'b0;
    defparam i1_4_lut_adj_321_LC_14_16_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_321_LC_14_16_7.LUT_INIT=16'b1111000000010000;
    LogicCell40 i1_4_lut_adj_321_LC_14_16_7 (
            .in0(N__51380),
            .in1(N__46486),
            .in2(N__63723),
            .in3(N__57693),
            .lcout(n13141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_1_i16_3_lut_LC_14_17_0.C_ON=1'b0;
    defparam mux_126_Mux_1_i16_3_lut_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_1_i16_3_lut_LC_14_17_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_126_Mux_1_i16_3_lut_LC_14_17_0 (
            .in0(N__42154),
            .in1(N__42132),
            .in2(_gnd_net_),
            .in3(N__59442),
            .lcout(n16_adj_1751),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_2_i16_3_lut_LC_14_17_2.C_ON=1'b0;
    defparam mux_126_Mux_2_i16_3_lut_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_2_i16_3_lut_LC_14_17_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_126_Mux_2_i16_3_lut_LC_14_17_2 (
            .in0(N__42103),
            .in1(N__42350),
            .in2(_gnd_net_),
            .in3(N__59443),
            .lcout(),
            .ltout(n16_adj_1746_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19221_3_lut_LC_14_17_3.C_ON=1'b0;
    defparam i19221_3_lut_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam i19221_3_lut_LC_14_17_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 i19221_3_lut_LC_14_17_3 (
            .in0(_gnd_net_),
            .in1(N__42069),
            .in2(N__42034),
            .in3(N__60599),
            .lcout(n22148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.MISO_48_12606_12607_set_LC_14_17_4 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12606_12607_set_LC_14_17_4 .SEQ_MODE=4'b1011;
    defparam \comm_spi.MISO_48_12606_12607_set_LC_14_17_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.MISO_48_12606_12607_set_LC_14_17_4  (
            .in0(N__42031),
            .in1(N__42007),
            .in2(_gnd_net_),
            .in3(N__41985),
            .lcout(\comm_spi.n15334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12606_12607_setC_net ),
            .ce(),
            .sr(N__41913));
    defparam mux_125_Mux_1_i112_3_lut_LC_14_17_7.C_ON=1'b0;
    defparam mux_125_Mux_1_i112_3_lut_LC_14_17_7.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_1_i112_3_lut_LC_14_17_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_125_Mux_1_i112_3_lut_LC_14_17_7 (
            .in0(N__41872),
            .in1(N__41836),
            .in2(_gnd_net_),
            .in3(N__60598),
            .lcout(n112_adj_1799),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4594_3_lut_LC_14_18_0.C_ON=1'b0;
    defparam i4594_3_lut_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam i4594_3_lut_LC_14_18_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 i4594_3_lut_LC_14_18_0 (
            .in0(N__49129),
            .in1(N__47813),
            .in2(_gnd_net_),
            .in3(N__56458),
            .lcout(n8_adj_1605),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_207_LC_14_18_1.C_ON=1'b0;
    defparam i1_4_lut_adj_207_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_207_LC_14_18_1.LUT_INIT=16'b1101000011011101;
    LogicCell40 i1_4_lut_adj_207_LC_14_18_1 (
            .in0(N__41824),
            .in1(N__63194),
            .in2(N__63784),
            .in3(N__57703),
            .lcout(),
            .ltout(n12056_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds0_307_LC_14_18_2.C_ON=1'b0;
    defparam trig_dds0_307_LC_14_18_2.SEQ_MODE=4'b1000;
    defparam trig_dds0_307_LC_14_18_2.LUT_INIT=16'b0101110000001100;
    LogicCell40 trig_dds0_307_LC_14_18_2 (
            .in0(N__57705),
            .in1(N__47575),
            .in2(N__41809),
            .in3(N__63777),
            .lcout(trig_dds0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61953),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i4_4_lut_LC_14_18_4 .C_ON=1'b0;
    defparam \SIG_DDS.i4_4_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i4_4_lut_LC_14_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \SIG_DDS.i4_4_lut_LC_14_18_4  (
            .in0(N__47662),
            .in1(N__44737),
            .in2(N__44763),
            .in3(N__50614),
            .lcout(\SIG_DDS.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i23_LC_14_18_5.C_ON=1'b0;
    defparam comm_test_buf_24_i23_LC_14_18_5.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i23_LC_14_18_5.LUT_INIT=16'b0000101011001010;
    LogicCell40 comm_test_buf_24_i23_LC_14_18_5 (
            .in0(N__42372),
            .in1(N__46647),
            .in2(N__45427),
            .in3(N__57706),
            .lcout(comm_test_buf_24_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61953),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i2_LC_14_18_6.C_ON=1'b0;
    defparam buf_dds0_i2_LC_14_18_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i2_LC_14_18_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_dds0_i2_LC_14_18_6 (
            .in0(N__57704),
            .in1(N__50776),
            .in2(N__52925),
            .in3(N__42351),
            .lcout(buf_dds0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61953),
            .ce(),
            .sr(_gnd_net_));
    defparam i6591_3_lut_LC_14_18_7.C_ON=1'b0;
    defparam i6591_3_lut_LC_14_18_7.SEQ_MODE=4'b0000;
    defparam i6591_3_lut_LC_14_18_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 i6591_3_lut_LC_14_18_7 (
            .in0(N__56459),
            .in1(_gnd_net_),
            .in2(N__55837),
            .in3(N__44999),
            .lcout(n8_adj_1619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6571_3_lut_LC_14_19_5.C_ON=1'b0;
    defparam i6571_3_lut_LC_14_19_5.SEQ_MODE=4'b0000;
    defparam i6571_3_lut_LC_14_19_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6571_3_lut_LC_14_19_5 (
            .in0(N__44632),
            .in1(N__42334),
            .in2(_gnd_net_),
            .in3(N__56460),
            .lcout(n8_adj_1615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6581_3_lut_LC_14_19_6.C_ON=1'b0;
    defparam i6581_3_lut_LC_14_19_6.SEQ_MODE=4'b0000;
    defparam i6581_3_lut_LC_14_19_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 i6581_3_lut_LC_14_19_6 (
            .in0(N__56461),
            .in1(N__43947),
            .in2(_gnd_net_),
            .in3(N__44940),
            .lcout(n8_adj_1617),
            .ltout(n8_adj_1617_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_8_i15_4_lut_LC_14_19_7.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_8_i15_4_lut_LC_14_19_7.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_8_i15_4_lut_LC_14_19_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_358_Mux_8_i15_4_lut_LC_14_19_7 (
            .in0(N__57702),
            .in1(N__63724),
            .in2(N__42301),
            .in3(N__44970),
            .lcout(data_index_9_N_236_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i2_LC_14_20_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i2_LC_14_20_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i2_LC_14_20_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \SIG_DDS.dds_state_i2_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__50460),
            .in2(_gnd_net_),
            .in3(N__50364),
            .lcout(dds_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61983),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i20129_4_lut_LC_14_20_4 .C_ON=1'b0;
    defparam \SIG_DDS.i20129_4_lut_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i20129_4_lut_LC_14_20_4 .LUT_INIT=16'b1100110001000110;
    LogicCell40 \SIG_DDS.i20129_4_lut_LC_14_20_4  (
            .in0(N__50592),
            .in1(N__50459),
            .in2(N__47584),
            .in3(N__50363),
            .lcout(\SIG_DDS.n13338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_15_1_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_15_1_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_15_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_90_2_lut_LC_15_1_1  (
            .in0(N__42489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57118),
            .lcout(\comm_spi.iclk_N_850 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_12602_12603_reset_LC_15_2_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12602_12603_reset_LC_15_2_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imosi_44_12602_12603_reset_LC_15_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.imosi_44_12602_12603_reset_LC_15_2_0  (
            .in0(N__50200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n15331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61825),
            .ce(),
            .sr(N__44794));
    defparam \comm_spi.iclk_40_12598_12599_reset_LC_15_3_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12598_12599_reset_LC_15_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.iclk_40_12598_12599_reset_LC_15_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12598_12599_reset_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42490),
            .lcout(\comm_spi.n15327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61827),
            .ce(),
            .sr(N__42442));
    defparam \comm_spi.data_rx_i0_12616_12617_reset_LC_15_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12616_12617_reset_LC_15_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i0_12616_12617_reset_LC_15_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_12616_12617_reset_LC_15_4_0  (
            .in0(N__47959),
            .in1(N__44785),
            .in2(_gnd_net_),
            .in3(N__45459),
            .lcout(\comm_spi.n15345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53634),
            .ce(),
            .sr(N__42511));
    defparam \ADC_VDC.genclk.t_clk_24_LC_15_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t_clk_24_LC_15_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t_clk_24_LC_15_5_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \ADC_VDC.genclk.t_clk_24_LC_15_5_4  (
            .in0(_gnd_net_),
            .in1(N__64227),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(VDC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t_clk_24C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_1_i4_3_lut_LC_15_5_5.C_ON=1'b0;
    defparam mux_134_Mux_1_i4_3_lut_LC_15_5_5.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_1_i4_3_lut_LC_15_5_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_134_Mux_1_i4_3_lut_LC_15_5_5 (
            .in0(N__43333),
            .in1(N__54709),
            .in2(_gnd_net_),
            .in3(N__54409),
            .lcout(n4_adj_1676),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_15_5_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_15_5_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_87_2_lut_LC_15_5_6  (
            .in0(N__57121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47542),
            .lcout(\comm_spi.DOUT_7__N_835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_15_5_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_15_5_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_91_2_lut_LC_15_5_7  (
            .in0(N__42491),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57120),
            .lcout(\comm_spi.iclk_N_851 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_15_6_0.C_ON=1'b0;
    defparam i9_4_lut_LC_15_6_0.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_15_6_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_15_6_0 (
            .in0(N__42429),
            .in1(N__42417),
            .in2(N__42406),
            .in3(N__42390),
            .lcout(),
            .ltout(n25_adj_1717_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_205_LC_15_6_1.C_ON=1'b0;
    defparam i15_4_lut_adj_205_LC_15_6_1.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_205_LC_15_6_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_205_LC_15_6_1 (
            .in0(N__45154),
            .in1(N__42853),
            .in2(N__42379),
            .in3(N__42910),
            .lcout(),
            .ltout(n20922_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_15_6_2.C_ON=1'b0;
    defparam i7_4_lut_LC_15_6_2.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_15_6_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 i7_4_lut_LC_15_6_2 (
            .in0(N__42967),
            .in1(N__43017),
            .in2(N__43006),
            .in3(N__43003),
            .lcout(n15420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_15_6_3.C_ON=1'b0;
    defparam i2_2_lut_LC_15_6_3.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_15_6_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2_2_lut_LC_15_6_3 (
            .in0(_gnd_net_),
            .in1(N__42993),
            .in2(_gnd_net_),
            .in3(N__42982),
            .lcout(n10_adj_1679),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_203_LC_15_6_4.C_ON=1'b0;
    defparam i11_4_lut_adj_203_LC_15_6_4.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_203_LC_15_6_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_203_LC_15_6_4 (
            .in0(N__42960),
            .in1(N__42948),
            .in2(N__42937),
            .in3(N__42921),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_15_6_5.C_ON=1'b0;
    defparam i10_4_lut_LC_15_6_5.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_15_6_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_LC_15_6_5 (
            .in0(N__42903),
            .in1(N__42891),
            .in2(N__42880),
            .in3(N__42864),
            .lcout(n26_adj_1715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SecClk_295_LC_15_7_2.C_ON=1'b0;
    defparam SecClk_295_LC_15_7_2.SEQ_MODE=4'b1000;
    defparam SecClk_295_LC_15_7_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 SecClk_295_LC_15_7_2 (
            .in0(_gnd_net_),
            .in1(N__42792),
            .in2(_gnd_net_),
            .in3(N__42826),
            .lcout(TEST_LED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_374_i9_2_lut_3_lut_LC_15_7_3.C_ON=1'b0;
    defparam comm_cmd_6__I_0_374_i9_2_lut_3_lut_LC_15_7_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_374_i9_2_lut_3_lut_LC_15_7_3.LUT_INIT=16'b1111111111101110;
    LogicCell40 comm_cmd_6__I_0_374_i9_2_lut_3_lut_LC_15_7_3 (
            .in0(N__59189),
            .in1(N__59969),
            .in2(_gnd_net_),
            .in3(N__60498),
            .lcout(n9_adj_1596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9640_1_lut_LC_15_7_4.C_ON=1'b0;
    defparam i9640_1_lut_LC_15_7_4.SEQ_MODE=4'b0000;
    defparam i9640_1_lut_LC_15_7_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i9640_1_lut_LC_15_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52658),
            .lcout(n12366),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19311_3_lut_LC_15_7_5.C_ON=1'b0;
    defparam i19311_3_lut_LC_15_7_5.SEQ_MODE=4'b0000;
    defparam i19311_3_lut_LC_15_7_5.LUT_INIT=16'b1100110010111011;
    LogicCell40 i19311_3_lut_LC_15_7_5 (
            .in0(N__58204),
            .in1(N__62637),
            .in2(_gnd_net_),
            .in3(N__63082),
            .lcout(n22238),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i7_LC_15_8_0.C_ON=1'b0;
    defparam comm_buf_6__i7_LC_15_8_0.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i7_LC_15_8_0.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i7_LC_15_8_0 (
            .in0(N__43072),
            .in1(N__63487),
            .in2(N__55941),
            .in3(N__45558),
            .lcout(comm_buf_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61843),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_test_buf_24_i17_LC_15_8_1.C_ON=1'b0;
    defparam comm_test_buf_24_i17_LC_15_8_1.SEQ_MODE=4'b1000;
    defparam comm_test_buf_24_i17_LC_15_8_1.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_test_buf_24_i17_LC_15_8_1 (
            .in0(N__57520),
            .in1(N__43056),
            .in2(N__44631),
            .in3(N__45372),
            .lcout(comm_test_buf_24_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61843),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i7_LC_15_8_3.C_ON=1'b0;
    defparam comm_cmd_i7_LC_15_8_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i7_LC_15_8_3.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i7_LC_15_8_3 (
            .in0(N__51165),
            .in1(N__55935),
            .in2(N__45955),
            .in3(N__45977),
            .lcout(comm_cmd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61843),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i0_LC_15_8_4.C_ON=1'b0;
    defparam comm_buf_6__i0_LC_15_8_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i0_LC_15_8_4.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_buf_6__i0_LC_15_8_4 (
            .in0(N__63489),
            .in1(N__53990),
            .in2(N__43042),
            .in3(N__45557),
            .lcout(comm_buf_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61843),
            .ce(),
            .sr(_gnd_net_));
    defparam i12808_3_lut_LC_15_8_6.C_ON=1'b0;
    defparam i12808_3_lut_LC_15_8_6.SEQ_MODE=4'b0000;
    defparam i12808_3_lut_LC_15_8_6.LUT_INIT=16'b1000100010101010;
    LogicCell40 i12808_3_lut_LC_15_8_6 (
            .in0(N__46390),
            .in1(N__63486),
            .in2(_gnd_net_),
            .in3(N__51164),
            .lcout(n15531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i5_LC_15_8_7.C_ON=1'b0;
    defparam comm_buf_6__i5_LC_15_8_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i5_LC_15_8_7.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_buf_6__i5_LC_15_8_7 (
            .in0(N__45556),
            .in1(N__45714),
            .in2(N__55193),
            .in3(N__63490),
            .lcout(comm_buf_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61843),
            .ce(),
            .sr(_gnd_net_));
    defparam i16114_3_lut_LC_15_9_0.C_ON=1'b0;
    defparam i16114_3_lut_LC_15_9_0.SEQ_MODE=4'b0000;
    defparam i16114_3_lut_LC_15_9_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i16114_3_lut_LC_15_9_0 (
            .in0(N__43041),
            .in1(N__43226),
            .in2(_gnd_net_),
            .in3(N__54588),
            .lcout(n18816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16116_3_lut_LC_15_9_1.C_ON=1'b0;
    defparam i16116_3_lut_LC_15_9_1.SEQ_MODE=4'b0000;
    defparam i16116_3_lut_LC_15_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i16116_3_lut_LC_15_9_1 (
            .in0(N__54587),
            .in1(N__43171),
            .in2(_gnd_net_),
            .in3(N__49122),
            .lcout(),
            .ltout(n18818_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_20434_LC_15_9_2.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_20434_LC_15_9_2.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_20434_LC_15_9_2.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_index_1__bdd_4_lut_20434_LC_15_9_2 (
            .in0(N__43240),
            .in1(N__54362),
            .in2(N__43024),
            .in3(N__51821),
            .lcout(),
            .ltout(n23372_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i0_LC_15_9_3.C_ON=1'b0;
    defparam comm_tx_buf_i0_LC_15_9_3.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i0_LC_15_9_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 comm_tx_buf_i0_LC_15_9_3 (
            .in0(N__54363),
            .in1(N__43234),
            .in2(N__43021),
            .in3(N__43294),
            .lcout(comm_tx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61849),
            .ce(N__46404),
            .sr(N__46352));
    defparam i19938_2_lut_LC_15_9_4.C_ON=1'b0;
    defparam i19938_2_lut_LC_15_9_4.SEQ_MODE=4'b0000;
    defparam i19938_2_lut_LC_15_9_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19938_2_lut_LC_15_9_4 (
            .in0(_gnd_net_),
            .in1(N__43249),
            .in2(_gnd_net_),
            .in3(N__54586),
            .lcout(n22338),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16113_3_lut_LC_15_9_5.C_ON=1'b0;
    defparam i16113_3_lut_LC_15_9_5.SEQ_MODE=4'b0000;
    defparam i16113_3_lut_LC_15_9_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 i16113_3_lut_LC_15_9_5 (
            .in0(N__54589),
            .in1(_gnd_net_),
            .in2(N__43956),
            .in3(N__53938),
            .lcout(n18815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16121_3_lut_LC_15_9_6.C_ON=1'b0;
    defparam i16121_3_lut_LC_15_9_6.SEQ_MODE=4'b0000;
    defparam i16121_3_lut_LC_15_9_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i16121_3_lut_LC_15_9_6 (
            .in0(N__43227),
            .in1(N__43948),
            .in2(_gnd_net_),
            .in3(N__46201),
            .lcout(n18823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_5__i0_LC_15_10_0.C_ON=1'b0;
    defparam comm_buf_5__i0_LC_15_10_0.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i0_LC_15_10_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_5__i0_LC_15_10_0 (
            .in0(N__43186),
            .in1(N__62629),
            .in2(_gnd_net_),
            .in3(N__54015),
            .lcout(comm_buf_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_buf_5__i7_LC_15_10_1.C_ON=1'b0;
    defparam comm_buf_5__i7_LC_15_10_1.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i7_LC_15_10_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_5__i7_LC_15_10_1 (
            .in0(N__62628),
            .in1(_gnd_net_),
            .in2(N__55931),
            .in3(N__43165),
            .lcout(comm_buf_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_buf_5__i6_LC_15_10_2.C_ON=1'b0;
    defparam comm_buf_5__i6_LC_15_10_2.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i6_LC_15_10_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i6_LC_15_10_2 (
            .in0(N__53856),
            .in1(N__43141),
            .in2(_gnd_net_),
            .in3(N__62632),
            .lcout(comm_buf_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_buf_5__i5_LC_15_10_3.C_ON=1'b0;
    defparam comm_buf_5__i5_LC_15_10_3.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i5_LC_15_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i5_LC_15_10_3 (
            .in0(N__62627),
            .in1(N__55160),
            .in2(_gnd_net_),
            .in3(N__43114),
            .lcout(comm_buf_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_buf_5__i4_LC_15_10_4.C_ON=1'b0;
    defparam comm_buf_5__i4_LC_15_10_4.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i4_LC_15_10_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i4_LC_15_10_4 (
            .in0(N__55067),
            .in1(N__43099),
            .in2(_gnd_net_),
            .in3(N__62631),
            .lcout(comm_buf_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_buf_5__i3_LC_15_10_5.C_ON=1'b0;
    defparam comm_buf_5__i3_LC_15_10_5.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i3_LC_15_10_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_5__i3_LC_15_10_5 (
            .in0(N__62626),
            .in1(_gnd_net_),
            .in2(N__62779),
            .in3(N__43387),
            .lcout(comm_buf_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_buf_5__i2_LC_15_10_6.C_ON=1'b0;
    defparam comm_buf_5__i2_LC_15_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i2_LC_15_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i2_LC_15_10_6 (
            .in0(N__54931),
            .in1(N__43369),
            .in2(_gnd_net_),
            .in3(N__62630),
            .lcout(comm_buf_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_buf_5__i1_LC_15_10_7.C_ON=1'b0;
    defparam comm_buf_5__i1_LC_15_10_7.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i1_LC_15_10_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i1_LC_15_10_7 (
            .in0(N__62625),
            .in1(N__54788),
            .in2(_gnd_net_),
            .in3(N__43348),
            .lcout(comm_buf_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61856),
            .ce(N__45886),
            .sr(N__45736));
    defparam comm_cmd_i0_LC_15_11_0.C_ON=1'b0;
    defparam comm_cmd_i0_LC_15_11_0.SEQ_MODE=4'b1000;
    defparam comm_cmd_i0_LC_15_11_0.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i0_LC_15_11_0 (
            .in0(N__58844),
            .in1(N__54020),
            .in2(N__45953),
            .in3(N__45996),
            .lcout(comm_cmd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61864),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i2_LC_15_11_1.C_ON=1'b0;
    defparam comm_cmd_i2_LC_15_11_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i2_LC_15_11_1.LUT_INIT=16'b1110001000100010;
    LogicCell40 comm_cmd_i2_LC_15_11_1 (
            .in0(N__59703),
            .in1(N__45998),
            .in2(N__45954),
            .in3(N__54930),
            .lcout(comm_cmd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61864),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i3_LC_15_11_2.C_ON=1'b0;
    defparam comm_cmd_i3_LC_15_11_2.SEQ_MODE=4'b1000;
    defparam comm_cmd_i3_LC_15_11_2.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i3_LC_15_11_2 (
            .in0(N__45942),
            .in1(N__45997),
            .in2(N__62794),
            .in3(N__60865),
            .lcout(comm_cmd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61864),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_188_i9_2_lut_3_lut_LC_15_11_3.C_ON=1'b0;
    defparam equal_188_i9_2_lut_3_lut_LC_15_11_3.SEQ_MODE=4'b0000;
    defparam equal_188_i9_2_lut_3_lut_LC_15_11_3.LUT_INIT=16'b1110111011111111;
    LogicCell40 equal_188_i9_2_lut_3_lut_LC_15_11_3 (
            .in0(N__59702),
            .in1(N__60248),
            .in2(_gnd_net_),
            .in3(N__58842),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_60_LC_15_11_4.C_ON=1'b0;
    defparam i1_2_lut_adj_60_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_60_LC_15_11_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_adj_60_LC_15_11_4 (
            .in0(N__61231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58614),
            .lcout(n8_adj_1504),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_20553_LC_15_11_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_20553_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_20553_LC_15_11_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_20553_LC_15_11_5 (
            .in0(N__48706),
            .in1(N__60249),
            .in2(N__43321),
            .in3(N__58843),
            .lcout(),
            .ltout(n23504_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23504_bdd_4_lut_LC_15_11_6.C_ON=1'b0;
    defparam n23504_bdd_4_lut_LC_15_11_6.SEQ_MODE=4'b0000;
    defparam n23504_bdd_4_lut_LC_15_11_6.LUT_INIT=16'b1110010111100000;
    LogicCell40 n23504_bdd_4_lut_LC_15_11_6 (
            .in0(N__60250),
            .in1(N__43543),
            .in2(N__43519),
            .in3(N__43509),
            .lcout(n22288),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i1_LC_15_11_7.C_ON=1'b0;
    defparam buf_control_i1_LC_15_11_7.SEQ_MODE=4'b1000;
    defparam buf_control_i1_LC_15_11_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i1_LC_15_11_7 (
            .in0(N__57620),
            .in1(N__46749),
            .in2(N__44617),
            .in3(N__49866),
            .lcout(DDS_RNG_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61864),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_315_LC_15_12_0.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_315_LC_15_12_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_315_LC_15_12_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_3_lut_4_lut_adj_315_LC_15_12_0 (
            .in0(N__63045),
            .in1(N__61300),
            .in2(N__43650),
            .in3(N__58608),
            .lcout(n21964),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_309_LC_15_12_1.C_ON=1'b0;
    defparam i1_4_lut_adj_309_LC_15_12_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_309_LC_15_12_1.LUT_INIT=16'b1010001010100000;
    LogicCell40 i1_4_lut_adj_309_LC_15_12_1 (
            .in0(N__54081),
            .in1(N__63046),
            .in2(N__54161),
            .in3(N__45865),
            .lcout(n12838),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20382_LC_15_12_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20382_LC_15_12_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20382_LC_15_12_2.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_20382_LC_15_12_2 (
            .in0(N__45829),
            .in1(N__60262),
            .in2(N__49012),
            .in3(N__59812),
            .lcout(n23306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19135_2_lut_3_lut_LC_15_12_3.C_ON=1'b0;
    defparam i19135_2_lut_3_lut_LC_15_12_3.SEQ_MODE=4'b0000;
    defparam i19135_2_lut_3_lut_LC_15_12_3.LUT_INIT=16'b1111111111101110;
    LogicCell40 i19135_2_lut_3_lut_LC_15_12_3 (
            .in0(N__58609),
            .in1(N__58365),
            .in2(_gnd_net_),
            .in3(N__61232),
            .lcout(n22061),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i4_LC_15_12_4.C_ON=1'b0;
    defparam comm_cmd_i4_LC_15_12_4.SEQ_MODE=4'b1000;
    defparam comm_cmd_i4_LC_15_12_4.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i4_LC_15_12_4 (
            .in0(N__58483),
            .in1(N__45941),
            .in2(N__55081),
            .in3(N__46008),
            .lcout(comm_cmd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61876),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_374_i10_2_lut_LC_15_12_5.C_ON=1'b0;
    defparam comm_cmd_6__I_0_374_i10_2_lut_LC_15_12_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_374_i10_2_lut_LC_15_12_5.LUT_INIT=16'b1111111100110011;
    LogicCell40 comm_cmd_6__I_0_374_i10_2_lut_LC_15_12_5 (
            .in0(_gnd_net_),
            .in1(N__58482),
            .in2(_gnd_net_),
            .in3(N__60879),
            .lcout(n6),
            .ltout(n6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_62_LC_15_12_6.C_ON=1'b0;
    defparam i1_4_lut_adj_62_LC_15_12_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_62_LC_15_12_6.LUT_INIT=16'b0000001100001011;
    LogicCell40 i1_4_lut_adj_62_LC_15_12_6 (
            .in0(N__43435),
            .in1(N__43633),
            .in2(N__43426),
            .in3(N__46481),
            .lcout(n21938),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i5_LC_15_12_7.C_ON=1'b0;
    defparam comm_cmd_i5_LC_15_12_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i5_LC_15_12_7.LUT_INIT=16'b1010110000001100;
    LogicCell40 comm_cmd_i5_LC_15_12_7 (
            .in0(N__45940),
            .in1(N__58615),
            .in2(N__46012),
            .in3(N__55189),
            .lcout(comm_cmd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61876),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20372_LC_15_13_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20372_LC_15_13_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20372_LC_15_13_1.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20372_LC_15_13_1 (
            .in0(N__59822),
            .in1(N__43699),
            .in2(N__43687),
            .in3(N__60353),
            .lcout(n23288),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i5_LC_15_13_2.C_ON=1'b0;
    defparam acadc_skipCount_i5_LC_15_13_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i5_LC_15_13_2.LUT_INIT=16'b0111001001010000;
    LogicCell40 acadc_skipCount_i5_LC_15_13_2 (
            .in0(N__46849),
            .in1(N__57619),
            .in2(N__51925),
            .in3(N__56577),
            .lcout(acadc_skipCount_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61888),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i1_LC_15_13_3.C_ON=1'b0;
    defparam acadc_skipCount_i1_LC_15_13_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i1_LC_15_13_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i1_LC_15_13_3 (
            .in0(N__57618),
            .in1(N__46850),
            .in2(N__52142),
            .in3(N__52233),
            .lcout(acadc_skipCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61888),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i2_LC_15_13_4.C_ON=1'b0;
    defparam req_data_cnt_i2_LC_15_13_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i2_LC_15_13_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 req_data_cnt_i2_LC_15_13_4 (
            .in0(N__51362),
            .in1(_gnd_net_),
            .in2(N__52842),
            .in3(N__47154),
            .lcout(req_data_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61888),
            .ce(),
            .sr(_gnd_net_));
    defparam i19814_3_lut_4_lut_LC_15_13_5.C_ON=1'b0;
    defparam i19814_3_lut_4_lut_LC_15_13_5.SEQ_MODE=4'b0000;
    defparam i19814_3_lut_4_lut_LC_15_13_5.LUT_INIT=16'b0000000000010000;
    LogicCell40 i19814_3_lut_4_lut_LC_15_13_5 (
            .in0(N__61267),
            .in1(N__60880),
            .in2(N__59973),
            .in3(N__58607),
            .lcout(),
            .ltout(n22396_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19906_4_lut_LC_15_13_6.C_ON=1'b0;
    defparam i19906_4_lut_LC_15_13_6.SEQ_MODE=4'b0000;
    defparam i19906_4_lut_LC_15_13_6.LUT_INIT=16'b1101100000000000;
    LogicCell40 i19906_4_lut_LC_15_13_6 (
            .in0(N__60352),
            .in1(N__56170),
            .in2(N__43654),
            .in3(N__58487),
            .lcout(n22397),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_56_LC_15_13_7.C_ON=1'b0;
    defparam i1_4_lut_adj_56_LC_15_13_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_56_LC_15_13_7.LUT_INIT=16'b0000001000001111;
    LogicCell40 i1_4_lut_adj_56_LC_15_13_7 (
            .in0(N__61268),
            .in1(N__46453),
            .in2(N__43651),
            .in3(N__43632),
            .lcout(n21929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_250_LC_15_14_0.C_ON=1'b0;
    defparam i6_4_lut_adj_250_LC_15_14_0.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_250_LC_15_14_0.LUT_INIT=16'b0110111111110110;
    LogicCell40 i6_4_lut_adj_250_LC_15_14_0 (
            .in0(N__55490),
            .in1(N__54658),
            .in2(N__52405),
            .in3(N__52832),
            .lcout(n22_adj_1801),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_1_i127_3_lut_LC_15_14_1.C_ON=1'b0;
    defparam mux_125_Mux_1_i127_3_lut_LC_15_14_1.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_1_i127_3_lut_LC_15_14_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_125_Mux_1_i127_3_lut_LC_15_14_1 (
            .in0(N__43567),
            .in1(N__61291),
            .in2(_gnd_net_),
            .in3(N__50965),
            .lcout(comm_buf_0_7_N_543_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_255_LC_15_14_2.C_ON=1'b0;
    defparam i2_4_lut_adj_255_LC_15_14_2.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_255_LC_15_14_2.LUT_INIT=16'b0110111111110110;
    LogicCell40 i2_4_lut_adj_255_LC_15_14_2 (
            .in0(N__52482),
            .in1(N__52549),
            .in2(N__52206),
            .in3(N__52258),
            .lcout(n18_adj_1699),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i1_LC_15_14_3.C_ON=1'b0;
    defparam req_data_cnt_i1_LC_15_14_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i1_LC_15_14_3.LUT_INIT=16'b1100101011001010;
    LogicCell40 req_data_cnt_i1_LC_15_14_3 (
            .in0(N__52205),
            .in1(N__47185),
            .in2(N__51338),
            .in3(_gnd_net_),
            .lcout(req_data_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61904),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_302_LC_15_14_5.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_302_LC_15_14_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_302_LC_15_14_5.LUT_INIT=16'b1111000000100000;
    LogicCell40 i1_3_lut_4_lut_adj_302_LC_15_14_5 (
            .in0(N__46203),
            .in1(N__63051),
            .in2(N__63762),
            .in3(N__57610),
            .lcout(n13257),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i7_LC_15_14_6.C_ON=1'b0;
    defparam req_data_cnt_i7_LC_15_14_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i7_LC_15_14_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 req_data_cnt_i7_LC_15_14_6 (
            .in0(_gnd_net_),
            .in1(N__47515),
            .in2(N__55497),
            .in3(N__51310),
            .lcout(req_data_cnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61904),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_235_LC_15_14_7.C_ON=1'b0;
    defparam i2_4_lut_adj_235_LC_15_14_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_235_LC_15_14_7.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_235_LC_15_14_7 (
            .in0(N__44017),
            .in1(N__52505),
            .in2(N__43996),
            .in3(N__52229),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_start_332_LC_15_15_0.C_ON=1'b0;
    defparam eis_start_332_LC_15_15_0.SEQ_MODE=4'b1000;
    defparam eis_start_332_LC_15_15_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_start_332_LC_15_15_0 (
            .in0(N__43960),
            .in1(N__43873),
            .in2(_gnd_net_),
            .in3(N__43828),
            .lcout(eis_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61918),
            .ce(),
            .sr(_gnd_net_));
    defparam i6621_3_lut_LC_15_15_1.C_ON=1'b0;
    defparam i6621_3_lut_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam i6621_3_lut_LC_15_15_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6621_3_lut_LC_15_15_1 (
            .in0(N__56065),
            .in1(N__44156),
            .in2(_gnd_net_),
            .in3(N__56451),
            .lcout(n8_adj_1625),
            .ltout(n8_adj_1625_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_4_i15_4_lut_LC_15_15_2.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_4_i15_4_lut_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_4_i15_4_lut_LC_15_15_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_state_3__I_0_358_Mux_4_i15_4_lut_LC_15_15_2 (
            .in0(N__63654),
            .in1(N__57582),
            .in2(N__43798),
            .in3(N__44181),
            .lcout(data_index_9_N_236_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i15_LC_15_15_3.C_ON=1'b0;
    defparam req_data_cnt_i15_LC_15_15_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i15_LC_15_15_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 req_data_cnt_i15_LC_15_15_3 (
            .in0(N__57583),
            .in1(N__51339),
            .in2(N__46658),
            .in3(N__44383),
            .lcout(req_data_cnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61918),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i0_LC_15_15_4.C_ON=1'b0;
    defparam req_data_cnt_i0_LC_15_15_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i0_LC_15_15_4.LUT_INIT=16'b0010001011100010;
    LogicCell40 req_data_cnt_i0_LC_15_15_4 (
            .in0(N__47014),
            .in1(N__51323),
            .in2(N__49133),
            .in3(N__57587),
            .lcout(req_data_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61918),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i4_LC_15_15_5.C_ON=1'b0;
    defparam data_index_i4_LC_15_15_5.SEQ_MODE=4'b1000;
    defparam data_index_i4_LC_15_15_5.LUT_INIT=16'b0000110010101010;
    LogicCell40 data_index_i4_LC_15_15_5 (
            .in0(N__44182),
            .in1(N__44170),
            .in2(N__57701),
            .in3(N__63655),
            .lcout(data_index_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61918),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20577_LC_15_15_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20577_LC_15_15_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20577_LC_15_15_6.LUT_INIT=16'b1110011011000100;
    LogicCell40 comm_cmd_1__bdd_4_lut_20577_LC_15_15_6 (
            .in0(N__59961),
            .in1(N__60478),
            .in2(N__56917),
            .in3(N__44350),
            .lcout(n23546),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_124_Mux_0_i30_4_lut_4_lut_LC_15_15_7.C_ON=1'b0;
    defparam mux_124_Mux_0_i30_4_lut_4_lut_LC_15_15_7.SEQ_MODE=4'b0000;
    defparam mux_124_Mux_0_i30_4_lut_4_lut_LC_15_15_7.LUT_INIT=16'b0000011110011010;
    LogicCell40 mux_124_Mux_0_i30_4_lut_4_lut_LC_15_15_7 (
            .in0(N__60479),
            .in1(N__59227),
            .in2(N__61018),
            .in3(N__59962),
            .lcout(n30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_259_LC_15_16_0.C_ON=1'b0;
    defparam i1_4_lut_adj_259_LC_15_16_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_259_LC_15_16_0.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_259_LC_15_16_0 (
            .in0(N__49396),
            .in1(N__49655),
            .in2(N__47013),
            .in3(N__49786),
            .lcout(n17_adj_1594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i6_LC_15_16_1.C_ON=1'b0;
    defparam req_data_cnt_i6_LC_15_16_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i6_LC_15_16_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 req_data_cnt_i6_LC_15_16_1 (
            .in0(N__49656),
            .in1(_gnd_net_),
            .in2(N__47076),
            .in3(N__51363),
            .lcout(req_data_cnt_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61938),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i8_LC_15_16_2.C_ON=1'b0;
    defparam acadc_skipCount_i8_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i8_LC_15_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_skipCount_i8_LC_15_16_2 (
            .in0(N__48872),
            .in1(N__46817),
            .in2(_gnd_net_),
            .in3(N__44115),
            .lcout(acadc_skipCount_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61938),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_249_LC_15_16_4.C_ON=1'b0;
    defparam i8_4_lut_adj_249_LC_15_16_4.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_249_LC_15_16_4.LUT_INIT=16'b0110111111110110;
    LogicCell40 i8_4_lut_adj_249_LC_15_16_4 (
            .in0(N__44381),
            .in1(N__50035),
            .in2(N__44079),
            .in3(N__50938),
            .lcout(n24_adj_1800),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i9_LC_15_16_5.C_ON=1'b0;
    defparam req_data_cnt_i9_LC_15_16_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i9_LC_15_16_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 req_data_cnt_i9_LC_15_16_5 (
            .in0(N__44078),
            .in1(N__51364),
            .in2(_gnd_net_),
            .in3(N__50808),
            .lcout(req_data_cnt_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61938),
            .ce(),
            .sr(_gnd_net_));
    defparam i20048_2_lut_LC_15_16_6.C_ON=1'b0;
    defparam i20048_2_lut_LC_15_16_6.SEQ_MODE=4'b0000;
    defparam i20048_2_lut_LC_15_16_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 i20048_2_lut_LC_15_16_6 (
            .in0(N__59010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44382),
            .lcout(n22314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19242_3_lut_LC_15_16_7.C_ON=1'b0;
    defparam i19242_3_lut_LC_15_16_7.SEQ_MODE=4'b0000;
    defparam i19242_3_lut_LC_15_16_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 i19242_3_lut_LC_15_16_7 (
            .in0(N__47391),
            .in1(_gnd_net_),
            .in2(N__50127),
            .in3(N__59009),
            .lcout(n22169),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20387_LC_15_17_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20387_LC_15_17_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20387_LC_15_17_0.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_20387_LC_15_17_0 (
            .in0(N__60496),
            .in1(N__59536),
            .in2(N__46447),
            .in3(N__59963),
            .lcout(),
            .ltout(n23312_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23312_bdd_4_lut_LC_15_17_1.C_ON=1'b0;
    defparam n23312_bdd_4_lut_LC_15_17_1.SEQ_MODE=4'b0000;
    defparam n23312_bdd_4_lut_LC_15_17_1.LUT_INIT=16'b1110010111100000;
    LogicCell40 n23312_bdd_4_lut_LC_15_17_1 (
            .in0(N__59965),
            .in1(N__44344),
            .in2(N__44320),
            .in3(N__44288),
            .lcout(),
            .ltout(n23315_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1665080_i1_3_lut_LC_15_17_2.C_ON=1'b0;
    defparam i1665080_i1_3_lut_LC_15_17_2.SEQ_MODE=4'b0000;
    defparam i1665080_i1_3_lut_LC_15_17_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1665080_i1_3_lut_LC_15_17_2 (
            .in0(_gnd_net_),
            .in1(N__44188),
            .in2(N__44317),
            .in3(N__60948),
            .lcout(),
            .ltout(n30_adj_1741_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_3_i127_3_lut_LC_15_17_3.C_ON=1'b0;
    defparam mux_126_Mux_3_i127_3_lut_LC_15_17_3.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_3_i127_3_lut_LC_15_17_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_126_Mux_3_i127_3_lut_LC_15_17_3 (
            .in0(_gnd_net_),
            .in1(N__44314),
            .in2(N__44299),
            .in3(N__61373),
            .lcout(comm_buf_1_7_N_559_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i3_LC_15_17_4.C_ON=1'b0;
    defparam acadc_skipCount_i3_LC_15_17_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i3_LC_15_17_4.LUT_INIT=16'b0100010011110000;
    LogicCell40 acadc_skipCount_i3_LC_15_17_4 (
            .in0(N__57617),
            .in1(N__49330),
            .in2(N__44295),
            .in3(N__46820),
            .lcout(acadc_skipCount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61954),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_LC_15_17_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_LC_15_17_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_LC_15_17_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_LC_15_17_5 (
            .in0(N__44272),
            .in1(N__59960),
            .in2(N__44260),
            .in3(N__60495),
            .lcout(),
            .ltout(n23558_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23558_bdd_4_lut_LC_15_17_6.C_ON=1'b0;
    defparam n23558_bdd_4_lut_LC_15_17_6.SEQ_MODE=4'b0000;
    defparam n23558_bdd_4_lut_LC_15_17_6.LUT_INIT=16'b1111000010101100;
    LogicCell40 n23558_bdd_4_lut_LC_15_17_6 (
            .in0(N__44230),
            .in1(N__44203),
            .in2(N__44191),
            .in3(N__59964),
            .lcout(n23561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i3_LC_15_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i3_LC_15_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i3_LC_15_18_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \SIG_DDS.bit_cnt_i3_LC_15_18_0  (
            .in0(N__44742),
            .in1(N__47661),
            .in2(N__44764),
            .in3(N__44527),
            .lcout(\SIG_DDS.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61971),
            .ce(N__50404),
            .sr(N__47674));
    defparam \SIG_DDS.bit_cnt_i2_LC_15_18_1 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i2_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i2_LC_15_18_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \SIG_DDS.bit_cnt_i2_LC_15_18_1  (
            .in0(N__47660),
            .in1(_gnd_net_),
            .in2(N__44743),
            .in3(N__44759),
            .lcout(\SIG_DDS.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61971),
            .ce(N__50404),
            .sr(N__47674));
    defparam \SIG_DDS.bit_cnt_i1_LC_15_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i1_LC_15_18_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i1_LC_15_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \SIG_DDS.bit_cnt_i1_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__44738),
            .in2(_gnd_net_),
            .in3(N__47659),
            .lcout(\SIG_DDS.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61971),
            .ce(N__50404),
            .sr(N__47674));
    defparam i16455_2_lut_3_lut_LC_15_18_3.C_ON=1'b0;
    defparam i16455_2_lut_3_lut_LC_15_18_3.SEQ_MODE=4'b0000;
    defparam i16455_2_lut_3_lut_LC_15_18_3.LUT_INIT=16'b0000000000100010;
    LogicCell40 i16455_2_lut_3_lut_LC_15_18_3 (
            .in0(N__44715),
            .in1(N__62678),
            .in2(_gnd_net_),
            .in3(N__64076),
            .lcout(n14_adj_1653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16463_2_lut_3_lut_LC_15_18_4.C_ON=1'b0;
    defparam i16463_2_lut_3_lut_LC_15_18_4.SEQ_MODE=4'b0000;
    defparam i16463_2_lut_3_lut_LC_15_18_4.LUT_INIT=16'b0000010000000100;
    LogicCell40 i16463_2_lut_3_lut_LC_15_18_4 (
            .in0(N__64077),
            .in1(N__55827),
            .in2(N__62690),
            .in3(_gnd_net_),
            .lcout(n14_adj_1609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16458_2_lut_3_lut_LC_15_18_6.C_ON=1'b0;
    defparam i16458_2_lut_3_lut_LC_15_18_6.SEQ_MODE=4'b0000;
    defparam i16458_2_lut_3_lut_LC_15_18_6.LUT_INIT=16'b0000010000000100;
    LogicCell40 i16458_2_lut_3_lut_LC_15_18_6 (
            .in0(N__64078),
            .in1(N__44642),
            .in2(N__62691),
            .in3(_gnd_net_),
            .lcout(n14_adj_1656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i6_LC_15_19_0.C_ON=1'b0;
    defparam data_index_i6_LC_15_19_0.SEQ_MODE=4'b1000;
    defparam data_index_i6_LC_15_19_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i6_LC_15_19_0 (
            .in0(N__45121),
            .in1(N__63742),
            .in2(N__57708),
            .in3(N__45112),
            .lcout(data_index_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61984),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19893_2_lut_LC_15_19_1 .C_ON=1'b0;
    defparam \SIG_DDS.i19893_2_lut_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19893_2_lut_LC_15_19_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \SIG_DDS.i19893_2_lut_LC_15_19_1  (
            .in0(N__44526),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50455),
            .lcout(\SIG_DDS.n22671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_9_i15_4_lut_LC_15_19_2.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_9_i15_4_lut_LC_15_19_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_9_i15_4_lut_LC_15_19_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_358_Mux_9_i15_4_lut_LC_15_19_2 (
            .in0(N__63738),
            .in1(N__44508),
            .in2(N__57707),
            .in3(N__44496),
            .lcout(data_index_9_N_236_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6601_3_lut_LC_15_19_3.C_ON=1'b0;
    defparam i6601_3_lut_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam i6601_3_lut_LC_15_19_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6601_3_lut_LC_15_19_3 (
            .in0(N__49221),
            .in1(N__45135),
            .in2(_gnd_net_),
            .in3(N__56473),
            .lcout(n8_adj_1621),
            .ltout(n8_adj_1621_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_6_i15_4_lut_LC_15_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_6_i15_4_lut_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_6_i15_4_lut_LC_15_19_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_358_Mux_6_i15_4_lut_LC_15_19_4 (
            .in0(N__57603),
            .in1(N__63740),
            .in2(N__45115),
            .in3(N__45111),
            .lcout(data_index_9_N_236_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i7_LC_15_19_5.C_ON=1'b0;
    defparam data_index_i7_LC_15_19_5.SEQ_MODE=4'b1000;
    defparam data_index_i7_LC_15_19_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i7_LC_15_19_5 (
            .in0(N__63741),
            .in1(N__44926),
            .in2(N__57711),
            .in3(N__44917),
            .lcout(data_index_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61984),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i8_LC_15_19_6.C_ON=1'b0;
    defparam data_index_i8_LC_15_19_6.SEQ_MODE=4'b1000;
    defparam data_index_i8_LC_15_19_6.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i8_LC_15_19_6 (
            .in0(N__44980),
            .in1(N__63743),
            .in2(N__57709),
            .in3(N__44971),
            .lcout(data_index_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61984),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_7_i15_4_lut_LC_15_19_7.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_7_i15_4_lut_LC_15_19_7.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_7_i15_4_lut_LC_15_19_7.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_358_Mux_7_i15_4_lut_LC_15_19_7 (
            .in0(N__63739),
            .in1(N__44925),
            .in2(N__57710),
            .in3(N__44916),
            .lcout(data_index_9_N_236_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i0_LC_15_20_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i0_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i0_LC_15_20_0 .LUT_INIT=16'b1100000001010101;
    LogicCell40 \SIG_DDS.dds_state_i0_LC_15_20_0  (
            .in0(N__50595),
            .in1(N__44812),
            .in2(N__44806),
            .in3(N__50330),
            .lcout(dds_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61996),
            .ce(N__47632),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_16_2_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_16_2_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_16_2_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_89_2_lut_LC_16_2_7  (
            .in0(_gnd_net_),
            .in1(N__50188),
            .in2(_gnd_net_),
            .in3(N__57119),
            .lcout(\comm_spi.imosi_N_841 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12616_12617_set_LC_16_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12616_12617_set_LC_16_3_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_rx_i0_12616_12617_set_LC_16_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_12616_12617_set_LC_16_3_0  (
            .in0(N__47958),
            .in1(N__44783),
            .in2(_gnd_net_),
            .in3(N__45460),
            .lcout(\comm_spi.n15344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53688),
            .ce(),
            .sr(N__47530));
    defparam \comm_spi.i12604_3_lut_LC_16_4_5 .C_ON=1'b0;
    defparam \comm_spi.i12604_3_lut_LC_16_4_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12604_3_lut_LC_16_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i12604_3_lut_LC_16_4_5  (
            .in0(N__47954),
            .in1(N__44784),
            .in2(_gnd_net_),
            .in3(N__45458),
            .lcout(\comm_spi.imosi ),
            .ltout(\comm_spi.imosi_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i20223_4_lut_3_lut_LC_16_4_6 .C_ON=1'b0;
    defparam \comm_spi.i20223_4_lut_3_lut_LC_16_4_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20223_4_lut_3_lut_LC_16_4_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \comm_spi.i20223_4_lut_3_lut_LC_16_4_6  (
            .in0(_gnd_net_),
            .in1(N__45244),
            .in2(N__45247),
            .in3(N__57070),
            .lcout(\comm_spi.n24019 ),
            .ltout(\comm_spi.n24019_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12618_3_lut_LC_16_4_7 .C_ON=1'b0;
    defparam \comm_spi.i12618_3_lut_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12618_3_lut_LC_16_4_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \comm_spi.i12618_3_lut_LC_16_4_7  (
            .in0(N__45238),
            .in1(N__45232),
            .in2(N__45226),
            .in3(_gnd_net_),
            .lcout(comm_rx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_112_LC_16_5_0.C_ON=1'b0;
    defparam i12_4_lut_adj_112_LC_16_5_0.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_112_LC_16_5_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_112_LC_16_5_0 (
            .in0(N__47919),
            .in1(N__48051),
            .in2(N__47833),
            .in3(N__48021),
            .lcout(n31_adj_1680),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_16_5_1.C_ON=1'b0;
    defparam i14_4_lut_LC_16_5_1.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_16_5_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_LC_16_5_1 (
            .in0(N__47937),
            .in1(N__47868),
            .in2(N__47890),
            .in3(N__48085),
            .lcout(n33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_adj_110_LC_16_5_2.C_ON=1'b0;
    defparam i13_4_lut_adj_110_LC_16_5_2.SEQ_MODE=4'b0000;
    defparam i13_4_lut_adj_110_LC_16_5_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_adj_110_LC_16_5_2 (
            .in0(N__47973),
            .in1(N__48235),
            .in2(N__48106),
            .in3(N__48202),
            .lcout(n32),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_202_LC_16_5_3.C_ON=1'b0;
    defparam i12_4_lut_adj_202_LC_16_5_3.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_202_LC_16_5_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_202_LC_16_5_3 (
            .in0(N__45222),
            .in1(N__45208),
            .in2(N__45190),
            .in3(N__45169),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_16_5_4.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_16_5_4.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_16_5_4.LUT_INIT=16'b1111111101110111;
    LogicCell40 i2_2_lut_3_lut_LC_16_5_4 (
            .in0(N__60063),
            .in1(N__60358),
            .in2(_gnd_net_),
            .in3(N__59185),
            .lcout(n11379),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_LC_16_6_0.C_ON=1'b0;
    defparam i11_4_lut_LC_16_6_0.SEQ_MODE=4'b0000;
    defparam i11_4_lut_LC_16_6_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_LC_16_6_0 (
            .in0(N__47904),
            .in1(N__48165),
            .in2(N__47854),
            .in3(N__48216),
            .lcout(n30_adj_1681),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_16_6_1.C_ON=1'b0;
    defparam i5_4_lut_LC_16_6_1.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_16_6_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i5_4_lut_LC_16_6_1 (
            .in0(N__48135),
            .in1(N__48120),
            .in2(N__48184),
            .in3(N__48150),
            .lcout(),
            .ltout(n12_adj_1760_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_16_6_2.C_ON=1'b0;
    defparam i6_4_lut_LC_16_6_2.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_16_6_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_LC_16_6_2 (
            .in0(N__48036),
            .in1(N__47991),
            .in2(N__45496),
            .in3(N__48436),
            .lcout(),
            .ltout(n20834_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_109_LC_16_6_3.C_ON=1'b0;
    defparam i15_4_lut_adj_109_LC_16_6_3.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_109_LC_16_6_3.LUT_INIT=16'b1111111111101111;
    LogicCell40 i15_4_lut_adj_109_LC_16_6_3 (
            .in0(N__48006),
            .in1(N__48066),
            .in2(N__45493),
            .in3(N__45490),
            .lcout(),
            .ltout(n34_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18_4_lut_LC_16_6_4.C_ON=1'b0;
    defparam i18_4_lut_LC_16_6_4.SEQ_MODE=4'b0000;
    defparam i18_4_lut_LC_16_6_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i18_4_lut_LC_16_6_4 (
            .in0(N__45484),
            .in1(N__45478),
            .in2(N__45472),
            .in3(N__45469),
            .lcout(n49),
            .ltout(n49_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam wdtick_flag_292_LC_16_6_5.C_ON=1'b0;
    defparam wdtick_flag_292_LC_16_6_5.SEQ_MODE=4'b1010;
    defparam wdtick_flag_292_LC_16_6_5.LUT_INIT=16'b1111111100001111;
    LogicCell40 wdtick_flag_292_LC_16_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45463),
            .in3(N__52659),
            .lcout(wdtick_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48405),
            .ce(),
            .sr(N__51225));
    defparam \comm_spi.i20208_4_lut_3_lut_LC_16_7_1 .C_ON=1'b0;
    defparam \comm_spi.i20208_4_lut_3_lut_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i20208_4_lut_3_lut_LC_16_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.i20208_4_lut_3_lut_LC_16_7_1  (
            .in0(N__45454),
            .in1(N__57049),
            .in2(_gnd_net_),
            .in3(N__50199),
            .lcout(\comm_spi.n24022 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_66_LC_16_7_6.C_ON=1'b0;
    defparam i1_2_lut_adj_66_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_66_LC_16_7_6.LUT_INIT=16'b0000000010101010;
    LogicCell40 i1_2_lut_adj_66_LC_16_7_6 (
            .in0(N__46199),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63073),
            .lcout(),
            .ltout(n8856_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_68_LC_16_7_7.C_ON=1'b0;
    defparam i1_4_lut_adj_68_LC_16_7_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_68_LC_16_7_7.LUT_INIT=16'b1100100010001000;
    LogicCell40 i1_4_lut_adj_68_LC_16_7_7 (
            .in0(N__57745),
            .in1(N__63601),
            .in2(N__45430),
            .in3(N__59190),
            .lcout(n13273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16182_3_lut_LC_16_8_0.C_ON=1'b0;
    defparam i16182_3_lut_LC_16_8_0.SEQ_MODE=4'b0000;
    defparam i16182_3_lut_LC_16_8_0.LUT_INIT=16'b1101100011011000;
    LogicCell40 i16182_3_lut_LC_16_8_0 (
            .in0(N__54527),
            .in1(N__55093),
            .in2(N__45328),
            .in3(_gnd_net_),
            .lcout(n18882),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19916_2_lut_LC_16_8_1.C_ON=1'b0;
    defparam i19916_2_lut_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam i19916_2_lut_LC_16_8_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19916_2_lut_LC_16_8_1 (
            .in0(_gnd_net_),
            .in1(N__45727),
            .in2(_gnd_net_),
            .in3(N__54525),
            .lcout(n22371),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16183_3_lut_LC_16_8_2.C_ON=1'b0;
    defparam i16183_3_lut_LC_16_8_2.SEQ_MODE=4'b0000;
    defparam i16183_3_lut_LC_16_8_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 i16183_3_lut_LC_16_8_2 (
            .in0(N__54528),
            .in1(_gnd_net_),
            .in2(N__45715),
            .in3(N__45700),
            .lcout(),
            .ltout(n18883_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i5_LC_16_8_3.C_ON=1'b0;
    defparam comm_tx_buf_i5_LC_16_8_3.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i5_LC_16_8_3.LUT_INIT=16'b1100110011100010;
    LogicCell40 comm_tx_buf_i5_LC_16_8_3 (
            .in0(N__45667),
            .in1(N__45607),
            .in2(N__45661),
            .in3(N__54307),
            .lcout(comm_tx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61850),
            .ce(N__46419),
            .sr(N__46341));
    defparam i16185_3_lut_LC_16_8_4.C_ON=1'b0;
    defparam i16185_3_lut_LC_16_8_4.SEQ_MODE=4'b0000;
    defparam i16185_3_lut_LC_16_8_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 i16185_3_lut_LC_16_8_4 (
            .in0(N__54526),
            .in1(N__45625),
            .in2(_gnd_net_),
            .in3(N__56578),
            .lcout(),
            .ltout(n18885_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_LC_16_8_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_LC_16_8_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_LC_16_8_5.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_index_1__bdd_4_lut_LC_16_8_5 (
            .in0(N__45616),
            .in1(N__54306),
            .in2(N__45610),
            .in3(N__51800),
            .lcout(n23414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20060_2_lut_LC_16_9_0.C_ON=1'b0;
    defparam i20060_2_lut_LC_16_9_0.SEQ_MODE=4'b0000;
    defparam i20060_2_lut_LC_16_9_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 i20060_2_lut_LC_16_9_0 (
            .in0(N__58949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51730),
            .lcout(n22618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i3_LC_16_9_1.C_ON=1'b0;
    defparam comm_buf_6__i3_LC_16_9_1.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i3_LC_16_9_1.LUT_INIT=16'b0000101011001010;
    LogicCell40 comm_buf_6__i3_LC_16_9_1 (
            .in0(N__46257),
            .in1(N__62784),
            .in2(N__45571),
            .in3(N__63595),
            .lcout(comm_buf_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61857),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_211_LC_16_9_2.C_ON=1'b0;
    defparam i1_4_lut_adj_211_LC_16_9_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_211_LC_16_9_2.LUT_INIT=16'b1110000010100000;
    LogicCell40 i1_4_lut_adj_211_LC_16_9_2 (
            .in0(N__63594),
            .in1(N__45586),
            .in2(N__63200),
            .in3(N__48301),
            .lcout(n12976),
            .ltout(n12976_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i2_LC_16_9_3.C_ON=1'b0;
    defparam comm_buf_6__i2_LC_16_9_3.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i2_LC_16_9_3.LUT_INIT=16'b0000110010101100;
    LogicCell40 comm_buf_6__i2_LC_16_9_3 (
            .in0(N__54925),
            .in1(N__45510),
            .in2(N__45520),
            .in3(N__63596),
            .lcout(comm_buf_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61857),
            .ce(),
            .sr(_gnd_net_));
    defparam i19807_4_lut_LC_16_9_4.C_ON=1'b0;
    defparam i19807_4_lut_LC_16_9_4.SEQ_MODE=4'b0000;
    defparam i19807_4_lut_LC_16_9_4.LUT_INIT=16'b0100000000000000;
    LogicCell40 i19807_4_lut_LC_16_9_4 (
            .in0(N__58950),
            .in1(N__60952),
            .in2(N__48271),
            .in3(N__60396),
            .lcout(),
            .ltout(n22375_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i2_LC_16_9_5.C_ON=1'b0;
    defparam comm_length_i2_LC_16_9_5.SEQ_MODE=4'b1000;
    defparam comm_length_i2_LC_16_9_5.LUT_INIT=16'b1111011110000000;
    LogicCell40 comm_length_i2_LC_16_9_5 (
            .in0(N__51514),
            .in1(N__63188),
            .in2(N__45847),
            .in3(N__48642),
            .lcout(comm_length_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61857),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_346_Mux_2_i4_3_lut_LC_16_9_6.C_ON=1'b0;
    defparam comm_state_3__I_0_346_Mux_2_i4_3_lut_LC_16_9_6.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_346_Mux_2_i4_3_lut_LC_16_9_6.LUT_INIT=16'b0011001110101010;
    LogicCell40 comm_state_3__I_0_346_Mux_2_i4_3_lut_LC_16_9_6 (
            .in0(N__45856),
            .in1(N__58210),
            .in2(_gnd_net_),
            .in3(N__62936),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20075_2_lut_LC_16_9_7.C_ON=1'b0;
    defparam i20075_2_lut_LC_16_9_7.SEQ_MODE=4'b0000;
    defparam i20075_2_lut_LC_16_9_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i20075_2_lut_LC_16_9_7 (
            .in0(_gnd_net_),
            .in1(N__45844),
            .in2(_gnd_net_),
            .in3(N__58948),
            .lcout(n22297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.bit_cnt_3787__i3_LC_16_10_0 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3787__i3_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3787__i3_LC_16_10_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \comm_spi.bit_cnt_3787__i3_LC_16_10_0  (
            .in0(N__51424),
            .in1(N__53771),
            .in2(N__51451),
            .in3(N__51472),
            .lcout(\comm_spi.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3787__i3C_net ),
            .ce(),
            .sr(N__57122));
    defparam \comm_spi.bit_cnt_3787__i2_LC_16_10_1 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3787__i2_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3787__i2_LC_16_10_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \comm_spi.bit_cnt_3787__i2_LC_16_10_1  (
            .in0(N__51471),
            .in1(N__51446),
            .in2(_gnd_net_),
            .in3(N__51423),
            .lcout(\comm_spi.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3787__i3C_net ),
            .ce(),
            .sr(N__57122));
    defparam \comm_spi.bit_cnt_3787__i1_LC_16_10_2 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3787__i1_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3787__i1_LC_16_10_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \comm_spi.bit_cnt_3787__i1_LC_16_10_2  (
            .in0(N__51445),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51470),
            .lcout(\comm_spi.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3787__i3C_net ),
            .ce(),
            .sr(N__57122));
    defparam \comm_spi.bit_cnt_3787__i0_LC_16_10_3 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3787__i0_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3787__i0_LC_16_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \comm_spi.bit_cnt_3787__i0_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51444),
            .lcout(\comm_spi.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3787__i3C_net ),
            .ce(),
            .sr(N__57122));
    defparam i12699_2_lut_LC_16_10_6.C_ON=1'b0;
    defparam i12699_2_lut_LC_16_10_6.SEQ_MODE=4'b0000;
    defparam i12699_2_lut_LC_16_10_6.LUT_INIT=16'b0011001100000000;
    LogicCell40 i12699_2_lut_LC_16_10_6 (
            .in0(_gnd_net_),
            .in1(N__45817),
            .in2(_gnd_net_),
            .in3(N__50020),
            .lcout(n15431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12794_2_lut_LC_16_10_7.C_ON=1'b0;
    defparam i12794_2_lut_LC_16_10_7.SEQ_MODE=4'b0000;
    defparam i12794_2_lut_LC_16_10_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12794_2_lut_LC_16_10_7 (
            .in0(_gnd_net_),
            .in1(N__63597),
            .in2(_gnd_net_),
            .in3(N__45885),
            .lcout(n15517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_226_LC_16_11_0.C_ON=1'b0;
    defparam i1_2_lut_adj_226_LC_16_11_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_226_LC_16_11_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_226_LC_16_11_0 (
            .in0(_gnd_net_),
            .in1(N__46474),
            .in2(_gnd_net_),
            .in3(N__46520),
            .lcout(n21966),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i1_LC_16_11_1.C_ON=1'b0;
    defparam comm_cmd_i1_LC_16_11_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i1_LC_16_11_1.LUT_INIT=16'b1011100000110000;
    LogicCell40 comm_cmd_i1_LC_16_11_1 (
            .in0(N__54792),
            .in1(N__46007),
            .in2(N__60357),
            .in3(N__45949),
            .lcout(comm_cmd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61877),
            .ce(),
            .sr(_gnd_net_));
    defparam i16279_2_lut_LC_16_11_2.C_ON=1'b0;
    defparam i16279_2_lut_LC_16_11_2.SEQ_MODE=4'b0000;
    defparam i16279_2_lut_LC_16_11_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i16279_2_lut_LC_16_11_2 (
            .in0(_gnd_net_),
            .in1(N__60233),
            .in2(_gnd_net_),
            .in3(N__58840),
            .lcout(n18955),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_332_LC_16_11_3.C_ON=1'b0;
    defparam i1_3_lut_adj_332_LC_16_11_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_332_LC_16_11_3.LUT_INIT=16'b1100110010001000;
    LogicCell40 i1_3_lut_adj_332_LC_16_11_3 (
            .in0(N__54171),
            .in1(N__54068),
            .in2(_gnd_net_),
            .in3(N__49348),
            .lcout(n12958),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i58_4_lut_LC_16_11_4.C_ON=1'b0;
    defparam i58_4_lut_LC_16_11_4.SEQ_MODE=4'b0000;
    defparam i58_4_lut_LC_16_11_4.LUT_INIT=16'b0100111001000100;
    LogicCell40 i58_4_lut_LC_16_11_4 (
            .in0(N__62530),
            .in1(N__45874),
            .in2(N__54418),
            .in3(N__48901),
            .lcout(n29_adj_1688),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_79_LC_16_11_5.C_ON=1'b0;
    defparam i1_2_lut_adj_79_LC_16_11_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_79_LC_16_11_5.LUT_INIT=16'b1111111101010101;
    LogicCell40 i1_2_lut_adj_79_LC_16_11_5 (
            .in0(N__58610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50858),
            .lcout(),
            .ltout(n11402_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_133_Mux_2_i127_4_lut_LC_16_11_6.C_ON=1'b0;
    defparam mux_133_Mux_2_i127_4_lut_LC_16_11_6.SEQ_MODE=4'b0000;
    defparam mux_133_Mux_2_i127_4_lut_LC_16_11_6.LUT_INIT=16'b0000101011001100;
    LogicCell40 mux_133_Mux_2_i127_4_lut_LC_16_11_6 (
            .in0(N__55598),
            .in1(N__58403),
            .in2(N__45859),
            .in3(N__61380),
            .lcout(comm_state_3_N_500_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19773_2_lut_4_lut_LC_16_11_7.C_ON=1'b0;
    defparam i19773_2_lut_4_lut_LC_16_11_7.SEQ_MODE=4'b0000;
    defparam i19773_2_lut_4_lut_LC_16_11_7.LUT_INIT=16'b0101000001000000;
    LogicCell40 i19773_2_lut_4_lut_LC_16_11_7 (
            .in0(N__60902),
            .in1(N__58841),
            .in2(N__58521),
            .in3(N__60247),
            .lcout(n22351),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16149_3_lut_LC_16_12_0.C_ON=1'b0;
    defparam i16149_3_lut_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam i16149_3_lut_LC_16_12_0.LUT_INIT=16'b1111101001010000;
    LogicCell40 i16149_3_lut_LC_16_12_0 (
            .in0(N__54542),
            .in1(_gnd_net_),
            .in2(N__62092),
            .in3(N__54949),
            .lcout(),
            .ltout(n18850_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i3_LC_16_12_1.C_ON=1'b0;
    defparam comm_tx_buf_i3_LC_16_12_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i3_LC_16_12_1.LUT_INIT=16'b1010101011011000;
    LogicCell40 comm_tx_buf_i3_LC_16_12_1 (
            .in0(N__46210),
            .in1(N__46237),
            .in2(N__46435),
            .in3(N__54331),
            .lcout(comm_tx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61889),
            .ce(N__46432),
            .sr(N__46353));
    defparam i19787_2_lut_LC_16_12_2.C_ON=1'b0;
    defparam i19787_2_lut_LC_16_12_2.SEQ_MODE=4'b0000;
    defparam i19787_2_lut_LC_16_12_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 i19787_2_lut_LC_16_12_2 (
            .in0(N__54539),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46276),
            .lcout(n22346),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16150_3_lut_LC_16_12_3.C_ON=1'b0;
    defparam i16150_3_lut_LC_16_12_3.SEQ_MODE=4'b0000;
    defparam i16150_3_lut_LC_16_12_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i16150_3_lut_LC_16_12_3 (
            .in0(N__46258),
            .in1(N__46109),
            .in2(_gnd_net_),
            .in3(N__54541),
            .lcout(n18851),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16152_3_lut_LC_16_12_4.C_ON=1'b0;
    defparam i16152_3_lut_LC_16_12_4.SEQ_MODE=4'b0000;
    defparam i16152_3_lut_LC_16_12_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 i16152_3_lut_LC_16_12_4 (
            .in0(N__54540),
            .in1(_gnd_net_),
            .in2(N__49292),
            .in3(N__46228),
            .lcout(),
            .ltout(n18853_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_20444_LC_16_12_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_20444_LC_16_12_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_20444_LC_16_12_5.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_index_1__bdd_4_lut_20444_LC_16_12_5 (
            .in0(N__46219),
            .in1(N__54330),
            .in2(N__46213),
            .in3(N__51829),
            .lcout(n23378),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16157_3_lut_LC_16_12_6.C_ON=1'b0;
    defparam i16157_3_lut_LC_16_12_6.SEQ_MODE=4'b0000;
    defparam i16157_3_lut_LC_16_12_6.LUT_INIT=16'b1110001011100010;
    LogicCell40 i16157_3_lut_LC_16_12_6 (
            .in0(N__62079),
            .in1(N__46200),
            .in2(N__46116),
            .in3(_gnd_net_),
            .lcout(n18858),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_16_12_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_16_12_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_104_2_lut_LC_16_12_7  (
            .in0(N__46058),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57129),
            .lcout(\comm_spi.data_tx_7__N_874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i7_LC_16_13_0.C_ON=1'b0;
    defparam buf_control_i7_LC_16_13_0.SEQ_MODE=4'b1000;
    defparam buf_control_i7_LC_16_13_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 buf_control_i7_LC_16_13_0 (
            .in0(N__46045),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buf_control_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61905),
            .ce(N__46687),
            .sr(N__51646));
    defparam i1_2_lut_adj_227_LC_16_13_1.C_ON=1'b0;
    defparam i1_2_lut_adj_227_LC_16_13_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_227_LC_16_13_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_adj_227_LC_16_13_1 (
            .in0(N__63050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64033),
            .lcout(),
            .ltout(n12021_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_291_LC_16_13_2.C_ON=1'b0;
    defparam i1_4_lut_adj_291_LC_16_13_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_291_LC_16_13_2.LUT_INIT=16'b1010101000001000;
    LogicCell40 i1_4_lut_adj_291_LC_16_13_2 (
            .in0(N__63196),
            .in1(N__62675),
            .in2(N__46690),
            .in3(N__63718),
            .lcout(n12614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i44_3_lut_LC_16_13_3.C_ON=1'b0;
    defparam i44_3_lut_LC_16_13_3.SEQ_MODE=4'b0000;
    defparam i44_3_lut_LC_16_13_3.LUT_INIT=16'b0110011000100010;
    LogicCell40 i44_3_lut_LC_16_13_3 (
            .in0(N__63049),
            .in1(N__64031),
            .in2(_gnd_net_),
            .in3(N__54198),
            .lcout(),
            .ltout(n25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_290_LC_16_13_4.C_ON=1'b0;
    defparam i1_4_lut_adj_290_LC_16_13_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_290_LC_16_13_4.LUT_INIT=16'b1010101000100000;
    LogicCell40 i1_4_lut_adj_290_LC_16_13_4 (
            .in0(N__63195),
            .in1(N__62673),
            .in2(N__46681),
            .in3(N__63717),
            .lcout(n12548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6984_2_lut_LC_16_13_6.C_ON=1'b0;
    defparam i6984_2_lut_LC_16_13_6.SEQ_MODE=4'b0000;
    defparam i6984_2_lut_LC_16_13_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 i6984_2_lut_LC_16_13_6 (
            .in0(N__62564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63048),
            .lcout(n9714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16459_2_lut_3_lut_LC_16_13_7.C_ON=1'b0;
    defparam i16459_2_lut_3_lut_LC_16_13_7.SEQ_MODE=4'b0000;
    defparam i16459_2_lut_3_lut_LC_16_13_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16459_2_lut_3_lut_LC_16_13_7 (
            .in0(N__62674),
            .in1(N__46642),
            .in2(_gnd_net_),
            .in3(N__64032),
            .lcout(n14_adj_1607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_306_LC_16_14_0.C_ON=1'b0;
    defparam i1_4_lut_adj_306_LC_16_14_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_306_LC_16_14_0.LUT_INIT=16'b1010101100000000;
    LogicCell40 i1_4_lut_adj_306_LC_16_14_0 (
            .in0(N__57712),
            .in1(N__46530),
            .in2(N__46504),
            .in3(N__63650),
            .lcout(n13129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19133_2_lut_LC_16_14_1.C_ON=1'b0;
    defparam i19133_2_lut_LC_16_14_1.SEQ_MODE=4'b0000;
    defparam i19133_2_lut_LC_16_14_1.LUT_INIT=16'b1100110011111111;
    LogicCell40 i19133_2_lut_LC_16_14_1 (
            .in0(_gnd_net_),
            .in1(N__46482),
            .in2(_gnd_net_),
            .in3(N__58624),
            .lcout(n22059),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_3_i26_3_lut_LC_16_14_2.C_ON=1'b0;
    defparam mux_126_Mux_3_i26_3_lut_LC_16_14_2.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_3_i26_3_lut_LC_16_14_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_126_Mux_3_i26_3_lut_LC_16_14_2 (
            .in0(N__59226),
            .in1(_gnd_net_),
            .in2(N__47137),
            .in3(N__49811),
            .lcout(n26_adj_1740),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_0_i26_3_lut_LC_16_14_3.C_ON=1'b0;
    defparam mux_126_Mux_0_i26_3_lut_LC_16_14_3.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_0_i26_3_lut_LC_16_14_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_126_Mux_0_i26_3_lut_LC_16_14_3 (
            .in0(N__47203),
            .in1(N__59225),
            .in2(_gnd_net_),
            .in3(N__49388),
            .lcout(),
            .ltout(n26_adj_1580_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20582_LC_16_14_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20582_LC_16_14_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20582_LC_16_14_4.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20582_LC_16_14_4 (
            .in0(N__58666),
            .in1(N__59974),
            .in2(N__47041),
            .in3(N__60395),
            .lcout(),
            .ltout(n23552_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23552_bdd_4_lut_LC_16_14_5.C_ON=1'b0;
    defparam n23552_bdd_4_lut_LC_16_14_5.SEQ_MODE=4'b0000;
    defparam n23552_bdd_4_lut_LC_16_14_5.LUT_INIT=16'b1111010010100100;
    LogicCell40 n23552_bdd_4_lut_LC_16_14_5 (
            .in0(N__59975),
            .in1(N__47038),
            .in2(N__47017),
            .in3(N__47009),
            .lcout(n23555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i4_LC_16_14_6.C_ON=1'b0;
    defparam req_data_cnt_i4_LC_16_14_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i4_LC_16_14_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i4_LC_16_14_6 (
            .in0(N__56022),
            .in1(N__51324),
            .in2(_gnd_net_),
            .in3(N__52481),
            .lcout(req_data_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61919),
            .ce(),
            .sr(_gnd_net_));
    defparam n23300_bdd_4_lut_LC_16_15_0.C_ON=1'b0;
    defparam n23300_bdd_4_lut_LC_16_15_0.SEQ_MODE=4'b0000;
    defparam n23300_bdd_4_lut_LC_16_15_0.LUT_INIT=16'b1100110011100010;
    LogicCell40 n23300_bdd_4_lut_LC_16_15_0 (
            .in0(N__46990),
            .in1(N__46975),
            .in2(N__46960),
            .in3(N__59976),
            .lcout(n23303),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19344_3_lut_LC_16_15_1.C_ON=1'b0;
    defparam i19344_3_lut_LC_16_15_1.SEQ_MODE=4'b0000;
    defparam i19344_3_lut_LC_16_15_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 i19344_3_lut_LC_16_15_1 (
            .in0(N__46920),
            .in1(N__46879),
            .in2(_gnd_net_),
            .in3(N__60497),
            .lcout(n22271),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19341_3_lut_LC_16_15_2.C_ON=1'b0;
    defparam i19341_3_lut_LC_16_15_2.SEQ_MODE=4'b0000;
    defparam i19341_3_lut_LC_16_15_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 i19341_3_lut_LC_16_15_2 (
            .in0(N__59209),
            .in1(N__47476),
            .in2(_gnd_net_),
            .in3(N__49742),
            .lcout(n22268),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i4_LC_16_15_4.C_ON=1'b0;
    defparam acadc_skipCount_i4_LC_16_15_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i4_LC_16_15_4.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i4_LC_16_15_4 (
            .in0(N__57853),
            .in1(N__46851),
            .in2(N__52513),
            .in3(N__56069),
            .lcout(acadc_skipCount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61939),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i0_LC_16_15_5.C_ON=1'b0;
    defparam buf_control_i0_LC_16_15_5.SEQ_MODE=4'b1000;
    defparam buf_control_i0_LC_16_15_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_control_i0_LC_16_15_5 (
            .in0(N__48879),
            .in1(N__46748),
            .in2(_gnd_net_),
            .in3(N__52625),
            .lcout(buf_control_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61939),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i4_LC_16_15_6.C_ON=1'b0;
    defparam buf_dds0_i4_LC_16_15_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i4_LC_16_15_6.LUT_INIT=16'b0111001001010000;
    LogicCell40 buf_dds0_i4_LC_16_15_6 (
            .in0(N__50769),
            .in1(N__57852),
            .in2(N__47267),
            .in3(N__56070),
            .lcout(buf_dds0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61939),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i0_LC_16_15_7.C_ON=1'b0;
    defparam buf_dds0_i0_LC_16_15_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i0_LC_16_15_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_dds0_i0_LC_16_15_7 (
            .in0(N__57851),
            .in1(N__50768),
            .in2(N__49140),
            .in3(N__47219),
            .lcout(buf_dds0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61939),
            .ce(),
            .sr(_gnd_net_));
    defparam data_idxvec_i0_LC_16_16_0.C_ON=1'b1;
    defparam data_idxvec_i0_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i0_LC_16_16_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i0_LC_16_16_0 (
            .in0(N__48250),
            .in1(N__47202),
            .in2(N__63763),
            .in3(N__47188),
            .lcout(data_idxvec_0),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(n20661),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i1_LC_16_16_1.C_ON=1'b1;
    defparam data_idxvec_i1_LC_16_16_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i1_LC_16_16_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i1_LC_16_16_1 (
            .in0(N__47175),
            .in1(N__52272),
            .in2(N__63767),
            .in3(N__47161),
            .lcout(data_idxvec_1),
            .ltout(),
            .carryin(n20661),
            .carryout(n20662),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i2_LC_16_16_2.C_ON=1'b1;
    defparam data_idxvec_i2_LC_16_16_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i2_LC_16_16_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i2_LC_16_16_2 (
            .in0(N__47158),
            .in1(N__52420),
            .in2(N__63764),
            .in3(N__47140),
            .lcout(data_idxvec_2),
            .ltout(),
            .carryin(n20662),
            .carryout(n20663),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i3_LC_16_16_3.C_ON=1'b1;
    defparam data_idxvec_i3_LC_16_16_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i3_LC_16_16_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i3_LC_16_16_3 (
            .in0(N__48942),
            .in1(N__47133),
            .in2(N__63768),
            .in3(N__47119),
            .lcout(data_idxvec_3),
            .ltout(),
            .carryin(n20663),
            .carryout(n20664),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i4_LC_16_16_4.C_ON=1'b1;
    defparam data_idxvec_i4_LC_16_16_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i4_LC_16_16_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i4_LC_16_16_4 (
            .in0(N__56023),
            .in1(N__52563),
            .in2(N__63765),
            .in3(N__47116),
            .lcout(data_idxvec_4),
            .ltout(),
            .carryin(n20664),
            .carryout(n20665),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i5_LC_16_16_5.C_ON=1'b1;
    defparam data_idxvec_i5_LC_16_16_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i5_LC_16_16_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i5_LC_16_16_5 (
            .in0(N__47099),
            .in1(N__51999),
            .in2(N__63769),
            .in3(N__47080),
            .lcout(data_idxvec_5),
            .ltout(),
            .carryin(n20665),
            .carryout(n20666),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i6_LC_16_16_6.C_ON=1'b1;
    defparam data_idxvec_i6_LC_16_16_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i6_LC_16_16_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i6_LC_16_16_6 (
            .in0(N__47069),
            .in1(N__49605),
            .in2(N__63766),
            .in3(N__47044),
            .lcout(data_idxvec_6),
            .ltout(),
            .carryin(n20666),
            .carryout(n20667),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i7_LC_16_16_7.C_ON=1'b1;
    defparam data_idxvec_i7_LC_16_16_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i7_LC_16_16_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i7_LC_16_16_7 (
            .in0(N__47516),
            .in1(N__54672),
            .in2(N__63770),
            .in3(N__47479),
            .lcout(data_idxvec_7),
            .ltout(),
            .carryin(n20667),
            .carryout(n20668),
            .clk(N__61955),
            .ce(N__47692),
            .sr(_gnd_net_));
    defparam data_idxvec_i8_LC_16_17_0.C_ON=1'b1;
    defparam data_idxvec_i8_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i8_LC_16_17_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i8_LC_16_17_0 (
            .in0(N__48871),
            .in1(N__47475),
            .in2(N__63779),
            .in3(N__47461),
            .lcout(data_idxvec_8),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(n20669),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_idxvec_i9_LC_16_17_1.C_ON=1'b1;
    defparam data_idxvec_i9_LC_16_17_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i9_LC_16_17_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i9_LC_16_17_1 (
            .in0(N__50797),
            .in1(N__63748),
            .in2(N__50953),
            .in3(N__47458),
            .lcout(data_idxvec_9),
            .ltout(),
            .carryin(n20669),
            .carryout(n20670),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_idxvec_i10_LC_16_17_2.C_ON=1'b1;
    defparam data_idxvec_i10_LC_16_17_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i10_LC_16_17_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i10_LC_16_17_2 (
            .in0(N__47451),
            .in1(N__47392),
            .in2(N__63780),
            .in3(N__47380),
            .lcout(data_idxvec_10),
            .ltout(),
            .carryin(n20670),
            .carryout(n20671),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_idxvec_i11_LC_16_17_3.C_ON=1'b1;
    defparam data_idxvec_i11_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i11_LC_16_17_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i11_LC_16_17_3 (
            .in0(N__56834),
            .in1(N__63752),
            .in2(N__56157),
            .in3(N__47377),
            .lcout(data_idxvec_11),
            .ltout(),
            .carryin(n20671),
            .carryout(n20672),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_idxvec_i12_LC_16_17_4.C_ON=1'b1;
    defparam data_idxvec_i12_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i12_LC_16_17_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i12_LC_16_17_4 (
            .in0(N__47352),
            .in1(N__49719),
            .in2(N__63781),
            .in3(N__47317),
            .lcout(data_idxvec_12),
            .ltout(),
            .carryin(n20672),
            .carryout(n20673),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_idxvec_i13_LC_16_17_5.C_ON=1'b1;
    defparam data_idxvec_i13_LC_16_17_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i13_LC_16_17_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i13_LC_16_17_5 (
            .in0(N__55287),
            .in1(N__63756),
            .in2(N__61095),
            .in3(N__47314),
            .lcout(data_idxvec_13),
            .ltout(),
            .carryin(n20673),
            .carryout(n20674),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_idxvec_i14_LC_16_17_6.C_ON=1'b1;
    defparam data_idxvec_i14_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i14_LC_16_17_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i14_LC_16_17_6 (
            .in0(N__51501),
            .in1(N__49026),
            .in2(N__63782),
            .in3(N__47311),
            .lcout(data_idxvec_14),
            .ltout(),
            .carryin(n20674),
            .carryout(n20675),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_idxvec_i15_LC_16_17_7.C_ON=1'b0;
    defparam data_idxvec_i15_LC_16_17_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i15_LC_16_17_7.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i15_LC_16_17_7 (
            .in0(N__47308),
            .in1(N__63760),
            .in2(N__47289),
            .in3(N__47296),
            .lcout(data_idxvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61972),
            .ce(N__47691),
            .sr(_gnd_net_));
    defparam data_index_i0_LC_16_18_1.C_ON=1'b0;
    defparam data_index_i0_LC_16_18_1.SEQ_MODE=4'b1000;
    defparam data_index_i0_LC_16_18_1.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i0_LC_16_18_1 (
            .in0(N__52587),
            .in1(N__63761),
            .in2(N__57855),
            .in3(N__53152),
            .lcout(data_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61985),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i20157_4_lut_LC_16_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.i20157_4_lut_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i20157_4_lut_LC_16_18_2 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \SIG_DDS.i20157_4_lut_LC_16_18_2  (
            .in0(N__50610),
            .in1(N__50536),
            .in2(N__47582),
            .in3(N__50314),
            .lcout(\SIG_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_LC_16_18_3.C_ON=1'b0;
    defparam i15_4_lut_LC_16_18_3.SEQ_MODE=4'b0000;
    defparam i15_4_lut_LC_16_18_3.LUT_INIT=16'b1010001011110111;
    LogicCell40 i15_4_lut_LC_16_18_3 (
            .in0(N__63744),
            .in1(N__56479),
            .in2(N__57854),
            .in3(N__47788),
            .lcout(n13052),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i12835_3_lut_LC_16_18_6 .C_ON=1'b0;
    defparam \SIG_DDS.i12835_3_lut_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i12835_3_lut_LC_16_18_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \SIG_DDS.i12835_3_lut_LC_16_18_6  (
            .in0(N__50609),
            .in1(N__50535),
            .in2(_gnd_net_),
            .in3(N__50315),
            .lcout(n15562),
            .ltout(n15562_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i0_LC_16_18_7 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i0_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i0_LC_16_18_7 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \SIG_DDS.bit_cnt_i0_LC_16_18_7  (
            .in0(N__50316),
            .in1(_gnd_net_),
            .in2(N__47665),
            .in3(N__47655),
            .lcout(bit_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61985),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i1_LC_16_19_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i1_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i1_LC_16_19_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \SIG_DDS.dds_state_i1_LC_16_19_0  (
            .in0(N__50599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50537),
            .lcout(dds_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61997),
            .ce(N__47625),
            .sr(N__50405));
    defparam \SIG_DDS.SCLK_27_LC_16_20_2 .C_ON=1'b0;
    defparam \SIG_DDS.SCLK_27_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.SCLK_27_LC_16_20_2 .LUT_INIT=16'b0011001010110001;
    LogicCell40 \SIG_DDS.SCLK_27_LC_16_20_2  (
            .in0(N__50594),
            .in1(N__50491),
            .in2(N__47601),
            .in3(N__50318),
            .lcout(DDS_SCK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62002),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i23_4_lut_LC_16_20_6 .C_ON=1'b0;
    defparam \SIG_DDS.i23_4_lut_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i23_4_lut_LC_16_20_6 .LUT_INIT=16'b1100110010011011;
    LogicCell40 \SIG_DDS.i23_4_lut_LC_16_20_6  (
            .in0(N__50593),
            .in1(N__50490),
            .in2(N__47583),
            .in3(N__50317),
            .lcout(\SIG_DDS.n9_adj_1490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_17_3_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_17_3_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_17_3_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_86_2_lut_LC_17_3_6  (
            .in0(N__47541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57096),
            .lcout(\comm_spi.DOUT_7__N_834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_12602_12603_set_LC_17_4_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12602_12603_set_LC_17_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imosi_44_12602_12603_set_LC_17_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_12602_12603_set_LC_17_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50198),
            .lcout(\comm_spi.n15330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61832),
            .ce(),
            .sr(N__50140));
    defparam wdtick_cnt_3783_3784__i1_LC_17_5_0.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i1_LC_17_5_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i1_LC_17_5_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i1_LC_17_5_0 (
            .in0(N__48541),
            .in1(N__47938),
            .in2(_gnd_net_),
            .in3(N__47923),
            .lcout(wdtick_cnt_0),
            .ltout(),
            .carryin(bfn_17_5_0_),
            .carryout(n20766),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i2_LC_17_5_1.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i2_LC_17_5_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i2_LC_17_5_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i2_LC_17_5_1 (
            .in0(N__48510),
            .in1(N__47920),
            .in2(_gnd_net_),
            .in3(N__47908),
            .lcout(wdtick_cnt_1),
            .ltout(),
            .carryin(n20766),
            .carryout(n20767),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i3_LC_17_5_2.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i3_LC_17_5_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i3_LC_17_5_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i3_LC_17_5_2 (
            .in0(N__48542),
            .in1(N__47905),
            .in2(_gnd_net_),
            .in3(N__47893),
            .lcout(wdtick_cnt_2),
            .ltout(),
            .carryin(n20767),
            .carryout(n20768),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i4_LC_17_5_3.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i4_LC_17_5_3.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i4_LC_17_5_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i4_LC_17_5_3 (
            .in0(N__48511),
            .in1(N__47883),
            .in2(_gnd_net_),
            .in3(N__47872),
            .lcout(wdtick_cnt_3),
            .ltout(),
            .carryin(n20768),
            .carryout(n20769),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i5_LC_17_5_4.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i5_LC_17_5_4.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i5_LC_17_5_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i5_LC_17_5_4 (
            .in0(N__48543),
            .in1(N__47869),
            .in2(_gnd_net_),
            .in3(N__47857),
            .lcout(wdtick_cnt_4),
            .ltout(),
            .carryin(n20769),
            .carryout(n20770),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i6_LC_17_5_5.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i6_LC_17_5_5.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i6_LC_17_5_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i6_LC_17_5_5 (
            .in0(N__48512),
            .in1(N__47847),
            .in2(_gnd_net_),
            .in3(N__47836),
            .lcout(wdtick_cnt_5),
            .ltout(),
            .carryin(n20770),
            .carryout(n20771),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i7_LC_17_5_6.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i7_LC_17_5_6.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i7_LC_17_5_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i7_LC_17_5_6 (
            .in0(N__48544),
            .in1(N__47832),
            .in2(_gnd_net_),
            .in3(N__47818),
            .lcout(wdtick_cnt_6),
            .ltout(),
            .carryin(n20771),
            .carryout(n20772),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i8_LC_17_5_7.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i8_LC_17_5_7.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i8_LC_17_5_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i8_LC_17_5_7 (
            .in0(N__48513),
            .in1(N__48099),
            .in2(_gnd_net_),
            .in3(N__48088),
            .lcout(wdtick_cnt_7),
            .ltout(),
            .carryin(n20772),
            .carryout(n20773),
            .clk(N__48406),
            .ce(N__48349),
            .sr(N__51226));
    defparam wdtick_cnt_3783_3784__i9_LC_17_6_0.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i9_LC_17_6_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i9_LC_17_6_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i9_LC_17_6_0 (
            .in0(N__48505),
            .in1(N__48084),
            .in2(_gnd_net_),
            .in3(N__48070),
            .lcout(wdtick_cnt_8),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(n20774),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i10_LC_17_6_1.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i10_LC_17_6_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i10_LC_17_6_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i10_LC_17_6_1 (
            .in0(N__48533),
            .in1(N__48067),
            .in2(_gnd_net_),
            .in3(N__48055),
            .lcout(wdtick_cnt_9),
            .ltout(),
            .carryin(n20774),
            .carryout(n20775),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i11_LC_17_6_2.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i11_LC_17_6_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i11_LC_17_6_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i11_LC_17_6_2 (
            .in0(N__48502),
            .in1(N__48052),
            .in2(_gnd_net_),
            .in3(N__48040),
            .lcout(wdtick_cnt_10),
            .ltout(),
            .carryin(n20775),
            .carryout(n20776),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i12_LC_17_6_3.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i12_LC_17_6_3.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i12_LC_17_6_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i12_LC_17_6_3 (
            .in0(N__48534),
            .in1(N__48037),
            .in2(_gnd_net_),
            .in3(N__48025),
            .lcout(wdtick_cnt_11),
            .ltout(),
            .carryin(n20776),
            .carryout(n20777),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i13_LC_17_6_4.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i13_LC_17_6_4.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i13_LC_17_6_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i13_LC_17_6_4 (
            .in0(N__48503),
            .in1(N__48022),
            .in2(_gnd_net_),
            .in3(N__48010),
            .lcout(wdtick_cnt_12),
            .ltout(),
            .carryin(n20777),
            .carryout(n20778),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i14_LC_17_6_5.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i14_LC_17_6_5.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i14_LC_17_6_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i14_LC_17_6_5 (
            .in0(N__48535),
            .in1(N__48007),
            .in2(_gnd_net_),
            .in3(N__47995),
            .lcout(wdtick_cnt_13),
            .ltout(),
            .carryin(n20778),
            .carryout(n20779),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i15_LC_17_6_6.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i15_LC_17_6_6.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i15_LC_17_6_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i15_LC_17_6_6 (
            .in0(N__48504),
            .in1(N__47992),
            .in2(_gnd_net_),
            .in3(N__47977),
            .lcout(wdtick_cnt_14),
            .ltout(),
            .carryin(n20779),
            .carryout(n20780),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i16_LC_17_6_7.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i16_LC_17_6_7.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i16_LC_17_6_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i16_LC_17_6_7 (
            .in0(N__48536),
            .in1(N__47974),
            .in2(_gnd_net_),
            .in3(N__47962),
            .lcout(wdtick_cnt_15),
            .ltout(),
            .carryin(n20780),
            .carryout(n20781),
            .clk(N__48407),
            .ce(N__48338),
            .sr(N__51224));
    defparam wdtick_cnt_3783_3784__i17_LC_17_7_0.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i17_LC_17_7_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i17_LC_17_7_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i17_LC_17_7_0 (
            .in0(N__48537),
            .in1(N__48234),
            .in2(_gnd_net_),
            .in3(N__48220),
            .lcout(wdtick_cnt_16),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(n20782),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i18_LC_17_7_1.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i18_LC_17_7_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i18_LC_17_7_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i18_LC_17_7_1 (
            .in0(N__48506),
            .in1(N__48217),
            .in2(_gnd_net_),
            .in3(N__48205),
            .lcout(wdtick_cnt_17),
            .ltout(),
            .carryin(n20782),
            .carryout(n20783),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i19_LC_17_7_2.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i19_LC_17_7_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i19_LC_17_7_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i19_LC_17_7_2 (
            .in0(N__48538),
            .in1(N__48201),
            .in2(_gnd_net_),
            .in3(N__48187),
            .lcout(wdtick_cnt_18),
            .ltout(),
            .carryin(n20783),
            .carryout(n20784),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i20_LC_17_7_3.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i20_LC_17_7_3.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i20_LC_17_7_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i20_LC_17_7_3 (
            .in0(N__48507),
            .in1(N__48183),
            .in2(_gnd_net_),
            .in3(N__48169),
            .lcout(wdtick_cnt_19),
            .ltout(),
            .carryin(n20784),
            .carryout(n20785),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i21_LC_17_7_4.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i21_LC_17_7_4.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i21_LC_17_7_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i21_LC_17_7_4 (
            .in0(N__48539),
            .in1(N__48166),
            .in2(_gnd_net_),
            .in3(N__48154),
            .lcout(wdtick_cnt_20),
            .ltout(),
            .carryin(n20785),
            .carryout(n20786),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i22_LC_17_7_5.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i22_LC_17_7_5.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i22_LC_17_7_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i22_LC_17_7_5 (
            .in0(N__48508),
            .in1(N__48151),
            .in2(_gnd_net_),
            .in3(N__48139),
            .lcout(wdtick_cnt_21),
            .ltout(),
            .carryin(n20786),
            .carryout(n20787),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i23_LC_17_7_6.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i23_LC_17_7_6.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i23_LC_17_7_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i23_LC_17_7_6 (
            .in0(N__48540),
            .in1(N__48136),
            .in2(_gnd_net_),
            .in3(N__48124),
            .lcout(wdtick_cnt_22),
            .ltout(),
            .carryin(n20787),
            .carryout(n20788),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i24_LC_17_7_7.C_ON=1'b1;
    defparam wdtick_cnt_3783_3784__i24_LC_17_7_7.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i24_LC_17_7_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3783_3784__i24_LC_17_7_7 (
            .in0(N__48509),
            .in1(N__48121),
            .in2(_gnd_net_),
            .in3(N__48109),
            .lcout(wdtick_cnt_23),
            .ltout(),
            .carryin(n20788),
            .carryout(n20789),
            .clk(N__48408),
            .ce(N__48337),
            .sr(N__51219));
    defparam wdtick_cnt_3783_3784__i25_LC_17_8_0.C_ON=1'b0;
    defparam wdtick_cnt_3783_3784__i25_LC_17_8_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3783_3784__i25_LC_17_8_0.LUT_INIT=16'b1000010001001000;
    LogicCell40 wdtick_cnt_3783_3784__i25_LC_17_8_0 (
            .in0(N__48435),
            .in1(N__48532),
            .in2(_gnd_net_),
            .in3(N__48439),
            .lcout(wdtick_cnt_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48410),
            .ce(N__48345),
            .sr(N__51223));
    defparam i2_2_lut_4_lut_LC_17_9_0.C_ON=1'b0;
    defparam i2_2_lut_4_lut_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam i2_2_lut_4_lut_LC_17_9_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 i2_2_lut_4_lut_LC_17_9_0 (
            .in0(N__51168),
            .in1(N__51784),
            .in2(N__62608),
            .in3(N__57353),
            .lcout(n7_adj_1757),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i1_LC_17_9_1.C_ON=1'b0;
    defparam comm_index_i1_LC_17_9_1.SEQ_MODE=4'b1000;
    defparam comm_index_i1_LC_17_9_1.LUT_INIT=16'b1101001011110000;
    LogicCell40 comm_index_i1_LC_17_9_1 (
            .in0(N__58042),
            .in1(N__58208),
            .in2(N__51808),
            .in3(N__54310),
            .lcout(comm_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61865),
            .ce(N__48262),
            .sr(N__48292));
    defparam i462_2_lut_LC_17_9_2.C_ON=1'b0;
    defparam i462_2_lut_LC_17_9_2.SEQ_MODE=4'b0000;
    defparam i462_2_lut_LC_17_9_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 i462_2_lut_LC_17_9_2 (
            .in0(N__58209),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58040),
            .lcout(n2562),
            .ltout(n2562_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i2_LC_17_9_3.C_ON=1'b0;
    defparam comm_index_i2_LC_17_9_3.SEQ_MODE=4'b1000;
    defparam comm_index_i2_LC_17_9_3.LUT_INIT=16'b0111111110000000;
    LogicCell40 comm_index_i2_LC_17_9_3 (
            .in0(N__51785),
            .in1(N__54309),
            .in2(N__48295),
            .in3(N__54572),
            .lcout(comm_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61865),
            .ce(N__48262),
            .sr(N__48292));
    defparam comm_index_i0_LC_17_9_4.C_ON=1'b0;
    defparam comm_index_i0_LC_17_9_4.SEQ_MODE=4'b1000;
    defparam comm_index_i0_LC_17_9_4.LUT_INIT=16'b1001100111001100;
    LogicCell40 comm_index_i0_LC_17_9_4 (
            .in0(N__58207),
            .in1(N__54308),
            .in2(_gnd_net_),
            .in3(N__58041),
            .lcout(comm_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61865),
            .ce(N__48262),
            .sr(N__48292));
    defparam i3_3_lut_4_lut_adj_284_LC_17_9_5.C_ON=1'b0;
    defparam i3_3_lut_4_lut_adj_284_LC_17_9_5.SEQ_MODE=4'b0000;
    defparam i3_3_lut_4_lut_adj_284_LC_17_9_5.LUT_INIT=16'b0000000001000000;
    LogicCell40 i3_3_lut_4_lut_adj_284_LC_17_9_5 (
            .in0(N__61381),
            .in1(N__60006),
            .in2(N__64066),
            .in3(N__63505),
            .lcout(n8_adj_1782),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_286_LC_17_9_6.C_ON=1'b0;
    defparam i1_3_lut_adj_286_LC_17_9_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_286_LC_17_9_6.LUT_INIT=16'b1110111000000000;
    LogicCell40 i1_3_lut_adj_286_LC_17_9_6 (
            .in0(N__63504),
            .in1(N__51175),
            .in2(_gnd_net_),
            .in3(N__63204),
            .lcout(n12540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_78_LC_17_9_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_78_LC_17_9_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_78_LC_17_9_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i1_2_lut_3_lut_adj_78_LC_17_9_7 (
            .in0(N__64034),
            .in1(N__49087),
            .in2(_gnd_net_),
            .in3(N__62449),
            .lcout(n14_adj_1606),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19313_4_lut_LC_17_10_0.C_ON=1'b0;
    defparam i19313_4_lut_LC_17_10_0.SEQ_MODE=4'b0000;
    defparam i19313_4_lut_LC_17_10_0.LUT_INIT=16'b1111101011011000;
    LogicCell40 i19313_4_lut_LC_17_10_0 (
            .in0(N__64023),
            .in1(N__53439),
            .in2(N__48673),
            .in3(N__48655),
            .lcout(),
            .ltout(n22240_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i0_LC_17_10_1.C_ON=1'b0;
    defparam comm_state_i0_LC_17_10_1.SEQ_MODE=4'b1000;
    defparam comm_state_i0_LC_17_10_1.LUT_INIT=16'b0011001111110000;
    LogicCell40 comm_state_i0_LC_17_10_1 (
            .in0(_gnd_net_),
            .in1(N__57739),
            .in2(N__48658),
            .in3(N__63494),
            .lcout(comm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61878),
            .ce(N__51235),
            .sr(_gnd_net_));
    defparam i20126_3_lut_LC_17_10_2.C_ON=1'b0;
    defparam i20126_3_lut_LC_17_10_2.SEQ_MODE=4'b0000;
    defparam i20126_3_lut_LC_17_10_2.LUT_INIT=16'b1010101010001000;
    LogicCell40 i20126_3_lut_LC_17_10_2 (
            .in0(N__62572),
            .in1(N__57300),
            .in2(_gnd_net_),
            .in3(N__51169),
            .lcout(n23053),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12533_2_lut_LC_17_10_4.C_ON=1'b0;
    defparam i12533_2_lut_LC_17_10_4.SEQ_MODE=4'b0000;
    defparam i12533_2_lut_LC_17_10_4.LUT_INIT=16'b1100110011111111;
    LogicCell40 i12533_2_lut_LC_17_10_4 (
            .in0(_gnd_net_),
            .in1(N__58153),
            .in2(_gnd_net_),
            .in3(N__62930),
            .lcout(n15261),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_128_LC_17_10_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_128_LC_17_10_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_128_LC_17_10_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_2_lut_3_lut_adj_128_LC_17_10_5 (
            .in0(N__62931),
            .in1(N__62570),
            .in2(_gnd_net_),
            .in3(N__64022),
            .lcout(),
            .ltout(n11280_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_228_LC_17_10_6.C_ON=1'b0;
    defparam i1_4_lut_adj_228_LC_17_10_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_228_LC_17_10_6.LUT_INIT=16'b1000110010101111;
    LogicCell40 i1_4_lut_adj_228_LC_17_10_6 (
            .in0(N__63492),
            .in1(N__63145),
            .in2(N__48649),
            .in3(N__56247),
            .lcout(n12509),
            .ltout(n12509_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_114_LC_17_10_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_114_LC_17_10_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_114_LC_17_10_7.LUT_INIT=16'b0001111100001111;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_114_LC_17_10_7 (
            .in0(N__64024),
            .in1(N__62571),
            .in2(N__48646),
            .in3(N__63493),
            .lcout(n18363),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_86_LC_17_11_0.C_ON=1'b0;
    defparam i1_4_lut_adj_86_LC_17_11_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_86_LC_17_11_0.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_86_LC_17_11_0 (
            .in0(N__54312),
            .in1(N__48643),
            .in2(N__48628),
            .in3(N__54537),
            .lcout(n4_adj_1745),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23486_bdd_4_lut_LC_17_11_1.C_ON=1'b0;
    defparam n23486_bdd_4_lut_LC_17_11_1.SEQ_MODE=4'b0000;
    defparam n23486_bdd_4_lut_LC_17_11_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 n23486_bdd_4_lut_LC_17_11_1 (
            .in0(N__48609),
            .in1(N__48586),
            .in2(N__48574),
            .in3(N__60309),
            .lcout(n22180),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_311_LC_17_11_2.C_ON=1'b0;
    defparam i1_2_lut_adj_311_LC_17_11_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_311_LC_17_11_2.LUT_INIT=16'b0000000011110000;
    LogicCell40 i1_2_lut_adj_311_LC_17_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51133),
            .in3(N__54538),
            .lcout(n4_adj_1749),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19973_2_lut_4_lut_LC_17_11_3.C_ON=1'b0;
    defparam i19973_2_lut_4_lut_LC_17_11_3.SEQ_MODE=4'b0000;
    defparam i19973_2_lut_4_lut_LC_17_11_3.LUT_INIT=16'b1111010111110111;
    LogicCell40 i19973_2_lut_4_lut_LC_17_11_3 (
            .in0(N__58650),
            .in1(N__60314),
            .in2(N__50885),
            .in3(N__59015),
            .lcout(n22330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i50_4_lut_LC_17_11_4.C_ON=1'b0;
    defparam i50_4_lut_LC_17_11_4.SEQ_MODE=4'b0000;
    defparam i50_4_lut_LC_17_11_4.LUT_INIT=16'b0011101101010000;
    LogicCell40 i50_4_lut_LC_17_11_4 (
            .in0(N__59014),
            .in1(N__59867),
            .in2(N__60463),
            .in3(N__60990),
            .lcout(),
            .ltout(n46_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19794_4_lut_LC_17_11_5.C_ON=1'b0;
    defparam i19794_4_lut_LC_17_11_5.SEQ_MODE=4'b0000;
    defparam i19794_4_lut_LC_17_11_5.LUT_INIT=16'b0101000001010001;
    LogicCell40 i19794_4_lut_LC_17_11_5 (
            .in0(N__58649),
            .in1(N__59887),
            .in2(N__48997),
            .in3(N__60313),
            .lcout(n22353),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_0_i111_3_lut_LC_17_11_6.C_ON=1'b0;
    defparam mux_126_Mux_0_i111_3_lut_LC_17_11_6.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_0_i111_3_lut_LC_17_11_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_126_Mux_0_i111_3_lut_LC_17_11_6 (
            .in0(N__59016),
            .in1(_gnd_net_),
            .in2(N__48994),
            .in3(N__48964),
            .lcout(n111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_323_LC_17_11_7.C_ON=1'b0;
    defparam i1_2_lut_adj_323_LC_17_11_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_323_LC_17_11_7.LUT_INIT=16'b0100010001000100;
    LogicCell40 i1_2_lut_adj_323_LC_17_11_7 (
            .in0(N__62905),
            .in1(N__54311),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16444_2_lut_3_lut_LC_17_12_0.C_ON=1'b0;
    defparam i16444_2_lut_3_lut_LC_17_12_0.SEQ_MODE=4'b0000;
    defparam i16444_2_lut_3_lut_LC_17_12_0.LUT_INIT=16'b0000000001000100;
    LogicCell40 i16444_2_lut_3_lut_LC_17_12_0 (
            .in0(N__62567),
            .in1(N__49273),
            .in2(_gnd_net_),
            .in3(N__64030),
            .lcout(n14_adj_1662),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_312_LC_17_12_1.C_ON=1'b0;
    defparam i19_4_lut_adj_312_LC_17_12_1.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_312_LC_17_12_1.LUT_INIT=16'b1101000100010001;
    LogicCell40 i19_4_lut_adj_312_LC_17_12_1 (
            .in0(N__51623),
            .in1(N__62565),
            .in2(N__49362),
            .in3(N__48900),
            .lcout(n12_adj_1684),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i0_LC_17_12_2.C_ON=1'b0;
    defparam buf_cfgRTD_i0_LC_17_12_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i0_LC_17_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i0_LC_17_12_2 (
            .in0(N__48880),
            .in1(N__48798),
            .in2(_gnd_net_),
            .in3(N__48692),
            .lcout(buf_cfgRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61906),
            .ce(),
            .sr(_gnd_net_));
    defparam i16282_2_lut_LC_17_12_3.C_ON=1'b0;
    defparam i16282_2_lut_LC_17_12_3.SEQ_MODE=4'b0000;
    defparam i16282_2_lut_LC_17_12_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i16282_2_lut_LC_17_12_3 (
            .in0(_gnd_net_),
            .in1(N__58515),
            .in2(_gnd_net_),
            .in3(N__58625),
            .lcout(n7148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_297_LC_17_12_4.C_ON=1'b0;
    defparam i1_2_lut_adj_297_LC_17_12_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_297_LC_17_12_4.LUT_INIT=16'b0000000010101010;
    LogicCell40 i1_2_lut_adj_297_LC_17_12_4 (
            .in0(N__58626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59936),
            .lcout(),
            .ltout(n4_adj_1709_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i45_4_lut_LC_17_12_5.C_ON=1'b0;
    defparam i45_4_lut_LC_17_12_5.SEQ_MODE=4'b0000;
    defparam i45_4_lut_LC_17_12_5.LUT_INIT=16'b1010000011001100;
    LogicCell40 i45_4_lut_LC_17_12_5 (
            .in0(N__49372),
            .in1(N__58399),
            .in2(N__49366),
            .in3(N__61379),
            .lcout(n30_adj_1720),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19163_2_lut_LC_17_12_6.C_ON=1'b0;
    defparam i19163_2_lut_LC_17_12_6.SEQ_MODE=4'b0000;
    defparam i19163_2_lut_LC_17_12_6.LUT_INIT=16'b1111111110101010;
    LogicCell40 i19163_2_lut_LC_17_12_6 (
            .in0(N__54326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62943),
            .lcout(n22089),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_330_LC_17_12_7.C_ON=1'b0;
    defparam i19_4_lut_adj_330_LC_17_12_7.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_330_LC_17_12_7.LUT_INIT=16'b1101000100010001;
    LogicCell40 i19_4_lut_adj_330_LC_17_12_7 (
            .in0(N__51624),
            .in1(N__62566),
            .in2(N__49363),
            .in3(N__51585),
            .lcout(n12_adj_1802),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i3_LC_17_13_0.C_ON=1'b0;
    defparam comm_buf_1__i3_LC_17_13_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i3_LC_17_13_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_1__i3_LC_17_13_0 (
            .in0(N__62598),
            .in1(N__62788),
            .in2(_gnd_net_),
            .in3(N__49342),
            .lcout(comm_buf_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61920),
            .ce(N__55769),
            .sr(N__55707));
    defparam comm_buf_1__i6_LC_17_13_1.C_ON=1'b0;
    defparam comm_buf_1__i6_LC_17_13_1.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i6_LC_17_13_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i6_LC_17_13_1 (
            .in0(N__53883),
            .in1(N__62599),
            .in2(_gnd_net_),
            .in3(N__49615),
            .lcout(comm_buf_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61920),
            .ce(N__55769),
            .sr(N__55707));
    defparam comm_buf_1__i0_LC_17_13_2.C_ON=1'b0;
    defparam comm_buf_1__i0_LC_17_13_2.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i0_LC_17_13_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_1__i0_LC_17_13_2 (
            .in0(N__62597),
            .in1(N__54023),
            .in2(_gnd_net_),
            .in3(N__51655),
            .lcout(comm_buf_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61920),
            .ce(N__55769),
            .sr(N__55707));
    defparam i19785_2_lut_LC_17_13_5.C_ON=1'b0;
    defparam i19785_2_lut_LC_17_13_5.SEQ_MODE=4'b0000;
    defparam i19785_2_lut_LC_17_13_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i19785_2_lut_LC_17_13_5 (
            .in0(_gnd_net_),
            .in1(N__49030),
            .in2(_gnd_net_),
            .in3(N__59191),
            .lcout(n22296),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19894_2_lut_LC_17_13_6.C_ON=1'b0;
    defparam i19894_2_lut_LC_17_13_6.SEQ_MODE=4'b0000;
    defparam i19894_2_lut_LC_17_13_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i19894_2_lut_LC_17_13_6 (
            .in0(N__59192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49723),
            .lcout(n22499),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23516_bdd_4_lut_LC_17_14_0.C_ON=1'b0;
    defparam n23516_bdd_4_lut_LC_17_14_0.SEQ_MODE=4'b0000;
    defparam n23516_bdd_4_lut_LC_17_14_0.LUT_INIT=16'b1111110000100010;
    LogicCell40 n23516_bdd_4_lut_LC_17_14_0 (
            .in0(N__49690),
            .in1(N__59978),
            .in2(N__49669),
            .in3(N__49588),
            .lcout(),
            .ltout(n23519_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1668899_i1_3_lut_LC_17_14_1.C_ON=1'b0;
    defparam i1668899_i1_3_lut_LC_17_14_1.SEQ_MODE=4'b0000;
    defparam i1668899_i1_3_lut_LC_17_14_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 i1668899_i1_3_lut_LC_17_14_1 (
            .in0(N__60976),
            .in1(_gnd_net_),
            .in2(N__49642),
            .in3(N__49639),
            .lcout(),
            .ltout(n30_adj_1724_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_6_i127_3_lut_LC_17_14_2.C_ON=1'b0;
    defparam mux_126_Mux_6_i127_3_lut_LC_17_14_2.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_6_i127_3_lut_LC_17_14_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_126_Mux_6_i127_3_lut_LC_17_14_2 (
            .in0(_gnd_net_),
            .in1(N__49627),
            .in2(N__49618),
            .in3(N__61383),
            .lcout(comm_buf_1_7_N_559_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_6_i26_3_lut_LC_17_14_3.C_ON=1'b0;
    defparam mux_126_Mux_6_i26_3_lut_LC_17_14_3.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_6_i26_3_lut_LC_17_14_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_126_Mux_6_i26_3_lut_LC_17_14_3 (
            .in0(N__49609),
            .in1(N__59502),
            .in2(_gnd_net_),
            .in3(N__49778),
            .lcout(),
            .ltout(n26_adj_1723_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20572_LC_17_14_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20572_LC_17_14_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20572_LC_17_14_4.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20572_LC_17_14_4 (
            .in0(N__55441),
            .in1(N__59977),
            .in2(N__49591),
            .in3(N__60603),
            .lcout(n23516),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16700105_i1_3_lut_LC_17_14_5.C_ON=1'b0;
    defparam i16700105_i1_3_lut_LC_17_14_5.SEQ_MODE=4'b0000;
    defparam i16700105_i1_3_lut_LC_17_14_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 i16700105_i1_3_lut_LC_17_14_5 (
            .in0(N__60975),
            .in1(N__49582),
            .in2(_gnd_net_),
            .in3(N__49576),
            .lcout(n30_adj_1579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i4_LC_17_14_6.C_ON=1'b0;
    defparam buf_dds1_i4_LC_17_14_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i4_LC_17_14_6.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i4_LC_17_14_6 (
            .in0(N__49457),
            .in1(N__55381),
            .in2(N__56086),
            .in3(N__49502),
            .lcout(buf_dds1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61940),
            .ce(),
            .sr(_gnd_net_));
    defparam data_cntvec_i0_i0_LC_17_15_0.C_ON=1'b1;
    defparam data_cntvec_i0_i0_LC_17_15_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i0_LC_17_15_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i0_LC_17_15_0 (
            .in0(_gnd_net_),
            .in1(N__49392),
            .in2(N__49438),
            .in3(_gnd_net_),
            .lcout(data_cntvec_0),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(n20622),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i1_LC_17_15_1.C_ON=1'b1;
    defparam data_cntvec_i0_i1_LC_17_15_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i1_LC_17_15_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i1_LC_17_15_1 (
            .in0(_gnd_net_),
            .in1(N__52257),
            .in2(_gnd_net_),
            .in3(N__49825),
            .lcout(data_cntvec_1),
            .ltout(),
            .carryin(n20622),
            .carryout(n20623),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i2_LC_17_15_2.C_ON=1'b1;
    defparam data_cntvec_i0_i2_LC_17_15_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i2_LC_17_15_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i2_LC_17_15_2 (
            .in0(_gnd_net_),
            .in1(N__52398),
            .in2(_gnd_net_),
            .in3(N__49822),
            .lcout(data_cntvec_2),
            .ltout(),
            .carryin(n20623),
            .carryout(n20624),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i3_LC_17_15_3.C_ON=1'b1;
    defparam data_cntvec_i0_i3_LC_17_15_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i3_LC_17_15_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i3_LC_17_15_3 (
            .in0(_gnd_net_),
            .in1(N__49815),
            .in2(_gnd_net_),
            .in3(N__49795),
            .lcout(data_cntvec_3),
            .ltout(),
            .carryin(n20624),
            .carryout(n20625),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i4_LC_17_15_4.C_ON=1'b1;
    defparam data_cntvec_i0_i4_LC_17_15_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i4_LC_17_15_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i4_LC_17_15_4 (
            .in0(_gnd_net_),
            .in1(N__52545),
            .in2(_gnd_net_),
            .in3(N__49792),
            .lcout(data_cntvec_4),
            .ltout(),
            .carryin(n20625),
            .carryout(n20626),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i5_LC_17_15_5.C_ON=1'b1;
    defparam data_cntvec_i0_i5_LC_17_15_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i5_LC_17_15_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i5_LC_17_15_5 (
            .in0(_gnd_net_),
            .in1(N__51980),
            .in2(_gnd_net_),
            .in3(N__49789),
            .lcout(data_cntvec_5),
            .ltout(),
            .carryin(n20626),
            .carryout(n20627),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i6_LC_17_15_6.C_ON=1'b1;
    defparam data_cntvec_i0_i6_LC_17_15_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i6_LC_17_15_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i6_LC_17_15_6 (
            .in0(_gnd_net_),
            .in1(N__49782),
            .in2(_gnd_net_),
            .in3(N__49762),
            .lcout(data_cntvec_6),
            .ltout(),
            .carryin(n20627),
            .carryout(n20628),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i7_LC_17_15_7.C_ON=1'b1;
    defparam data_cntvec_i0_i7_LC_17_15_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i7_LC_17_15_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i7_LC_17_15_7 (
            .in0(_gnd_net_),
            .in1(N__54650),
            .in2(_gnd_net_),
            .in3(N__49759),
            .lcout(data_cntvec_7),
            .ltout(),
            .carryin(n20628),
            .carryout(n20629),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__50018),
            .sr(N__49942));
    defparam data_cntvec_i0_i8_LC_17_16_0.C_ON=1'b1;
    defparam data_cntvec_i0_i8_LC_17_16_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i8_LC_17_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i8_LC_17_16_0 (
            .in0(_gnd_net_),
            .in1(N__49746),
            .in2(_gnd_net_),
            .in3(N__49726),
            .lcout(data_cntvec_8),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(n20630),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam data_cntvec_i0_i9_LC_17_16_1.C_ON=1'b1;
    defparam data_cntvec_i0_i9_LC_17_16_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i9_LC_17_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i9_LC_17_16_1 (
            .in0(_gnd_net_),
            .in1(N__50937),
            .in2(_gnd_net_),
            .in3(N__50131),
            .lcout(data_cntvec_9),
            .ltout(),
            .carryin(n20630),
            .carryout(n20631),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam data_cntvec_i0_i10_LC_17_16_2.C_ON=1'b1;
    defparam data_cntvec_i0_i10_LC_17_16_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i10_LC_17_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i10_LC_17_16_2 (
            .in0(_gnd_net_),
            .in1(N__50117),
            .in2(_gnd_net_),
            .in3(N__50092),
            .lcout(data_cntvec_10),
            .ltout(),
            .carryin(n20631),
            .carryout(n20632),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam data_cntvec_i0_i11_LC_17_16_3.C_ON=1'b1;
    defparam data_cntvec_i0_i11_LC_17_16_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i11_LC_17_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i11_LC_17_16_3 (
            .in0(_gnd_net_),
            .in1(N__56132),
            .in2(_gnd_net_),
            .in3(N__50089),
            .lcout(data_cntvec_11),
            .ltout(),
            .carryin(n20632),
            .carryout(n20633),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam data_cntvec_i0_i12_LC_17_16_4.C_ON=1'b1;
    defparam data_cntvec_i0_i12_LC_17_16_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i12_LC_17_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i12_LC_17_16_4 (
            .in0(_gnd_net_),
            .in1(N__50082),
            .in2(_gnd_net_),
            .in3(N__50068),
            .lcout(data_cntvec_12),
            .ltout(),
            .carryin(n20633),
            .carryout(n20634),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam data_cntvec_i0_i13_LC_17_16_5.C_ON=1'b1;
    defparam data_cntvec_i0_i13_LC_17_16_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i13_LC_17_16_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i13_LC_17_16_5 (
            .in0(_gnd_net_),
            .in1(N__50058),
            .in2(_gnd_net_),
            .in3(N__50044),
            .lcout(data_cntvec_13),
            .ltout(),
            .carryin(n20634),
            .carryout(n20635),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam data_cntvec_i0_i14_LC_17_16_6.C_ON=1'b1;
    defparam data_cntvec_i0_i14_LC_17_16_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i14_LC_17_16_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i14_LC_17_16_6 (
            .in0(_gnd_net_),
            .in1(N__51699),
            .in2(_gnd_net_),
            .in3(N__50041),
            .lcout(data_cntvec_14),
            .ltout(),
            .carryin(n20635),
            .carryout(n20636),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam data_cntvec_i0_i15_LC_17_16_7.C_ON=1'b0;
    defparam data_cntvec_i0_i15_LC_17_16_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i15_LC_17_16_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i15_LC_17_16_7 (
            .in0(_gnd_net_),
            .in1(N__50034),
            .in2(_gnd_net_),
            .in3(N__50038),
            .lcout(data_cntvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__50017),
            .sr(N__49943));
    defparam n23480_bdd_4_lut_LC_17_17_0.C_ON=1'b0;
    defparam n23480_bdd_4_lut_LC_17_17_0.SEQ_MODE=4'b0000;
    defparam n23480_bdd_4_lut_LC_17_17_0.LUT_INIT=16'b1011101010011000;
    LogicCell40 n23480_bdd_4_lut_LC_17_17_0 (
            .in0(N__49909),
            .in1(N__60592),
            .in2(N__49884),
            .in3(N__49852),
            .lcout(),
            .ltout(n22183_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_20528_LC_17_17_1.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_20528_LC_17_17_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_20528_LC_17_17_1.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_2__bdd_4_lut_20528_LC_17_17_1 (
            .in0(N__61022),
            .in1(N__60059),
            .in2(N__49828),
            .in3(N__50899),
            .lcout(),
            .ltout(n23462_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23462_bdd_4_lut_LC_17_17_2.C_ON=1'b0;
    defparam n23462_bdd_4_lut_LC_17_17_2.SEQ_MODE=4'b0000;
    defparam n23462_bdd_4_lut_LC_17_17_2.LUT_INIT=16'b1111000011001010;
    LogicCell40 n23462_bdd_4_lut_LC_17_17_2 (
            .in0(N__50986),
            .in1(N__50977),
            .in2(N__50968),
            .in3(N__61023),
            .lcout(n23465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19257_3_lut_LC_17_17_3.C_ON=1'b0;
    defparam i19257_3_lut_LC_17_17_3.SEQ_MODE=4'b0000;
    defparam i19257_3_lut_LC_17_17_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 i19257_3_lut_LC_17_17_3 (
            .in0(N__50949),
            .in1(N__59408),
            .in2(_gnd_net_),
            .in3(N__50933),
            .lcout(),
            .ltout(n22184_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19259_4_lut_LC_17_17_4.C_ON=1'b0;
    defparam i19259_4_lut_LC_17_17_4.SEQ_MODE=4'b0000;
    defparam i19259_4_lut_LC_17_17_4.LUT_INIT=16'b1110111011110000;
    LogicCell40 i19259_4_lut_LC_17_17_4 (
            .in0(N__59409),
            .in1(N__50917),
            .in2(N__50902),
            .in3(N__60591),
            .lcout(n22186),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_285_LC_17_17_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_285_LC_17_17_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_285_LC_17_17_6.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_285_LC_17_17_6 (
            .in0(N__60058),
            .in1(N__58528),
            .in2(_gnd_net_),
            .in3(N__61021),
            .lcout(n21997),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i9_LC_17_18_3.C_ON=1'b0;
    defparam buf_dds0_i9_LC_17_18_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i9_LC_17_18_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 buf_dds0_i9_LC_17_18_3 (
            .in0(N__50807),
            .in1(N__50633),
            .in2(_gnd_net_),
            .in3(N__50775),
            .lcout(buf_dds0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61998),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.CS_28_LC_17_20_7 .C_ON=1'b0;
    defparam \SIG_DDS.CS_28_LC_17_20_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.CS_28_LC_17_20_7 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \SIG_DDS.CS_28_LC_17_20_7  (
            .in0(N__50608),
            .in1(N__50538),
            .in2(_gnd_net_),
            .in3(N__50329),
            .lcout(DDS_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__62008),
            .ce(N__50245),
            .sr(_gnd_net_));
    defparam i20042_2_lut_LC_18_3_7.C_ON=1'b0;
    defparam i20042_2_lut_LC_18_3_7.SEQ_MODE=4'b0000;
    defparam i20042_2_lut_LC_18_3_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i20042_2_lut_LC_18_3_7 (
            .in0(_gnd_net_),
            .in1(N__50233),
            .in2(_gnd_net_),
            .in3(N__59427),
            .lcout(n22595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_18_4_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_18_4_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_18_4_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_88_2_lut_LC_18_4_2  (
            .in0(N__50168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57077),
            .lcout(\comm_spi.imosi_N_840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_12628_12629_reset_LC_18_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12628_12629_reset_LC_18_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i3_12628_12629_reset_LC_18_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_12628_12629_reset_LC_18_7_0  (
            .in0(N__51124),
            .in1(N__51103),
            .in2(_gnd_net_),
            .in3(N__51079),
            .lcout(\comm_spi.n15357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53670),
            .ce(),
            .sr(N__51022));
    defparam i19790_2_lut_LC_18_8_0.C_ON=1'b0;
    defparam i19790_2_lut_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam i19790_2_lut_LC_18_8_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19790_2_lut_LC_18_8_0 (
            .in0(_gnd_net_),
            .in1(N__56871),
            .in2(_gnd_net_),
            .in3(N__63030),
            .lcout(),
            .ltout(n22489_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i3_LC_18_8_1.C_ON=1'b0;
    defparam comm_state_i3_LC_18_8_1.SEQ_MODE=4'b1000;
    defparam comm_state_i3_LC_18_8_1.LUT_INIT=16'b0010000001110101;
    LogicCell40 comm_state_i3_LC_18_8_1 (
            .in0(N__63358),
            .in1(N__57521),
            .in2(N__51004),
            .in3(N__50992),
            .lcout(comm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61866),
            .ce(N__50998),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_18_8_2.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_18_8_2.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_18_8_2.LUT_INIT=16'b1111101111111111;
    LogicCell40 i2_3_lut_4_lut_LC_18_8_2 (
            .in0(N__62485),
            .in1(N__63029),
            .in2(N__54183),
            .in3(N__57354),
            .lcout(),
            .ltout(n20959_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_88_LC_18_8_3.C_ON=1'b0;
    defparam i1_4_lut_adj_88_LC_18_8_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_88_LC_18_8_3.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_adj_88_LC_18_8_3 (
            .in0(N__57970),
            .in1(N__51566),
            .in2(N__51001),
            .in3(N__53349),
            .lcout(n21883),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_70_LC_18_8_4.C_ON=1'b0;
    defparam i1_2_lut_adj_70_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_70_LC_18_8_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_70_LC_18_8_4 (
            .in0(_gnd_net_),
            .in1(N__64006),
            .in2(_gnd_net_),
            .in3(N__63357),
            .lcout(n12951),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_346_Mux_3_i7_4_lut_LC_18_8_6.C_ON=1'b0;
    defparam comm_state_3__I_0_346_Mux_3_i7_4_lut_LC_18_8_6.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_346_Mux_3_i7_4_lut_LC_18_8_6.LUT_INIT=16'b1101110111110000;
    LogicCell40 comm_state_3__I_0_346_Mux_3_i7_4_lut_LC_18_8_6 (
            .in0(N__62486),
            .in1(N__51406),
            .in2(N__53416),
            .in3(N__64007),
            .lcout(n19241),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19824_2_lut_3_lut_LC_18_9_0.C_ON=1'b0;
    defparam i19824_2_lut_3_lut_LC_18_9_0.SEQ_MODE=4'b0000;
    defparam i19824_2_lut_3_lut_LC_18_9_0.LUT_INIT=16'b0000000001000100;
    LogicCell40 i19824_2_lut_3_lut_LC_18_9_0 (
            .in0(N__58117),
            .in1(N__62421),
            .in2(_gnd_net_),
            .in3(N__58036),
            .lcout(n22339),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_LC_18_9_1.C_ON=1'b0;
    defparam i2_4_lut_4_lut_LC_18_9_1.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_LC_18_9_1.LUT_INIT=16'b0100111111101111;
    LogicCell40 i2_4_lut_4_lut_LC_18_9_1 (
            .in0(N__58037),
            .in1(N__58118),
            .in2(N__62601),
            .in3(N__62933),
            .lcout(n22033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_304_LC_18_9_2.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_304_LC_18_9_2.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_304_LC_18_9_2.LUT_INIT=16'b1111111011111111;
    LogicCell40 i2_3_lut_4_lut_adj_304_LC_18_9_2 (
            .in0(N__53438),
            .in1(N__62427),
            .in2(N__54184),
            .in3(N__58038),
            .lcout(),
            .ltout(n12064_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_143_LC_18_9_3.C_ON=1'b0;
    defparam i1_4_lut_adj_143_LC_18_9_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_143_LC_18_9_3.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_adj_143_LC_18_9_3 (
            .in0(N__51244),
            .in1(N__51567),
            .in2(N__51238),
            .in3(N__53350),
            .lcout(n21885),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19147_2_lut_LC_18_9_4.C_ON=1'b0;
    defparam i19147_2_lut_LC_18_9_4.SEQ_MODE=4'b0000;
    defparam i19147_2_lut_LC_18_9_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 i19147_2_lut_LC_18_9_4 (
            .in0(N__62934),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62426),
            .lcout(),
            .ltout(n22073_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_224_LC_18_9_5.C_ON=1'b0;
    defparam i1_4_lut_adj_224_LC_18_9_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_224_LC_18_9_5.LUT_INIT=16'b1100110000000100;
    LogicCell40 i1_4_lut_adj_224_LC_18_9_5 (
            .in0(N__64011),
            .in1(N__63173),
            .in2(N__51229),
            .in3(N__63378),
            .lcout(n12050),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam flagcntwd_306_LC_18_9_6.C_ON=1'b0;
    defparam flagcntwd_306_LC_18_9_6.SEQ_MODE=4'b1000;
    defparam flagcntwd_306_LC_18_9_6.LUT_INIT=16'b1111111101010101;
    LogicCell40 flagcntwd_306_LC_18_9_6 (
            .in0(N__62935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62428),
            .lcout(flagcntwd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61879),
            .ce(N__51184),
            .sr(N__51645));
    defparam i17_3_lut_3_lut_LC_18_9_7.C_ON=1'b0;
    defparam i17_3_lut_3_lut_LC_18_9_7.SEQ_MODE=4'b0000;
    defparam i17_3_lut_3_lut_LC_18_9_7.LUT_INIT=16'b0000010110100000;
    LogicCell40 i17_3_lut_3_lut_LC_18_9_7 (
            .in0(N__62422),
            .in1(_gnd_net_),
            .in2(N__64050),
            .in3(N__62932),
            .lcout(n10_adj_1602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_106_LC_18_10_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_106_LC_18_10_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_106_LC_18_10_0.LUT_INIT=16'b0000000100000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_106_LC_18_10_0 (
            .in0(N__51780),
            .in1(N__51166),
            .in2(N__58181),
            .in3(N__58018),
            .lcout(n21956),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_107_LC_18_10_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_107_LC_18_10_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_107_LC_18_10_1.LUT_INIT=16'b0001000000000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_107_LC_18_10_1 (
            .in0(N__51167),
            .in1(N__58151),
            .in2(N__58039),
            .in3(N__51779),
            .lcout(n29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12123_2_lut_LC_18_10_2.C_ON=1'b0;
    defparam i12123_2_lut_LC_18_10_2.SEQ_MODE=4'b0000;
    defparam i12123_2_lut_LC_18_10_2.LUT_INIT=16'b1110111011101110;
    LogicCell40 i12123_2_lut_LC_18_10_2 (
            .in0(N__62569),
            .in1(N__62906),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n14851),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_3_lut_LC_18_10_3.C_ON=1'b0;
    defparam i3_3_lut_LC_18_10_3.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_18_10_3.LUT_INIT=16'b1111111111011101;
    LogicCell40 i3_3_lut_LC_18_10_3 (
            .in0(N__58152),
            .in1(N__62568),
            .in2(_gnd_net_),
            .in3(N__51568),
            .lcout(n21981),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_132_LC_18_10_4.C_ON=1'b0;
    defparam i1_4_lut_adj_132_LC_18_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_132_LC_18_10_4.LUT_INIT=16'b1111111110111000;
    LogicCell40 i1_4_lut_adj_132_LC_18_10_4 (
            .in0(N__53398),
            .in1(N__63985),
            .in2(N__51547),
            .in3(N__63613),
            .lcout(n11_adj_1585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i14_LC_18_10_5.C_ON=1'b0;
    defparam req_data_cnt_i14_LC_18_10_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i14_LC_18_10_5.LUT_INIT=16'b1011100010111000;
    LogicCell40 req_data_cnt_i14_LC_18_10_5 (
            .in0(N__51502),
            .in1(N__51283),
            .in2(N__51729),
            .in3(_gnd_net_),
            .lcout(req_data_cnt_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61890),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i2_3_lut_LC_18_10_6 .C_ON=1'b0;
    defparam \comm_spi.i2_3_lut_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i2_3_lut_LC_18_10_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \comm_spi.i2_3_lut_LC_18_10_6  (
            .in0(N__51469),
            .in1(N__51450),
            .in2(_gnd_net_),
            .in3(N__51422),
            .lcout(\comm_spi.n18536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19781_2_lut_3_lut_LC_18_10_7.C_ON=1'b0;
    defparam i19781_2_lut_3_lut_LC_18_10_7.SEQ_MODE=4'b0000;
    defparam i19781_2_lut_3_lut_LC_18_10_7.LUT_INIT=16'b1111111111011101;
    LogicCell40 i19781_2_lut_3_lut_LC_18_10_7 (
            .in0(N__62907),
            .in1(N__58147),
            .in2(_gnd_net_),
            .in3(N__57299),
            .lcout(n22487),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_52_LC_18_11_0.C_ON=1'b0;
    defparam i1_4_lut_adj_52_LC_18_11_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_52_LC_18_11_0.LUT_INIT=16'b1010000010100010;
    LogicCell40 i1_4_lut_adj_52_LC_18_11_0 (
            .in0(N__63393),
            .in1(N__51397),
            .in2(N__57763),
            .in3(N__58369),
            .lcout(n13171),
            .ltout(n13171_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i11_LC_18_11_1.C_ON=1'b0;
    defparam req_data_cnt_i11_LC_18_11_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i11_LC_18_11_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 req_data_cnt_i11_LC_18_11_1 (
            .in0(_gnd_net_),
            .in1(N__57953),
            .in2(N__51247),
            .in3(N__56838),
            .lcout(req_data_cnt_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61907),
            .ce(),
            .sr(_gnd_net_));
    defparam i20051_2_lut_LC_18_11_2.C_ON=1'b0;
    defparam i20051_2_lut_LC_18_11_2.SEQ_MODE=4'b0000;
    defparam i20051_2_lut_LC_18_11_2.LUT_INIT=16'b1111111100110011;
    LogicCell40 i20051_2_lut_LC_18_11_2 (
            .in0(_gnd_net_),
            .in1(N__58526),
            .in2(_gnd_net_),
            .in3(N__58651),
            .lcout(n22329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_326_LC_18_11_3.C_ON=1'b0;
    defparam i1_2_lut_adj_326_LC_18_11_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_326_LC_18_11_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_326_LC_18_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54445),
            .in3(N__54546),
            .lcout(n20318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_130_LC_18_11_4.C_ON=1'b0;
    defparam i1_4_lut_adj_130_LC_18_11_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_130_LC_18_11_4.LUT_INIT=16'b1000100011000000;
    LogicCell40 i1_4_lut_adj_130_LC_18_11_4 (
            .in0(N__51877),
            .in1(N__58527),
            .in2(N__51865),
            .in3(N__61362),
            .lcout(comm_state_3_N_484_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_87_LC_18_11_5.C_ON=1'b0;
    defparam i2_3_lut_adj_87_LC_18_11_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_87_LC_18_11_5.LUT_INIT=16'b1101110111101110;
    LogicCell40 i2_3_lut_adj_87_LC_18_11_5 (
            .in0(N__51856),
            .in1(N__51844),
            .in2(_gnd_net_),
            .in3(N__51807),
            .lcout(n5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_251_LC_18_11_6.C_ON=1'b0;
    defparam i7_4_lut_adj_251_LC_18_11_6.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_251_LC_18_11_6.LUT_INIT=16'b0110111111110110;
    LogicCell40 i7_4_lut_adj_251_LC_18_11_6 (
            .in0(N__51725),
            .in1(N__51703),
            .in2(N__57957),
            .in3(N__56137),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11570_3_lut_LC_18_11_7.C_ON=1'b0;
    defparam i11570_3_lut_LC_18_11_7.SEQ_MODE=4'b0000;
    defparam i11570_3_lut_LC_18_11_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i11570_3_lut_LC_18_11_7 (
            .in0(N__61363),
            .in1(N__51670),
            .in2(_gnd_net_),
            .in3(N__51664),
            .lcout(comm_buf_1_7_N_559_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_82_LC_18_12_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_82_LC_18_12_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_82_LC_18_12_0.LUT_INIT=16'b1110111000000000;
    LogicCell40 i1_2_lut_3_lut_adj_82_LC_18_12_0 (
            .in0(N__62481),
            .in1(N__63994),
            .in2(_gnd_net_),
            .in3(N__63382),
            .lcout(n21271),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_317_LC_18_12_1.C_ON=1'b0;
    defparam i19_4_lut_adj_317_LC_18_12_1.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_317_LC_18_12_1.LUT_INIT=16'b0001101100010001;
    LogicCell40 i19_4_lut_adj_317_LC_18_12_1 (
            .in0(N__62596),
            .in1(N__51625),
            .in2(N__51601),
            .in3(N__51589),
            .lcout(),
            .ltout(n12_adj_1677_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_318_LC_18_12_2.C_ON=1'b0;
    defparam i1_3_lut_adj_318_LC_18_12_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_318_LC_18_12_2.LUT_INIT=16'b1111101000000000;
    LogicCell40 i1_3_lut_adj_318_LC_18_12_2 (
            .in0(N__54160),
            .in1(_gnd_net_),
            .in2(N__51574),
            .in3(N__54066),
            .lcout(n12892),
            .ltout(n12892_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12787_2_lut_LC_18_12_3.C_ON=1'b0;
    defparam i12787_2_lut_LC_18_12_3.SEQ_MODE=4'b0000;
    defparam i12787_2_lut_LC_18_12_3.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12787_2_lut_LC_18_12_3 (
            .in0(N__63381),
            .in1(_gnd_net_),
            .in2(N__51571),
            .in3(_gnd_net_),
            .lcout(n15510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_209_LC_18_12_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_209_LC_18_12_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_209_LC_18_12_4.LUT_INIT=16'b1110111011111111;
    LogicCell40 i1_2_lut_3_lut_adj_209_LC_18_12_4 (
            .in0(N__62480),
            .in1(N__63993),
            .in2(_gnd_net_),
            .in3(N__63379),
            .lcout(n12966),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i72_4_lut_LC_18_12_5.C_ON=1'b0;
    defparam i72_4_lut_LC_18_12_5.SEQ_MODE=4'b0000;
    defparam i72_4_lut_LC_18_12_5.LUT_INIT=16'b1110010001000100;
    LogicCell40 i72_4_lut_LC_18_12_5 (
            .in0(N__62595),
            .in1(N__58378),
            .in2(N__54417),
            .in3(N__54430),
            .lcout(),
            .ltout(n37_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_301_LC_18_12_6.C_ON=1'b0;
    defparam i1_4_lut_adj_301_LC_18_12_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_301_LC_18_12_6.LUT_INIT=16'b1000100011001000;
    LogicCell40 i1_4_lut_adj_301_LC_18_12_6 (
            .in0(N__54159),
            .in1(N__54067),
            .in2(N__52009),
            .in3(N__62969),
            .lcout(n12761),
            .ltout(n12761_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12766_2_lut_LC_18_12_7.C_ON=1'b0;
    defparam i12766_2_lut_LC_18_12_7.SEQ_MODE=4'b0000;
    defparam i12766_2_lut_LC_18_12_7.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12766_2_lut_LC_18_12_7 (
            .in0(N__63380),
            .in1(_gnd_net_),
            .in2(N__52006),
            .in3(_gnd_net_),
            .lcout(n15489),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_5_i26_3_lut_LC_18_13_0.C_ON=1'b0;
    defparam mux_126_Mux_5_i26_3_lut_LC_18_13_0.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_5_i26_3_lut_LC_18_13_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_126_Mux_5_i26_3_lut_LC_18_13_0 (
            .in0(N__59505),
            .in1(N__52003),
            .in2(_gnd_net_),
            .in3(N__51981),
            .lcout(),
            .ltout(n26_adj_1730_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20414_LC_18_13_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20414_LC_18_13_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20414_LC_18_13_1.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20414_LC_18_13_1 (
            .in0(N__59554),
            .in1(N__59982),
            .in2(N__51958),
            .in3(N__60521),
            .lcout(),
            .ltout(n23336_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23336_bdd_4_lut_LC_18_13_2.C_ON=1'b0;
    defparam n23336_bdd_4_lut_LC_18_13_2.SEQ_MODE=4'b0000;
    defparam n23336_bdd_4_lut_LC_18_13_2.LUT_INIT=16'b1110010111100000;
    LogicCell40 n23336_bdd_4_lut_LC_18_13_2 (
            .in0(N__59984),
            .in1(N__51955),
            .in2(N__51928),
            .in3(N__51924),
            .lcout(),
            .ltout(n23339_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1668296_i1_3_lut_LC_18_13_3.C_ON=1'b0;
    defparam i1668296_i1_3_lut_LC_18_13_3.SEQ_MODE=4'b0000;
    defparam i1668296_i1_3_lut_LC_18_13_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1668296_i1_3_lut_LC_18_13_3 (
            .in0(_gnd_net_),
            .in1(N__52282),
            .in2(N__51901),
            .in3(N__60957),
            .lcout(),
            .ltout(n30_adj_1731_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_5_i127_3_lut_LC_18_13_4.C_ON=1'b0;
    defparam mux_126_Mux_5_i127_3_lut_LC_18_13_4.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_5_i127_3_lut_LC_18_13_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 mux_126_Mux_5_i127_3_lut_LC_18_13_4 (
            .in0(_gnd_net_),
            .in1(N__61408),
            .in2(N__51898),
            .in3(N__51895),
            .lcout(),
            .ltout(comm_buf_1_7_N_559_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i5_LC_18_13_5.C_ON=1'b0;
    defparam comm_buf_1__i5_LC_18_13_5.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i5_LC_18_13_5.LUT_INIT=16'b1011100010111000;
    LogicCell40 comm_buf_1__i5_LC_18_13_5 (
            .in0(N__55170),
            .in1(N__62600),
            .in2(N__52363),
            .in3(_gnd_net_),
            .lcout(comm_buf_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61941),
            .ce(N__55751),
            .sr(N__55714));
    defparam n23354_bdd_4_lut_LC_18_13_6.C_ON=1'b0;
    defparam n23354_bdd_4_lut_LC_18_13_6.SEQ_MODE=4'b0000;
    defparam n23354_bdd_4_lut_LC_18_13_6.LUT_INIT=16'b1111101001000100;
    LogicCell40 n23354_bdd_4_lut_LC_18_13_6 (
            .in0(N__59983),
            .in1(N__52360),
            .in2(N__52342),
            .in3(N__52297),
            .lcout(n23357),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_1_i26_3_lut_LC_18_14_0.C_ON=1'b0;
    defparam mux_126_Mux_1_i26_3_lut_LC_18_14_0.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_1_i26_3_lut_LC_18_14_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_126_Mux_1_i26_3_lut_LC_18_14_0 (
            .in0(N__52276),
            .in1(N__59503),
            .in2(_gnd_net_),
            .in3(N__52247),
            .lcout(n26_adj_1753),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19215_3_lut_LC_18_14_1.C_ON=1'b0;
    defparam i19215_3_lut_LC_18_14_1.SEQ_MODE=4'b0000;
    defparam i19215_3_lut_LC_18_14_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 i19215_3_lut_LC_18_14_1 (
            .in0(N__60519),
            .in1(N__52234),
            .in2(_gnd_net_),
            .in3(N__52207),
            .lcout(),
            .ltout(n22142_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_20468_LC_18_14_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_20468_LC_18_14_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_20468_LC_18_14_2.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_2__bdd_4_lut_20468_LC_18_14_2 (
            .in0(N__60977),
            .in1(N__59987),
            .in2(N__52183),
            .in3(N__52015),
            .lcout(),
            .ltout(n23408_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23408_bdd_4_lut_LC_18_14_3.C_ON=1'b0;
    defparam n23408_bdd_4_lut_LC_18_14_3.SEQ_MODE=4'b0000;
    defparam n23408_bdd_4_lut_LC_18_14_3.LUT_INIT=16'b1111000010101100;
    LogicCell40 n23408_bdd_4_lut_LC_18_14_3 (
            .in0(N__52180),
            .in1(N__52681),
            .in2(N__52162),
            .in3(N__60978),
            .lcout(),
            .ltout(n23411_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_1_i127_3_lut_LC_18_14_4.C_ON=1'b0;
    defparam mux_126_Mux_1_i127_3_lut_LC_18_14_4.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_1_i127_3_lut_LC_18_14_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 mux_126_Mux_1_i127_3_lut_LC_18_14_4 (
            .in0(_gnd_net_),
            .in1(N__61407),
            .in2(N__52159),
            .in3(N__52156),
            .lcout(),
            .ltout(comm_buf_1_7_N_559_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i1_LC_18_14_5.C_ON=1'b0;
    defparam comm_buf_1__i1_LC_18_14_5.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i1_LC_18_14_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i1_LC_18_14_5 (
            .in0(N__54796),
            .in1(_gnd_net_),
            .in2(N__52147),
            .in3(N__62671),
            .lcout(comm_buf_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61957),
            .ce(N__55767),
            .sr(N__55709));
    defparam i19216_4_lut_LC_18_14_6.C_ON=1'b0;
    defparam i19216_4_lut_LC_18_14_6.SEQ_MODE=4'b0000;
    defparam i19216_4_lut_LC_18_14_6.LUT_INIT=16'b1111110010111000;
    LogicCell40 i19216_4_lut_LC_18_14_6 (
            .in0(N__52039),
            .in1(N__60518),
            .in2(N__52024),
            .in3(N__59504),
            .lcout(n22143),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_4_i26_3_lut_LC_18_15_0.C_ON=1'b0;
    defparam mux_126_Mux_4_i26_3_lut_LC_18_15_0.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_4_i26_3_lut_LC_18_15_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_126_Mux_4_i26_3_lut_LC_18_15_0 (
            .in0(N__52567),
            .in1(N__59506),
            .in2(_gnd_net_),
            .in3(N__52541),
            .lcout(),
            .ltout(n26_adj_1735_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20400_LC_18_15_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20400_LC_18_15_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20400_LC_18_15_1.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_20400_LC_18_15_1 (
            .in0(N__52525),
            .in1(N__59985),
            .in2(N__52516),
            .in3(N__60520),
            .lcout(),
            .ltout(n23318_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23318_bdd_4_lut_LC_18_15_2.C_ON=1'b0;
    defparam n23318_bdd_4_lut_LC_18_15_2.SEQ_MODE=4'b0000;
    defparam n23318_bdd_4_lut_LC_18_15_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n23318_bdd_4_lut_LC_18_15_2 (
            .in0(N__59986),
            .in1(N__52512),
            .in2(N__52489),
            .in3(N__52486),
            .lcout(),
            .ltout(n23321_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1667693_i1_3_lut_LC_18_15_3.C_ON=1'b0;
    defparam i1667693_i1_3_lut_LC_18_15_3.SEQ_MODE=4'b0000;
    defparam i1667693_i1_3_lut_LC_18_15_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1667693_i1_3_lut_LC_18_15_3 (
            .in0(_gnd_net_),
            .in1(N__52462),
            .in2(N__52447),
            .in3(N__60979),
            .lcout(),
            .ltout(n30_adj_1736_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_4_i127_3_lut_LC_18_15_4.C_ON=1'b0;
    defparam mux_126_Mux_4_i127_3_lut_LC_18_15_4.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_4_i127_3_lut_LC_18_15_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_126_Mux_4_i127_3_lut_LC_18_15_4 (
            .in0(_gnd_net_),
            .in1(N__52444),
            .in2(N__52426),
            .in3(N__61352),
            .lcout(),
            .ltout(comm_buf_1_7_N_559_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i4_LC_18_15_5.C_ON=1'b0;
    defparam comm_buf_1__i4_LC_18_15_5.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i4_LC_18_15_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i4_LC_18_15_5 (
            .in0(N__55060),
            .in1(_gnd_net_),
            .in2(N__52423),
            .in3(N__62670),
            .lcout(comm_buf_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61974),
            .ce(N__55768),
            .sr(N__55700));
    defparam mux_126_Mux_2_i26_3_lut_LC_18_16_0.C_ON=1'b0;
    defparam mux_126_Mux_2_i26_3_lut_LC_18_16_0.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_2_i26_3_lut_LC_18_16_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_126_Mux_2_i26_3_lut_LC_18_16_0 (
            .in0(N__52419),
            .in1(N__59507),
            .in2(_gnd_net_),
            .in3(N__52397),
            .lcout(),
            .ltout(n26_adj_1748_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19225_4_lut_LC_18_16_1.C_ON=1'b0;
    defparam i19225_4_lut_LC_18_16_1.SEQ_MODE=4'b0000;
    defparam i19225_4_lut_LC_18_16_1.LUT_INIT=16'b0100010011110000;
    LogicCell40 i19225_4_lut_LC_18_16_1 (
            .in0(N__59508),
            .in1(N__52378),
            .in2(N__52366),
            .in3(N__60647),
            .lcout(),
            .ltout(n22152_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_20493_LC_18_16_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_20493_LC_18_16_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_20493_LC_18_16_2.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_2__bdd_4_lut_20493_LC_18_16_2 (
            .in0(N__52786),
            .in1(N__60065),
            .in2(N__52993),
            .in3(N__61024),
            .lcout(),
            .ltout(n23444_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23444_bdd_4_lut_LC_18_16_3.C_ON=1'b0;
    defparam n23444_bdd_4_lut_LC_18_16_3.SEQ_MODE=4'b0000;
    defparam n23444_bdd_4_lut_LC_18_16_3.LUT_INIT=16'b1110010111100000;
    LogicCell40 n23444_bdd_4_lut_LC_18_16_3 (
            .in0(N__61025),
            .in1(N__52990),
            .in2(N__52972),
            .in3(N__52969),
            .lcout(),
            .ltout(n23447_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_2_i127_3_lut_LC_18_16_4.C_ON=1'b0;
    defparam mux_126_Mux_2_i127_3_lut_LC_18_16_4.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_2_i127_3_lut_LC_18_16_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_126_Mux_2_i127_3_lut_LC_18_16_4 (
            .in0(_gnd_net_),
            .in1(N__52957),
            .in2(N__52942),
            .in3(N__61411),
            .lcout(),
            .ltout(comm_buf_1_7_N_559_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i2_LC_18_16_5.C_ON=1'b0;
    defparam comm_buf_1__i2_LC_18_16_5.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i2_LC_18_16_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i2_LC_18_16_5 (
            .in0(_gnd_net_),
            .in1(N__54929),
            .in2(N__52939),
            .in3(N__62672),
            .lcout(comm_buf_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61986),
            .ce(N__55774),
            .sr(N__55708));
    defparam i19224_3_lut_LC_18_16_6.C_ON=1'b0;
    defparam i19224_3_lut_LC_18_16_6.SEQ_MODE=4'b0000;
    defparam i19224_3_lut_LC_18_16_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i19224_3_lut_LC_18_16_6 (
            .in0(N__60646),
            .in1(N__52843),
            .in2(_gnd_net_),
            .in3(N__52812),
            .lcout(n22151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i23_3_lut_LC_18_17_2.C_ON=1'b0;
    defparam mux_125_Mux_3_i23_3_lut_LC_18_17_2.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i23_3_lut_LC_18_17_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_125_Mux_3_i23_3_lut_LC_18_17_2 (
            .in0(N__52779),
            .in1(N__59410),
            .in2(_gnd_net_),
            .in3(N__52744),
            .lcout(n23_adj_1791),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19209_3_lut_LC_18_17_7.C_ON=1'b0;
    defparam i19209_3_lut_LC_18_17_7.SEQ_MODE=4'b0000;
    defparam i19209_3_lut_LC_18_17_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i19209_3_lut_LC_18_17_7 (
            .in0(N__52716),
            .in1(N__52690),
            .in2(_gnd_net_),
            .in3(N__60593),
            .lcout(n22136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16252_2_lut_2_lut_LC_18_18_5.C_ON=1'b0;
    defparam i16252_2_lut_2_lut_LC_18_18_5.SEQ_MODE=4'b0000;
    defparam i16252_2_lut_2_lut_LC_18_18_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i16252_2_lut_2_lut_LC_18_18_5 (
            .in0(_gnd_net_),
            .in1(N__52669),
            .in2(_gnd_net_),
            .in3(N__52638),
            .lcout(CONT_SD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_0_i15_4_lut_LC_18_19_6.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_0_i15_4_lut_LC_18_19_6.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_0_i15_4_lut_LC_18_19_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_358_Mux_0_i15_4_lut_LC_18_19_6 (
            .in0(N__63525),
            .in1(N__52588),
            .in2(N__57872),
            .in3(N__53151),
            .lcout(data_index_9_N_236_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20091_2_lut_LC_19_4_7.C_ON=1'b0;
    defparam i20091_2_lut_LC_19_4_7.SEQ_MODE=4'b0000;
    defparam i20091_2_lut_LC_19_4_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i20091_2_lut_LC_19_4_7 (
            .in0(_gnd_net_),
            .in1(N__53035),
            .in2(_gnd_net_),
            .in3(N__59399),
            .lcout(n22500),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0on_i0_LC_19_5_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i0_LC_19_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i0_LC_19_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i0_LC_19_5_0  (
            .in0(_gnd_net_),
            .in1(N__56722),
            .in2(_gnd_net_),
            .in3(N__53014),
            .lcout(\ADC_VDC.genclk.t0on_0 ),
            .ltout(),
            .carryin(bfn_19_5_0_),
            .carryout(\ADC_VDC.genclk.n20751 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i1_LC_19_5_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i1_LC_19_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i1_LC_19_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i1_LC_19_5_1  (
            .in0(_gnd_net_),
            .in1(N__56752),
            .in2(N__64844),
            .in3(N__53011),
            .lcout(\ADC_VDC.genclk.t0on_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20751 ),
            .carryout(\ADC_VDC.genclk.n20752 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i2_LC_19_5_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i2_LC_19_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i2_LC_19_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i2_LC_19_5_2  (
            .in0(_gnd_net_),
            .in1(N__64780),
            .in2(N__56692),
            .in3(N__53008),
            .lcout(\ADC_VDC.genclk.t0on_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20752 ),
            .carryout(\ADC_VDC.genclk.n20753 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i3_LC_19_5_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i3_LC_19_5_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0on_i3_LC_19_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i3_LC_19_5_3  (
            .in0(_gnd_net_),
            .in1(N__57244),
            .in2(N__64845),
            .in3(N__53005),
            .lcout(\ADC_VDC.genclk.t0on_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20753 ),
            .carryout(\ADC_VDC.genclk.n20754 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i4_LC_19_5_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i4_LC_19_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i4_LC_19_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i4_LC_19_5_4  (
            .in0(_gnd_net_),
            .in1(N__64784),
            .in2(N__56740),
            .in3(N__53002),
            .lcout(\ADC_VDC.genclk.t0on_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20754 ),
            .carryout(\ADC_VDC.genclk.n20755 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i5_LC_19_5_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i5_LC_19_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i5_LC_19_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i5_LC_19_5_5  (
            .in0(_gnd_net_),
            .in1(N__57231),
            .in2(N__64846),
            .in3(N__52999),
            .lcout(\ADC_VDC.genclk.t0on_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20755 ),
            .carryout(\ADC_VDC.genclk.n20756 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i6_LC_19_5_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i6_LC_19_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i6_LC_19_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i6_LC_19_5_6  (
            .in0(_gnd_net_),
            .in1(N__64788),
            .in2(N__56767),
            .in3(N__52996),
            .lcout(\ADC_VDC.genclk.t0on_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20756 ),
            .carryout(\ADC_VDC.genclk.n20757 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i7_LC_19_5_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i7_LC_19_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i7_LC_19_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i7_LC_19_5_7  (
            .in0(_gnd_net_),
            .in1(N__56676),
            .in2(N__64847),
            .in3(N__53179),
            .lcout(\ADC_VDC.genclk.t0on_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20757 ),
            .carryout(\ADC_VDC.genclk.n20758 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57199),
            .sr(N__64447));
    defparam \ADC_VDC.genclk.t0on_i8_LC_19_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i8_LC_19_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i8_LC_19_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i8_LC_19_6_0  (
            .in0(_gnd_net_),
            .in1(N__57217),
            .in2(N__64696),
            .in3(N__53176),
            .lcout(\ADC_VDC.genclk.t0on_8 ),
            .ltout(),
            .carryin(bfn_19_6_0_),
            .carryout(\ADC_VDC.genclk.n20759 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam \ADC_VDC.genclk.t0on_i9_LC_19_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i9_LC_19_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i9_LC_19_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i9_LC_19_6_1  (
            .in0(_gnd_net_),
            .in1(N__64641),
            .in2(N__56632),
            .in3(N__53173),
            .lcout(\ADC_VDC.genclk.t0on_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20759 ),
            .carryout(\ADC_VDC.genclk.n20760 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam \ADC_VDC.genclk.t0on_i10_LC_19_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i10_LC_19_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i10_LC_19_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i10_LC_19_6_2  (
            .in0(_gnd_net_),
            .in1(N__56662),
            .in2(N__64693),
            .in3(N__53170),
            .lcout(\ADC_VDC.genclk.t0on_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20760 ),
            .carryout(\ADC_VDC.genclk.n20761 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam \ADC_VDC.genclk.t0on_i11_LC_19_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i11_LC_19_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i11_LC_19_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i11_LC_19_6_3  (
            .in0(_gnd_net_),
            .in1(N__64629),
            .in2(N__56602),
            .in3(N__53167),
            .lcout(\ADC_VDC.genclk.t0on_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20761 ),
            .carryout(\ADC_VDC.genclk.n20762 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam \ADC_VDC.genclk.t0on_i12_LC_19_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i12_LC_19_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i12_LC_19_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i12_LC_19_6_4  (
            .in0(_gnd_net_),
            .in1(N__56706),
            .in2(N__64694),
            .in3(N__53164),
            .lcout(\ADC_VDC.genclk.t0on_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20762 ),
            .carryout(\ADC_VDC.genclk.n20763 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam \ADC_VDC.genclk.t0on_i13_LC_19_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i13_LC_19_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i13_LC_19_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i13_LC_19_6_5  (
            .in0(_gnd_net_),
            .in1(N__64633),
            .in2(N__57262),
            .in3(N__53161),
            .lcout(\ADC_VDC.genclk.t0on_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20763 ),
            .carryout(\ADC_VDC.genclk.n20764 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam \ADC_VDC.genclk.t0on_i14_LC_19_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i14_LC_19_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i14_LC_19_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i14_LC_19_6_6  (
            .in0(_gnd_net_),
            .in1(N__56644),
            .in2(N__64695),
            .in3(N__53158),
            .lcout(\ADC_VDC.genclk.t0on_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20764 ),
            .carryout(\ADC_VDC.genclk.n20765 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam \ADC_VDC.genclk.t0on_i15_LC_19_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0on_i15_LC_19_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i15_LC_19_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0on_i15_LC_19_6_7  (
            .in0(N__56616),
            .in1(N__64637),
            .in2(_gnd_net_),
            .in3(N__53155),
            .lcout(\ADC_VDC.genclk.t0on_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57195),
            .sr(N__64457));
    defparam dds0_mclkcnt_i7_3792__i0_LC_19_7_0.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3792__i0_LC_19_7_0.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i0_LC_19_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i0_LC_19_7_0 (
            .in0(_gnd_net_),
            .in1(N__53245),
            .in2(_gnd_net_),
            .in3(N__53209),
            .lcout(dds0_mclkcnt_0),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(n20819),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3792__i1_LC_19_7_1.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3792__i1_LC_19_7_1.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i1_LC_19_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i1_LC_19_7_1 (
            .in0(_gnd_net_),
            .in1(N__53286),
            .in2(_gnd_net_),
            .in3(N__53206),
            .lcout(dds0_mclkcnt_1),
            .ltout(),
            .carryin(n20819),
            .carryout(n20820),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3792__i2_LC_19_7_2.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3792__i2_LC_19_7_2.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i2_LC_19_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i2_LC_19_7_2 (
            .in0(_gnd_net_),
            .in1(N__53230),
            .in2(_gnd_net_),
            .in3(N__53203),
            .lcout(dds0_mclkcnt_2),
            .ltout(),
            .carryin(n20820),
            .carryout(n20821),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3792__i3_LC_19_7_3.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3792__i3_LC_19_7_3.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i3_LC_19_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i3_LC_19_7_3 (
            .in0(_gnd_net_),
            .in1(N__53314),
            .in2(_gnd_net_),
            .in3(N__53200),
            .lcout(dds0_mclkcnt_3),
            .ltout(),
            .carryin(n20821),
            .carryout(n20822),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3792__i4_LC_19_7_4.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3792__i4_LC_19_7_4.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i4_LC_19_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i4_LC_19_7_4 (
            .in0(_gnd_net_),
            .in1(N__53272),
            .in2(_gnd_net_),
            .in3(N__53197),
            .lcout(dds0_mclkcnt_4),
            .ltout(),
            .carryin(n20822),
            .carryout(n20823),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3792__i5_LC_19_7_5.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3792__i5_LC_19_7_5.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i5_LC_19_7_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i5_LC_19_7_5 (
            .in0(_gnd_net_),
            .in1(N__53302),
            .in2(_gnd_net_),
            .in3(N__53194),
            .lcout(dds0_mclkcnt_5),
            .ltout(),
            .carryin(n20823),
            .carryout(n20824),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3792__i6_LC_19_7_6.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3792__i6_LC_19_7_6.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i6_LC_19_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i6_LC_19_7_6 (
            .in0(_gnd_net_),
            .in1(N__53185),
            .in2(_gnd_net_),
            .in3(N__53191),
            .lcout(dds0_mclkcnt_6),
            .ltout(),
            .carryin(n20824),
            .carryout(n20825),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3792__i7_LC_19_7_7.C_ON=1'b0;
    defparam dds0_mclkcnt_i7_3792__i7_LC_19_7_7.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3792__i7_LC_19_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3792__i7_LC_19_7_7 (
            .in0(_gnd_net_),
            .in1(N__53259),
            .in2(_gnd_net_),
            .in3(N__53188),
            .lcout(dds0_mclkcnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclkcnt_i7_3792__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i16388_2_lut_LC_19_8_0.C_ON=1'b0;
    defparam i16388_2_lut_LC_19_8_0.SEQ_MODE=4'b0000;
    defparam i16388_2_lut_LC_19_8_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 i16388_2_lut_LC_19_8_0 (
            .in0(_gnd_net_),
            .in1(N__53391),
            .in2(_gnd_net_),
            .in3(N__53217),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclk_297_LC_19_8_1.C_ON=1'b0;
    defparam dds0_mclk_297_LC_19_8_1.SEQ_MODE=4'b1000;
    defparam dds0_mclk_297_LC_19_8_1.LUT_INIT=16'b1001100111001100;
    LogicCell40 dds0_mclk_297_LC_19_8_1 (
            .in0(N__53218),
            .in1(N__53364),
            .in2(_gnd_net_),
            .in3(N__53392),
            .lcout(DDS_MCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclk_297C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i4170_2_lut_LC_19_8_2.C_ON=1'b0;
    defparam i4170_2_lut_LC_19_8_2.SEQ_MODE=4'b0000;
    defparam i4170_2_lut_LC_19_8_2.LUT_INIT=16'b1111111110101010;
    LogicCell40 i4170_2_lut_LC_19_8_2 (
            .in0(N__58193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58030),
            .lcout(),
            .ltout(n6888_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_72_LC_19_8_3.C_ON=1'b0;
    defparam i1_4_lut_adj_72_LC_19_8_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_72_LC_19_8_3.LUT_INIT=16'b1111111000000000;
    LogicCell40 i1_4_lut_adj_72_LC_19_8_3 (
            .in0(N__53320),
            .in1(N__54175),
            .in2(N__53353),
            .in3(N__53326),
            .lcout(n21865),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_71_LC_19_8_4.C_ON=1'b0;
    defparam i1_4_lut_adj_71_LC_19_8_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_71_LC_19_8_4.LUT_INIT=16'b1111001110110011;
    LogicCell40 i1_4_lut_adj_71_LC_19_8_4 (
            .in0(N__63190),
            .in1(N__63056),
            .in2(N__53338),
            .in3(N__57905),
            .lcout(n22027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_75_LC_19_8_5.C_ON=1'b0;
    defparam i1_2_lut_adj_75_LC_19_8_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_75_LC_19_8_5.LUT_INIT=16'b1010101011111111;
    LogicCell40 i1_2_lut_adj_75_LC_19_8_5 (
            .in0(N__63055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62290),
            .lcout(n22018),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_243_LC_19_8_6.C_ON=1'b0;
    defparam i5_4_lut_adj_243_LC_19_8_6.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_243_LC_19_8_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_adj_243_LC_19_8_6 (
            .in0(N__53313),
            .in1(N__53301),
            .in2(N__53290),
            .in3(N__53271),
            .lcout(),
            .ltout(n12_adj_1685_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_248_LC_19_8_7.C_ON=1'b0;
    defparam i6_4_lut_adj_248_LC_19_8_7.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_248_LC_19_8_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_248_LC_19_8_7 (
            .in0(N__53260),
            .in1(N__53244),
            .in2(N__53233),
            .in3(N__53229),
            .lcout(n21857),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_valid_85_LC_19_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_valid_85_LC_19_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_valid_85_LC_19_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.data_valid_85_LC_19_9_0  (
            .in0(_gnd_net_),
            .in1(N__53785),
            .in2(_gnd_net_),
            .in3(N__53740),
            .lcout(comm_data_vld),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.data_valid_85C_net ),
            .ce(),
            .sr(N__57078));
    defparam \comm_spi.data_rx_i7_LC_19_10_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i7_LC_19_10_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i7_LC_19_10_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i7_LC_19_10_0  (
            .in0(N__53781),
            .in1(N__53837),
            .in2(_gnd_net_),
            .in3(N__53739),
            .lcout(comm_rx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53677),
            .ce(),
            .sr(N__57092));
    defparam \comm_spi.data_rx_i6_LC_19_10_1 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i6_LC_19_10_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i6_LC_19_10_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i6_LC_19_10_1  (
            .in0(N__53738),
            .in1(N__55132),
            .in2(_gnd_net_),
            .in3(N__53780),
            .lcout(comm_rx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53677),
            .ce(),
            .sr(N__57092));
    defparam \comm_spi.data_rx_i5_LC_19_10_2 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i5_LC_19_10_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i5_LC_19_10_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i5_LC_19_10_2  (
            .in0(N__53779),
            .in1(N__55016),
            .in2(_gnd_net_),
            .in3(N__53737),
            .lcout(comm_rx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53677),
            .ce(),
            .sr(N__57092));
    defparam \comm_spi.data_rx_i4_LC_19_10_3 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i4_LC_19_10_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i4_LC_19_10_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i4_LC_19_10_3  (
            .in0(N__53736),
            .in1(N__62727),
            .in2(_gnd_net_),
            .in3(N__53778),
            .lcout(comm_rx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53677),
            .ce(),
            .sr(N__57092));
    defparam \comm_spi.data_rx_i3_LC_19_10_4 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i3_LC_19_10_4 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i3_LC_19_10_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i3_LC_19_10_4  (
            .in0(N__53777),
            .in1(N__54878),
            .in2(_gnd_net_),
            .in3(N__53735),
            .lcout(comm_rx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53677),
            .ce(),
            .sr(N__57092));
    defparam \comm_spi.data_rx_i2_LC_19_10_5 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i2_LC_19_10_5 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i2_LC_19_10_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i2_LC_19_10_5  (
            .in0(N__53734),
            .in1(N__54750),
            .in2(_gnd_net_),
            .in3(N__53776),
            .lcout(comm_rx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53677),
            .ce(),
            .sr(N__57092));
    defparam \comm_spi.data_rx_i1_LC_19_10_6 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i1_LC_19_10_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i1_LC_19_10_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \comm_spi.data_rx_i1_LC_19_10_6  (
            .in0(N__53775),
            .in1(N__53733),
            .in2(_gnd_net_),
            .in3(N__54022),
            .lcout(comm_rx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53677),
            .ce(),
            .sr(N__57092));
    defparam i19760_4_lut_LC_19_11_0.C_ON=1'b0;
    defparam i19760_4_lut_LC_19_11_0.SEQ_MODE=4'b0000;
    defparam i19760_4_lut_LC_19_11_0.LUT_INIT=16'b1110111011111010;
    LogicCell40 i19760_4_lut_LC_19_11_0 (
            .in0(N__63084),
            .in1(N__53464),
            .in2(N__53455),
            .in3(N__61405),
            .lcout(),
            .ltout(n22321_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_1__bdd_4_lut_LC_19_11_1.C_ON=1'b0;
    defparam comm_state_1__bdd_4_lut_LC_19_11_1.SEQ_MODE=4'b0000;
    defparam comm_state_1__bdd_4_lut_LC_19_11_1.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_state_1__bdd_4_lut_LC_19_11_1 (
            .in0(N__62369),
            .in1(N__53446),
            .in2(N__53419),
            .in3(N__63889),
            .lcout(n23342),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20000_4_lut_LC_19_11_2.C_ON=1'b0;
    defparam i20000_4_lut_LC_19_11_2.SEQ_MODE=4'b0000;
    defparam i20000_4_lut_LC_19_11_2.LUT_INIT=16'b0101010000000100;
    LogicCell40 i20000_4_lut_LC_19_11_2 (
            .in0(N__53409),
            .in1(N__58411),
            .in2(N__61414),
            .in3(N__55558),
            .lcout(n22352),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_299_LC_19_11_3.C_ON=1'b0;
    defparam i1_2_lut_adj_299_LC_19_11_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_299_LC_19_11_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_299_LC_19_11_3 (
            .in0(_gnd_net_),
            .in1(N__54585),
            .in2(_gnd_net_),
            .in3(N__54444),
            .lcout(n21862),
            .ltout(n21862_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i44_4_lut_LC_19_11_4.C_ON=1'b0;
    defparam i44_4_lut_LC_19_11_4.SEQ_MODE=4'b0000;
    defparam i44_4_lut_LC_19_11_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 i44_4_lut_LC_19_11_4 (
            .in0(N__54419),
            .in1(N__62368),
            .in2(N__54205),
            .in3(N__54202),
            .lcout(),
            .ltout(n22_adj_1725_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_294_LC_19_11_5.C_ON=1'b0;
    defparam i1_4_lut_adj_294_LC_19_11_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_294_LC_19_11_5.LUT_INIT=16'b1011101000000000;
    LogicCell40 i1_4_lut_adj_294_LC_19_11_5 (
            .in0(N__54182),
            .in1(N__63083),
            .in2(N__54091),
            .in3(N__54065),
            .lcout(n12677),
            .ltout(n12677_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12759_2_lut_LC_19_11_6.C_ON=1'b0;
    defparam i12759_2_lut_LC_19_11_6.SEQ_MODE=4'b0000;
    defparam i12759_2_lut_LC_19_11_6.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12759_2_lut_LC_19_11_6 (
            .in0(N__63528),
            .in1(_gnd_net_),
            .in2(N__54088),
            .in3(_gnd_net_),
            .lcout(n15482),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_19_11_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_19_11_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_19_11_7.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_LC_19_11_7 (
            .in0(N__63110),
            .in1(N__63888),
            .in2(_gnd_net_),
            .in3(N__63527),
            .lcout(n21895),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i0_LC_19_12_0.C_ON=1'b0;
    defparam comm_buf_4__i0_LC_19_12_0.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i0_LC_19_12_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_4__i0_LC_19_12_0 (
            .in0(N__54037),
            .in1(N__62525),
            .in2(_gnd_net_),
            .in3(N__54021),
            .lcout(comm_buf_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam comm_buf_4__i7_LC_19_12_1.C_ON=1'b0;
    defparam comm_buf_4__i7_LC_19_12_1.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i7_LC_19_12_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i7_LC_19_12_1 (
            .in0(N__62524),
            .in1(N__55884),
            .in2(_gnd_net_),
            .in3(N__53920),
            .lcout(comm_buf_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam comm_buf_4__i6_LC_19_12_2.C_ON=1'b0;
    defparam comm_buf_4__i6_LC_19_12_2.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i6_LC_19_12_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i6_LC_19_12_2 (
            .in0(N__53855),
            .in1(N__53812),
            .in2(_gnd_net_),
            .in3(N__62528),
            .lcout(comm_buf_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam comm_buf_4__i5_LC_19_12_3.C_ON=1'b0;
    defparam comm_buf_4__i5_LC_19_12_3.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i5_LC_19_12_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_4__i5_LC_19_12_3 (
            .in0(N__62523),
            .in1(_gnd_net_),
            .in2(N__55169),
            .in3(N__55105),
            .lcout(comm_buf_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam comm_buf_4__i4_LC_19_12_4.C_ON=1'b0;
    defparam comm_buf_4__i4_LC_19_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i4_LC_19_12_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i4_LC_19_12_4 (
            .in0(N__55038),
            .in1(N__54991),
            .in2(_gnd_net_),
            .in3(N__62527),
            .lcout(comm_buf_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam comm_buf_4__i3_LC_19_12_5.C_ON=1'b0;
    defparam comm_buf_4__i3_LC_19_12_5.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i3_LC_19_12_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_4__i3_LC_19_12_5 (
            .in0(N__62522),
            .in1(_gnd_net_),
            .in2(N__62775),
            .in3(N__54964),
            .lcout(comm_buf_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam comm_buf_4__i2_LC_19_12_6.C_ON=1'b0;
    defparam comm_buf_4__i2_LC_19_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i2_LC_19_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i2_LC_19_12_6 (
            .in0(N__54896),
            .in1(N__54850),
            .in2(_gnd_net_),
            .in3(N__62526),
            .lcout(comm_buf_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam comm_buf_4__i1_LC_19_12_7.C_ON=1'b0;
    defparam comm_buf_4__i1_LC_19_12_7.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i1_LC_19_12_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i1_LC_19_12_7 (
            .in0(N__62521),
            .in1(N__54769),
            .in2(_gnd_net_),
            .in3(N__54724),
            .lcout(comm_buf_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61942),
            .ce(N__54694),
            .sr(N__54688));
    defparam mux_126_Mux_7_i26_3_lut_LC_19_13_0.C_ON=1'b0;
    defparam mux_126_Mux_7_i26_3_lut_LC_19_13_0.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_7_i26_3_lut_LC_19_13_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_126_Mux_7_i26_3_lut_LC_19_13_0 (
            .in0(N__54676),
            .in1(N__59425),
            .in2(_gnd_net_),
            .in3(N__54657),
            .lcout(),
            .ltout(n26_adj_1716_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19336_4_lut_LC_19_13_1.C_ON=1'b0;
    defparam i19336_4_lut_LC_19_13_1.SEQ_MODE=4'b0000;
    defparam i19336_4_lut_LC_19_13_1.LUT_INIT=16'b1110111011110000;
    LogicCell40 i19336_4_lut_LC_19_13_1 (
            .in0(N__59426),
            .in1(N__54628),
            .in2(N__54619),
            .in3(N__60522),
            .lcout(),
            .ltout(n22263_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_20488_LC_19_13_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_20488_LC_19_13_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_20488_LC_19_13_2.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_2__bdd_4_lut_20488_LC_19_13_2 (
            .in0(N__59904),
            .in1(N__55456),
            .in2(N__54616),
            .in3(N__60955),
            .lcout(),
            .ltout(n23420_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23420_bdd_4_lut_LC_19_13_3.C_ON=1'b0;
    defparam n23420_bdd_4_lut_LC_19_13_3.SEQ_MODE=4'b0000;
    defparam n23420_bdd_4_lut_LC_19_13_3.LUT_INIT=16'b1110010111100000;
    LogicCell40 n23420_bdd_4_lut_LC_19_13_3 (
            .in0(N__60956),
            .in1(N__55999),
            .in2(N__55981),
            .in3(N__55978),
            .lcout(),
            .ltout(n23423_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_126_Mux_7_i127_3_lut_LC_19_13_4.C_ON=1'b0;
    defparam mux_126_Mux_7_i127_3_lut_LC_19_13_4.SEQ_MODE=4'b0000;
    defparam mux_126_Mux_7_i127_3_lut_LC_19_13_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_126_Mux_7_i127_3_lut_LC_19_13_4 (
            .in0(_gnd_net_),
            .in1(N__55966),
            .in2(N__55948),
            .in3(N__61409),
            .lcout(),
            .ltout(comm_buf_1_7_N_559_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i7_LC_19_13_5.C_ON=1'b0;
    defparam comm_buf_1__i7_LC_19_13_5.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i7_LC_19_13_5.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_1__i7_LC_19_13_5 (
            .in0(N__62529),
            .in1(N__55899),
            .in2(N__55852),
            .in3(_gnd_net_),
            .lcout(comm_buf_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61958),
            .ce(N__55770),
            .sr(N__55710));
    defparam i19746_3_lut_LC_19_14_0.C_ON=1'b0;
    defparam i19746_3_lut_LC_19_14_0.SEQ_MODE=4'b0000;
    defparam i19746_3_lut_LC_19_14_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 i19746_3_lut_LC_19_14_0 (
            .in0(N__55630),
            .in1(N__56185),
            .in2(_gnd_net_),
            .in3(N__58522),
            .lcout(n22356),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23348_bdd_4_lut_LC_19_14_1.C_ON=1'b0;
    defparam n23348_bdd_4_lut_LC_19_14_1.SEQ_MODE=4'b0000;
    defparam n23348_bdd_4_lut_LC_19_14_1.LUT_INIT=16'b1110111001010000;
    LogicCell40 n23348_bdd_4_lut_LC_19_14_1 (
            .in0(N__60516),
            .in1(N__55223),
            .in2(N__55548),
            .in3(N__55510),
            .lcout(n23351),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19335_3_lut_LC_19_14_3.C_ON=1'b0;
    defparam i19335_3_lut_LC_19_14_3.SEQ_MODE=4'b0000;
    defparam i19335_3_lut_LC_19_14_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i19335_3_lut_LC_19_14_3 (
            .in0(N__60517),
            .in1(N__55501),
            .in2(_gnd_net_),
            .in3(N__55477),
            .lcout(n22262),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20112_2_lut_LC_19_14_6.C_ON=1'b0;
    defparam i20112_2_lut_LC_19_14_6.SEQ_MODE=4'b0000;
    defparam i20112_2_lut_LC_19_14_6.LUT_INIT=16'b0000101000001010;
    LogicCell40 i20112_2_lut_LC_19_14_6 (
            .in0(N__55450),
            .in1(_gnd_net_),
            .in2(N__59517),
            .in3(_gnd_net_),
            .lcout(n22391),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i13_LC_19_14_7.C_ON=1'b0;
    defparam buf_dds1_i13_LC_19_14_7.SEQ_MODE=4'b1000;
    defparam buf_dds1_i13_LC_19_14_7.LUT_INIT=16'b1110111000101110;
    LogicCell40 buf_dds1_i13_LC_19_14_7 (
            .in0(N__55227),
            .in1(N__55380),
            .in2(N__63737),
            .in3(N__55288),
            .lcout(buf_dds1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61975),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i5_LC_19_15_0.C_ON=1'b0;
    defparam data_index_i5_LC_19_15_0.SEQ_MODE=4'b1000;
    defparam data_index_i5_LC_19_15_0.LUT_INIT=16'b0101000011011000;
    LogicCell40 data_index_i5_LC_19_15_0 (
            .in0(N__63643),
            .in1(N__56389),
            .in2(N__56380),
            .in3(N__57730),
            .lcout(data_index_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61987),
            .ce(),
            .sr(_gnd_net_));
    defparam i16198_3_lut_LC_19_15_1.C_ON=1'b0;
    defparam i16198_3_lut_LC_19_15_1.SEQ_MODE=4'b0000;
    defparam i16198_3_lut_LC_19_15_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i16198_3_lut_LC_19_15_1 (
            .in0(N__56532),
            .in1(N__56495),
            .in2(_gnd_net_),
            .in3(N__56478),
            .lcout(n8_adj_1623),
            .ltout(n8_adj_1623_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_358_Mux_5_i15_4_lut_LC_19_15_2.C_ON=1'b0;
    defparam comm_state_3__I_0_358_Mux_5_i15_4_lut_LC_19_15_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_358_Mux_5_i15_4_lut_LC_19_15_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_state_3__I_0_358_Mux_5_i15_4_lut_LC_19_15_2 (
            .in0(N__63642),
            .in1(N__57728),
            .in2(N__56383),
            .in3(N__56376),
            .lcout(data_index_9_N_236_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds1_308_LC_19_15_3.C_ON=1'b0;
    defparam trig_dds1_308_LC_19_15_3.SEQ_MODE=4'b1000;
    defparam trig_dds1_308_LC_19_15_3.LUT_INIT=16'b0110000001100100;
    LogicCell40 trig_dds1_308_LC_19_15_3 (
            .in0(N__57729),
            .in1(N__63644),
            .in2(N__56205),
            .in3(N__56257),
            .lcout(trig_dds1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61987),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_298_LC_19_15_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_298_LC_19_15_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_298_LC_19_15_4.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_adj_298_LC_19_15_4 (
            .in0(N__60953),
            .in1(N__59900),
            .in2(_gnd_net_),
            .in3(N__58641),
            .lcout(n21920),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19888_4_lut_LC_19_15_5.C_ON=1'b0;
    defparam i19888_4_lut_LC_19_15_5.SEQ_MODE=4'b0000;
    defparam i19888_4_lut_LC_19_15_5.LUT_INIT=16'b0000000101000000;
    LogicCell40 i19888_4_lut_LC_19_15_5 (
            .in0(N__58642),
            .in1(N__60954),
            .in2(N__60014),
            .in3(N__59400),
            .lcout(),
            .ltout(n22399_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i59_4_lut_LC_19_15_6.C_ON=1'b0;
    defparam i59_4_lut_LC_19_15_6.SEQ_MODE=4'b0000;
    defparam i59_4_lut_LC_19_15_6.LUT_INIT=16'b1000100011110000;
    LogicCell40 i59_4_lut_LC_19_15_6 (
            .in0(N__59401),
            .in1(N__56184),
            .in2(N__56173),
            .in3(N__61401),
            .lcout(n40_adj_1689),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i26_3_lut_LC_19_16_4.C_ON=1'b0;
    defparam mux_125_Mux_3_i26_3_lut_LC_19_16_4.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i26_3_lut_LC_19_16_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_125_Mux_3_i26_3_lut_LC_19_16_4 (
            .in0(N__59497),
            .in1(N__56158),
            .in2(_gnd_net_),
            .in3(N__56133),
            .lcout(n26_adj_1792),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16465_2_lut_3_lut_LC_19_17_2.C_ON=1'b0;
    defparam i16465_2_lut_3_lut_LC_19_17_2.SEQ_MODE=4'b0000;
    defparam i16465_2_lut_3_lut_LC_19_17_2.LUT_INIT=16'b0000000000100010;
    LogicCell40 i16465_2_lut_3_lut_LC_19_17_2 (
            .in0(N__56074),
            .in1(N__62646),
            .in2(_gnd_net_),
            .in3(N__64049),
            .lcout(n14_adj_1611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16456_2_lut_3_lut_LC_19_17_4.C_ON=1'b0;
    defparam i16456_2_lut_3_lut_LC_19_17_4.SEQ_MODE=4'b0000;
    defparam i16456_2_lut_3_lut_LC_19_17_4.LUT_INIT=16'b0000000000100010;
    LogicCell40 i16456_2_lut_3_lut_LC_19_17_4 (
            .in0(N__62056),
            .in1(N__62645),
            .in2(_gnd_net_),
            .in3(N__64048),
            .lcout(n14_adj_1654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i20146_2_lut_4_lut_LC_20_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i20146_2_lut_4_lut_LC_20_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i20146_2_lut_4_lut_LC_20_5_0 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \ADC_VDC.genclk.i20146_2_lut_4_lut_LC_20_5_0  (
            .in0(N__64219),
            .in1(N__64179),
            .in2(N__64168),
            .in3(N__64237),
            .lcout(\ADC_VDC.genclk.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i1_LC_20_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i1_LC_20_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i1_LC_20_5_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ADC_VDC.genclk.div_state_i1_LC_20_5_1  (
            .in0(_gnd_net_),
            .in1(N__64167),
            .in2(_gnd_net_),
            .in3(N__64220),
            .lcout(\ADC_VDC.genclk.div_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i1C_net ),
            .ce(N__56776),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i20156_2_lut_LC_20_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i20156_2_lut_LC_20_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i20156_2_lut_LC_20_5_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ADC_VDC.genclk.i20156_2_lut_LC_20_5_2  (
            .in0(_gnd_net_),
            .in1(N__64162),
            .in2(_gnd_net_),
            .in3(N__64216),
            .lcout(\ADC_VDC.genclk.n15418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i20142_2_lut_LC_20_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i20142_2_lut_LC_20_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i20142_2_lut_LC_20_5_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ADC_VDC.genclk.i20142_2_lut_LC_20_5_3  (
            .in0(N__64217),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64163),
            .lcout(\ADC_VDC.genclk.n12361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19910_4_lut_LC_20_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19910_4_lut_LC_20_6_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19910_4_lut_LC_20_6_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i19910_4_lut_LC_20_6_0  (
            .in0(N__56763),
            .in1(N__56751),
            .in2(N__56739),
            .in3(N__56721),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n22308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i20049_4_lut_LC_20_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i20049_4_lut_LC_20_6_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i20049_4_lut_LC_20_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i20049_4_lut_LC_20_6_1  (
            .in0(N__57268),
            .in1(N__57205),
            .in2(N__56710),
            .in3(N__56650),
            .lcout(\ADC_VDC.genclk.n22302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_adj_5_LC_20_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_5_LC_20_6_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_5_LC_20_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_adj_5_LC_20_6_2  (
            .in0(N__56707),
            .in1(N__56688),
            .in2(N__56677),
            .in3(N__56661),
            .lcout(\ADC_VDC.genclk.n27_adj_1483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_adj_3_LC_20_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_3_LC_20_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_3_LC_20_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_adj_3_LC_20_6_3  (
            .in0(N__56643),
            .in1(N__56628),
            .in2(N__56617),
            .in3(N__56598),
            .lcout(\ADC_VDC.genclk.n28_adj_1481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_adj_4_LC_20_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_4_LC_20_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_4_LC_20_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_adj_4_LC_20_6_4  (
            .in0(N__57261),
            .in1(N__57243),
            .in2(N__57232),
            .in3(N__57216),
            .lcout(\ADC_VDC.genclk.n26_adj_1482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_20_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_20_6_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_20_6_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_20_6_6  (
            .in0(_gnd_net_),
            .in1(N__64218),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.genclk.div_state_1__N_1480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_clear_304_LC_20_7_0.C_ON=1'b0;
    defparam comm_clear_304_LC_20_7_0.SEQ_MODE=4'b1000;
    defparam comm_clear_304_LC_20_7_0.LUT_INIT=16'b0111011101010101;
    LogicCell40 comm_clear_304_LC_20_7_0 (
            .in0(N__62450),
            .in1(N__63602),
            .in2(_gnd_net_),
            .in3(N__63072),
            .lcout(comm_clear),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61880),
            .ce(N__56896),
            .sr(_gnd_net_));
    defparam i7121_2_lut_LC_20_8_1.C_ON=1'b0;
    defparam i7121_2_lut_LC_20_8_1.SEQ_MODE=4'b0000;
    defparam i7121_2_lut_LC_20_8_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 i7121_2_lut_LC_20_8_1 (
            .in0(_gnd_net_),
            .in1(N__62240),
            .in2(_gnd_net_),
            .in3(N__63966),
            .lcout(n9837),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20104_2_lut_LC_20_8_2.C_ON=1'b0;
    defparam i20104_2_lut_LC_20_8_2.SEQ_MODE=4'b0000;
    defparam i20104_2_lut_LC_20_8_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i20104_2_lut_LC_20_8_2 (
            .in0(_gnd_net_),
            .in1(N__56926),
            .in2(_gnd_net_),
            .in3(N__59420),
            .lcout(n22170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_adj_144_LC_20_8_5.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_144_LC_20_8_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_144_LC_20_8_5.LUT_INIT=16'b1110111011111111;
    LogicCell40 i2_2_lut_3_lut_adj_144_LC_20_8_5 (
            .in0(N__63028),
            .in1(N__62242),
            .in2(_gnd_net_),
            .in3(N__63488),
            .lcout(n12035),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i22_3_lut_4_lut_LC_20_8_6.C_ON=1'b0;
    defparam i22_3_lut_4_lut_LC_20_8_6.SEQ_MODE=4'b0000;
    defparam i22_3_lut_4_lut_LC_20_8_6.LUT_INIT=16'b0100011001000100;
    LogicCell40 i22_3_lut_4_lut_LC_20_8_6 (
            .in0(N__62241),
            .in1(N__63027),
            .in2(N__58132),
            .in3(N__58031),
            .lcout(n7_adj_1687),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_346_Mux_1_i8_3_lut_4_lut_LC_20_9_0.C_ON=1'b0;
    defparam comm_state_3__I_0_346_Mux_1_i8_3_lut_4_lut_LC_20_9_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_346_Mux_1_i8_3_lut_4_lut_LC_20_9_0.LUT_INIT=16'b0101001100000011;
    LogicCell40 comm_state_3__I_0_346_Mux_1_i8_3_lut_4_lut_LC_20_9_0 (
            .in0(N__57907),
            .in1(N__56875),
            .in2(N__63085),
            .in3(N__62296),
            .lcout(n8_adj_1659),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i228_2_lut_LC_20_9_2.C_ON=1'b0;
    defparam i228_2_lut_LC_20_9_2.SEQ_MODE=4'b0000;
    defparam i228_2_lut_LC_20_9_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i228_2_lut_LC_20_9_2 (
            .in0(_gnd_net_),
            .in1(N__58186),
            .in2(_gnd_net_),
            .in3(N__58022),
            .lcout(n1373),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_346_Mux_1_i2_3_lut_4_lut_LC_20_9_3.C_ON=1'b0;
    defparam comm_state_3__I_0_346_Mux_1_i2_3_lut_4_lut_LC_20_9_3.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_346_Mux_1_i2_3_lut_4_lut_LC_20_9_3.LUT_INIT=16'b0011000010111000;
    LogicCell40 comm_state_3__I_0_346_Mux_1_i2_3_lut_4_lut_LC_20_9_3 (
            .in0(N__62297),
            .in1(N__63070),
            .in2(N__58205),
            .in3(N__57906),
            .lcout(),
            .ltout(n2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23342_bdd_4_lut_LC_20_9_4.C_ON=1'b0;
    defparam n23342_bdd_4_lut_LC_20_9_4.SEQ_MODE=4'b0000;
    defparam n23342_bdd_4_lut_LC_20_9_4.LUT_INIT=16'b1111110000100010;
    LogicCell40 n23342_bdd_4_lut_LC_20_9_4 (
            .in0(N__63071),
            .in1(N__63910),
            .in2(N__57892),
            .in3(N__57889),
            .lcout(),
            .ltout(n23345_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i1_LC_20_9_5.C_ON=1'b0;
    defparam comm_state_i1_LC_20_9_5.SEQ_MODE=4'b1000;
    defparam comm_state_i1_LC_20_9_5.LUT_INIT=16'b0111010000110000;
    LogicCell40 comm_state_i1_LC_20_9_5 (
            .in0(N__57468),
            .in1(N__63540),
            .in2(N__57367),
            .in3(N__57364),
            .lcout(comm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61908),
            .ce(N__57325),
            .sr(_gnd_net_));
    defparam i20047_4_lut_LC_20_9_6.C_ON=1'b0;
    defparam i20047_4_lut_LC_20_9_6.SEQ_MODE=4'b0000;
    defparam i20047_4_lut_LC_20_9_6.LUT_INIT=16'b0101010000000100;
    LogicCell40 i20047_4_lut_LC_20_9_6 (
            .in0(N__62293),
            .in1(N__58185),
            .in2(N__64029),
            .in3(N__57358),
            .lcout(),
            .ltout(n22340_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20168_4_lut_LC_20_9_7.C_ON=1'b0;
    defparam i20168_4_lut_LC_20_9_7.SEQ_MODE=4'b0000;
    defparam i20168_4_lut_LC_20_9_7.LUT_INIT=16'b1100111111011101;
    LogicCell40 i20168_4_lut_LC_20_9_7 (
            .in0(N__57337),
            .in1(N__63539),
            .in2(N__57328),
            .in3(N__63066),
            .lcout(n14_adj_1593),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19903_2_lut_3_lut_LC_20_10_0.C_ON=1'b0;
    defparam i19903_2_lut_3_lut_LC_20_10_0.SEQ_MODE=4'b0000;
    defparam i19903_2_lut_3_lut_LC_20_10_0.LUT_INIT=16'b0011001000110010;
    LogicCell40 i19903_2_lut_3_lut_LC_20_10_0 (
            .in0(N__58035),
            .in1(N__63059),
            .in2(N__63987),
            .in3(_gnd_net_),
            .lcout(n22492),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7001_3_lut_4_lut_LC_20_10_1.C_ON=1'b0;
    defparam i7001_3_lut_4_lut_LC_20_10_1.SEQ_MODE=4'b0000;
    defparam i7001_3_lut_4_lut_LC_20_10_1.LUT_INIT=16'b1111010111100100;
    LogicCell40 i7001_3_lut_4_lut_LC_20_10_1 (
            .in0(N__63060),
            .in1(N__63908),
            .in2(N__57310),
            .in3(N__58032),
            .lcout(),
            .ltout(n9725_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_346_Mux_2_i6_4_lut_LC_20_10_2.C_ON=1'b0;
    defparam comm_state_3__I_0_346_Mux_2_i6_4_lut_LC_20_10_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_346_Mux_2_i6_4_lut_LC_20_10_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_state_3__I_0_346_Mux_2_i6_4_lut_LC_20_10_2 (
            .in0(N__62292),
            .in1(N__58187),
            .in2(N__57283),
            .in3(N__57280),
            .lcout(),
            .ltout(n6_adj_1657_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i2_LC_20_10_3.C_ON=1'b0;
    defparam comm_state_i2_LC_20_10_3.SEQ_MODE=4'b1000;
    defparam comm_state_i2_LC_20_10_3.LUT_INIT=16'b1111000010001000;
    LogicCell40 comm_state_i2_LC_20_10_3 (
            .in0(N__58216),
            .in1(N__58237),
            .in2(N__58231),
            .in3(N__63909),
            .lcout(comm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61921),
            .ce(N__58225),
            .sr(N__63617));
    defparam i1_4_lut_adj_283_LC_20_10_4.C_ON=1'b0;
    defparam i1_4_lut_adj_283_LC_20_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_283_LC_20_10_4.LUT_INIT=16'b0000101100101100;
    LogicCell40 i1_4_lut_adj_283_LC_20_10_4 (
            .in0(N__58034),
            .in1(N__58192),
            .in2(N__63986),
            .in3(N__62294),
            .lcout(),
            .ltout(n26_adj_1597_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20171_2_lut_3_lut_LC_20_10_5.C_ON=1'b0;
    defparam i20171_2_lut_3_lut_LC_20_10_5.SEQ_MODE=4'b0000;
    defparam i20171_2_lut_3_lut_LC_20_10_5.LUT_INIT=16'b1111111101011111;
    LogicCell40 i20171_2_lut_3_lut_LC_20_10_5 (
            .in0(N__63058),
            .in1(_gnd_net_),
            .in2(N__58228),
            .in3(N__63541),
            .lcout(n18_adj_1595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_147_LC_20_10_6.C_ON=1'b0;
    defparam i1_2_lut_adj_147_LC_20_10_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_147_LC_20_10_6.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_147_LC_20_10_6 (
            .in0(_gnd_net_),
            .in1(N__58188),
            .in2(_gnd_net_),
            .in3(N__62295),
            .lcout(n21908),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_281_LC_20_10_7.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_281_LC_20_10_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_281_LC_20_10_7.LUT_INIT=16'b0111011111110011;
    LogicCell40 i1_4_lut_4_lut_adj_281_LC_20_10_7 (
            .in0(N__63057),
            .in1(N__62291),
            .in2(N__58206),
            .in3(N__58033),
            .lcout(n4_adj_1718),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20087_2_lut_LC_20_11_0.C_ON=1'b0;
    defparam i20087_2_lut_LC_20_11_0.SEQ_MODE=4'b0000;
    defparam i20087_2_lut_LC_20_11_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 i20087_2_lut_LC_20_11_0 (
            .in0(_gnd_net_),
            .in1(N__58915),
            .in2(_gnd_net_),
            .in3(N__57958),
            .lcout(n22642),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_5_i127_3_lut_LC_20_11_6.C_ON=1'b0;
    defparam mux_125_Mux_5_i127_3_lut_LC_20_11_6.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_5_i127_3_lut_LC_20_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_125_Mux_5_i127_3_lut_LC_20_11_6 (
            .in0(N__57937),
            .in1(N__58318),
            .in2(_gnd_net_),
            .in3(N__61406),
            .lcout(comm_buf_0_7_N_543_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_300_LC_20_12_0.C_ON=1'b0;
    defparam i1_4_lut_adj_300_LC_20_12_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_300_LC_20_12_0.LUT_INIT=16'b1110001011111011;
    LogicCell40 i1_4_lut_adj_300_LC_20_12_0 (
            .in0(N__59421),
            .in1(N__61034),
            .in2(N__60044),
            .in3(N__60499),
            .lcout(n48),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19784_2_lut_3_lut_4_lut_LC_20_12_2.C_ON=1'b0;
    defparam i19784_2_lut_3_lut_4_lut_LC_20_12_2.SEQ_MODE=4'b0000;
    defparam i19784_2_lut_3_lut_4_lut_LC_20_12_2.LUT_INIT=16'b0000000000001000;
    LogicCell40 i19784_2_lut_3_lut_4_lut_LC_20_12_2 (
            .in0(N__58653),
            .in1(N__58492),
            .in2(N__60043),
            .in3(N__61033),
            .lcout(n22365),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19803_3_lut_4_lut_LC_20_12_3.C_ON=1'b0;
    defparam i19803_3_lut_4_lut_LC_20_12_3.SEQ_MODE=4'b0000;
    defparam i19803_3_lut_4_lut_LC_20_12_3.LUT_INIT=16'b0000000000100000;
    LogicCell40 i19803_3_lut_4_lut_LC_20_12_3 (
            .in0(N__61035),
            .in1(N__58654),
            .in2(N__58511),
            .in3(N__59423),
            .lcout(),
            .ltout(n22364_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20094_4_lut_LC_20_12_4.C_ON=1'b0;
    defparam i20094_4_lut_LC_20_12_4.SEQ_MODE=4'b0000;
    defparam i20094_4_lut_LC_20_12_4.LUT_INIT=16'b1011100000000000;
    LogicCell40 i20094_4_lut_LC_20_12_4 (
            .in0(N__58429),
            .in1(N__61374),
            .in2(N__58423),
            .in3(N__60501),
            .lcout(),
            .ltout(n22370_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19802_4_lut_LC_20_12_5.C_ON=1'b0;
    defparam i19802_4_lut_LC_20_12_5.SEQ_MODE=4'b0000;
    defparam i19802_4_lut_LC_20_12_5.LUT_INIT=16'b1111010011110000;
    LogicCell40 i19802_4_lut_LC_20_12_5 (
            .in0(N__61375),
            .in1(N__58420),
            .in2(N__58414),
            .in3(N__58407),
            .lcout(n22368),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_185_i9_2_lut_3_lut_LC_20_12_6.C_ON=1'b0;
    defparam equal_185_i9_2_lut_3_lut_LC_20_12_6.SEQ_MODE=4'b0000;
    defparam equal_185_i9_2_lut_3_lut_LC_20_12_6.LUT_INIT=16'b1110111011111111;
    LogicCell40 equal_185_i9_2_lut_3_lut_LC_20_12_6 (
            .in0(N__59422),
            .in1(N__59954),
            .in2(_gnd_net_),
            .in3(N__60500),
            .lcout(n9_adj_1507),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23492_bdd_4_lut_LC_20_12_7.C_ON=1'b0;
    defparam n23492_bdd_4_lut_LC_20_12_7.SEQ_MODE=4'b0000;
    defparam n23492_bdd_4_lut_LC_20_12_7.LUT_INIT=16'b1110111001010000;
    LogicCell40 n23492_bdd_4_lut_LC_20_12_7 (
            .in0(N__61036),
            .in1(N__58348),
            .in2(N__58330),
            .in3(N__60721),
            .lcout(n23495),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19755_2_lut_LC_20_13_5.C_ON=1'b0;
    defparam i19755_2_lut_LC_20_13_5.SEQ_MODE=4'b0000;
    defparam i19755_2_lut_LC_20_13_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i19755_2_lut_LC_20_13_5 (
            .in0(_gnd_net_),
            .in1(N__58312),
            .in2(_gnd_net_),
            .in3(N__59424),
            .lcout(n22316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n23456_bdd_4_lut_LC_20_14_1.C_ON=1'b0;
    defparam n23456_bdd_4_lut_LC_20_14_1.SEQ_MODE=4'b0000;
    defparam n23456_bdd_4_lut_LC_20_14_1.LUT_INIT=16'b1110111001010000;
    LogicCell40 n23456_bdd_4_lut_LC_20_14_1 (
            .in0(N__60093),
            .in1(N__58300),
            .in2(N__58291),
            .in3(N__59566),
            .lcout(),
            .ltout(n23459_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1661462_i1_3_lut_LC_20_14_2.C_ON=1'b0;
    defparam i1661462_i1_3_lut_LC_20_14_2.SEQ_MODE=4'b0000;
    defparam i1661462_i1_3_lut_LC_20_14_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1661462_i1_3_lut_LC_20_14_2 (
            .in0(_gnd_net_),
            .in1(N__58276),
            .in2(N__58258),
            .in3(N__61020),
            .lcout(),
            .ltout(n30_adj_1793_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_3_i127_3_lut_LC_20_14_3.C_ON=1'b0;
    defparam mux_125_Mux_3_i127_3_lut_LC_20_14_3.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_3_i127_3_lut_LC_20_14_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_125_Mux_3_i127_3_lut_LC_20_14_3 (
            .in0(_gnd_net_),
            .in1(N__58255),
            .in2(N__61417),
            .in3(N__61410),
            .lcout(comm_buf_0_7_N_543_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_5_i28_4_lut_LC_20_14_5.C_ON=1'b0;
    defparam mux_125_Mux_5_i28_4_lut_LC_20_14_5.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_5_i28_4_lut_LC_20_14_5.LUT_INIT=16'b0110001001000000;
    LogicCell40 mux_125_Mux_5_i28_4_lut_LC_20_14_5 (
            .in0(N__60601),
            .in1(N__59406),
            .in2(N__61102),
            .in3(N__61075),
            .lcout(),
            .ltout(n28_adj_1775_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_LC_20_14_6.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_LC_20_14_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_LC_20_14_6.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_2__bdd_4_lut_LC_20_14_6 (
            .in0(N__60676),
            .in1(N__60092),
            .in2(N__61060),
            .in3(N__61019),
            .lcout(n23492),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_125_Mux_5_i25_4_lut_LC_20_14_7.C_ON=1'b0;
    defparam mux_125_Mux_5_i25_4_lut_LC_20_14_7.SEQ_MODE=4'b0000;
    defparam mux_125_Mux_5_i25_4_lut_LC_20_14_7.LUT_INIT=16'b0111001001010000;
    LogicCell40 mux_125_Mux_5_i25_4_lut_LC_20_14_7 (
            .in0(N__60600),
            .in1(N__59405),
            .in2(N__60712),
            .in3(N__60697),
            .lcout(n25_adj_1774),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_20508_LC_20_15_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_20508_LC_20_15_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_20508_LC_20_15_5.LUT_INIT=16'b1110011010100010;
    LogicCell40 comm_cmd_1__bdd_4_lut_20508_LC_20_15_5 (
            .in0(N__60602),
            .in1(N__60064),
            .in2(N__59584),
            .in3(N__59572),
            .lcout(n23456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19937_2_lut_LC_20_15_6.C_ON=1'b0;
    defparam i19937_2_lut_LC_20_15_6.SEQ_MODE=4'b0000;
    defparam i19937_2_lut_LC_20_15_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i19937_2_lut_LC_20_15_6 (
            .in0(_gnd_net_),
            .in1(N__59560),
            .in2(_gnd_net_),
            .in3(N__59501),
            .lcout(n22313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19751_2_lut_LC_20_17_3.C_ON=1'b0;
    defparam i19751_2_lut_LC_20_17_3.SEQ_MODE=4'b0000;
    defparam i19751_2_lut_LC_20_17_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19751_2_lut_LC_20_17_3 (
            .in0(_gnd_net_),
            .in1(N__59542),
            .in2(_gnd_net_),
            .in3(N__59407),
            .lcout(n22300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20099_2_lut_LC_20_18_2.C_ON=1'b0;
    defparam i20099_2_lut_LC_20_18_2.SEQ_MODE=4'b0000;
    defparam i20099_2_lut_LC_20_18_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i20099_2_lut_LC_20_18_2 (
            .in0(_gnd_net_),
            .in1(N__59527),
            .in2(_gnd_net_),
            .in3(N__59496),
            .lcout(n22649),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_LC_22_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_22_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_22_5_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_LC_22_5_2  (
            .in0(N__64902),
            .in1(N__64341),
            .in2(N__64984),
            .in3(N__64302),
            .lcout(\ADC_VDC.genclk.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_LC_22_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_22_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_22_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_LC_22_5_3  (
            .in0(N__64917),
            .in1(N__64359),
            .in2(N__64270),
            .in3(N__64947),
            .lcout(\ADC_VDC.genclk.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i20011_4_lut_LC_22_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i20011_4_lut_LC_22_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i20011_4_lut_LC_22_5_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i20011_4_lut_LC_22_5_5  (
            .in0(N__64284),
            .in1(N__64377),
            .in2(N__64327),
            .in3(N__64392),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n22305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19909_4_lut_LC_22_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19909_4_lut_LC_22_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19909_4_lut_LC_22_5_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i19909_4_lut_LC_22_5_6  (
            .in0(N__64138),
            .in1(N__64252),
            .in2(N__64246),
            .in3(N__64243),
            .lcout(\ADC_VDC.genclk.n22303 ),
            .ltout(\ADC_VDC.genclk.n22303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i0_LC_22_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i0_LC_22_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i0_LC_22_5_7 .LUT_INIT=16'b1111011111010101;
    LogicCell40 \ADC_VDC.genclk.div_state_i0_LC_22_5_7  (
            .in0(N__64161),
            .in1(N__64228),
            .in2(N__64189),
            .in3(N__64186),
            .lcout(\ADC_VDC.genclk.div_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_LC_22_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_22_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_22_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_LC_22_6_4  (
            .in0(N__64887),
            .in1(N__64962),
            .in2(N__64498),
            .in3(N__64932),
            .lcout(\ADC_VDC.genclk.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_response_305_LC_22_8_7.C_ON=1'b0;
    defparam comm_response_305_LC_22_8_7.SEQ_MODE=4'b1000;
    defparam comm_response_305_LC_22_8_7.LUT_INIT=16'b0000010000110100;
    LogicCell40 comm_response_305_LC_22_8_7 (
            .in0(N__64025),
            .in1(N__63491),
            .in2(N__62633),
            .in3(N__63077),
            .lcout(ICE_GPMI_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61924),
            .ce(N__62803),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_22_10_5.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_22_10_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_22_10_5.LUT_INIT=16'b1101110111010000;
    LogicCell40 i1_3_lut_4_lut_LC_22_10_5 (
            .in0(N__63959),
            .in1(N__63722),
            .in2(N__63205),
            .in3(N__63074),
            .lcout(n12045),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i3_LC_22_11_4.C_ON=1'b0;
    defparam comm_buf_0__i3_LC_22_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i3_LC_22_11_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i3_LC_22_11_4 (
            .in0(N__62780),
            .in1(N__62602),
            .in2(_gnd_net_),
            .in3(N__62113),
            .lcout(comm_buf_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__61976),
            .ce(N__61437),
            .sr(N__64416));
    defparam \ADC_VDC.genclk.t0off_i0_LC_23_5_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i0_LC_23_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i0_LC_23_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i0_LC_23_5_0  (
            .in0(_gnd_net_),
            .in1(N__64393),
            .in2(_gnd_net_),
            .in3(N__64381),
            .lcout(\ADC_VDC.genclk.t0off_0 ),
            .ltout(),
            .carryin(bfn_23_5_0_),
            .carryout(\ADC_VDC.genclk.n20736 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i1_LC_23_5_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i1_LC_23_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i1_LC_23_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i1_LC_23_5_1  (
            .in0(_gnd_net_),
            .in1(N__64378),
            .in2(N__64848),
            .in3(N__64366),
            .lcout(\ADC_VDC.genclk.t0off_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20736 ),
            .carryout(\ADC_VDC.genclk.n20737 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i2_LC_23_5_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i2_LC_23_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i2_LC_23_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i2_LC_23_5_2  (
            .in0(_gnd_net_),
            .in1(N__64795),
            .in2(N__64363),
            .in3(N__64345),
            .lcout(\ADC_VDC.genclk.t0off_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20737 ),
            .carryout(\ADC_VDC.genclk.n20738 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i3_LC_23_5_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i3_LC_23_5_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0off_i3_LC_23_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i3_LC_23_5_3  (
            .in0(_gnd_net_),
            .in1(N__64342),
            .in2(N__64849),
            .in3(N__64330),
            .lcout(\ADC_VDC.genclk.t0off_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20738 ),
            .carryout(\ADC_VDC.genclk.n20739 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i4_LC_23_5_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i4_LC_23_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i4_LC_23_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i4_LC_23_5_4  (
            .in0(_gnd_net_),
            .in1(N__64799),
            .in2(N__64326),
            .in3(N__64306),
            .lcout(\ADC_VDC.genclk.t0off_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20739 ),
            .carryout(\ADC_VDC.genclk.n20740 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i5_LC_23_5_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i5_LC_23_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i5_LC_23_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i5_LC_23_5_5  (
            .in0(_gnd_net_),
            .in1(N__64303),
            .in2(N__64850),
            .in3(N__64291),
            .lcout(\ADC_VDC.genclk.t0off_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20740 ),
            .carryout(\ADC_VDC.genclk.n20741 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i6_LC_23_5_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i6_LC_23_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i6_LC_23_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i6_LC_23_5_6  (
            .in0(_gnd_net_),
            .in1(N__64803),
            .in2(N__64288),
            .in3(N__64273),
            .lcout(\ADC_VDC.genclk.t0off_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20741 ),
            .carryout(\ADC_VDC.genclk.n20742 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i7_LC_23_5_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i7_LC_23_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i7_LC_23_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i7_LC_23_5_7  (
            .in0(_gnd_net_),
            .in1(N__64269),
            .in2(N__64851),
            .in3(N__64255),
            .lcout(\ADC_VDC.genclk.t0off_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20742 ),
            .carryout(\ADC_VDC.genclk.n20743 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__64479),
            .sr(N__64459));
    defparam \ADC_VDC.genclk.t0off_i8_LC_23_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i8_LC_23_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i8_LC_23_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i8_LC_23_6_0  (
            .in0(_gnd_net_),
            .in1(N__64980),
            .in2(N__64730),
            .in3(N__64966),
            .lcout(\ADC_VDC.genclk.t0off_8 ),
            .ltout(),
            .carryin(bfn_23_6_0_),
            .carryout(\ADC_VDC.genclk.n20744 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
    defparam \ADC_VDC.genclk.t0off_i9_LC_23_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i9_LC_23_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i9_LC_23_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i9_LC_23_6_1  (
            .in0(_gnd_net_),
            .in1(N__64963),
            .in2(N__64733),
            .in3(N__64951),
            .lcout(\ADC_VDC.genclk.t0off_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20744 ),
            .carryout(\ADC_VDC.genclk.n20745 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
    defparam \ADC_VDC.genclk.t0off_i10_LC_23_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i10_LC_23_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i10_LC_23_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i10_LC_23_6_2  (
            .in0(_gnd_net_),
            .in1(N__64948),
            .in2(N__64727),
            .in3(N__64936),
            .lcout(\ADC_VDC.genclk.t0off_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20745 ),
            .carryout(\ADC_VDC.genclk.n20746 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
    defparam \ADC_VDC.genclk.t0off_i11_LC_23_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i11_LC_23_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i11_LC_23_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i11_LC_23_6_3  (
            .in0(_gnd_net_),
            .in1(N__64933),
            .in2(N__64731),
            .in3(N__64921),
            .lcout(\ADC_VDC.genclk.t0off_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20746 ),
            .carryout(\ADC_VDC.genclk.n20747 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
    defparam \ADC_VDC.genclk.t0off_i12_LC_23_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i12_LC_23_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i12_LC_23_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i12_LC_23_6_4  (
            .in0(_gnd_net_),
            .in1(N__64918),
            .in2(N__64728),
            .in3(N__64906),
            .lcout(\ADC_VDC.genclk.t0off_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20747 ),
            .carryout(\ADC_VDC.genclk.n20748 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
    defparam \ADC_VDC.genclk.t0off_i13_LC_23_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i13_LC_23_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i13_LC_23_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i13_LC_23_6_5  (
            .in0(_gnd_net_),
            .in1(N__64903),
            .in2(N__64732),
            .in3(N__64891),
            .lcout(\ADC_VDC.genclk.t0off_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20748 ),
            .carryout(\ADC_VDC.genclk.n20749 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
    defparam \ADC_VDC.genclk.t0off_i14_LC_23_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i14_LC_23_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i14_LC_23_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i14_LC_23_6_6  (
            .in0(_gnd_net_),
            .in1(N__64888),
            .in2(N__64729),
            .in3(N__64876),
            .lcout(\ADC_VDC.genclk.t0off_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n20749 ),
            .carryout(\ADC_VDC.genclk.n20750 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
    defparam \ADC_VDC.genclk.t0off_i15_LC_23_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0off_i15_LC_23_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i15_LC_23_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0off_i15_LC_23_6_7  (
            .in0(N__64666),
            .in1(N__64497),
            .in2(_gnd_net_),
            .in3(N__64501),
            .lcout(\ADC_VDC.genclk.t0off_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__64483),
            .sr(N__64458));
endmodule // zim
