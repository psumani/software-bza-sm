// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 3 2023 14:37:23

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "zim" view "INTERFACE"

module zim (
    VAC_DRDY,
    IAC_FLT1,
    DDS_SCK,
    ICE_IOR_166,
    ICE_IOR_119,
    DDS_MOSI,
    VAC_MISO,
    DDS_MOSI1,
    ICE_IOR_146,
    VDC_CLK,
    ICE_IOT_222,
    IAC_CS,
    ICE_IOL_18B,
    ICE_IOL_13A,
    ICE_IOB_81,
    VAC_OSR1,
    IAC_MOSI,
    DDS_CS1,
    ICE_IOL_4B,
    ICE_IOB_94,
    VAC_CS,
    VAC_CLK,
    ICE_SPI_CE0,
    ICE_IOR_167,
    ICE_IOR_118,
    RTD_SDO,
    IAC_OSR0,
    VDC_SCLK,
    VAC_FLT1,
    ICE_SPI_MOSI,
    ICE_IOR_165,
    ICE_IOR_147,
    ICE_IOL_14A,
    ICE_IOL_13B,
    ICE_IOB_91,
    ICE_GPMO_0,
    DDS_RNG_0,
    VDC_RNG0,
    ICE_SPI_SCLK,
    ICE_IOR_152,
    ICE_IOL_12A,
    RTD_DRDY,
    ICE_SPI_MISO,
    ICE_IOT_177,
    ICE_IOR_141,
    ICE_IOB_80,
    ICE_IOB_102,
    ICE_GPMO_2,
    ICE_GPMI_0,
    IAC_MISO,
    VAC_OSR0,
    VAC_MOSI,
    TEST_LED,
    ICE_IOR_148,
    STAT_COMM,
    ICE_SYSCLK,
    ICE_IOR_161,
    ICE_IOB_95,
    ICE_IOB_82,
    ICE_IOB_104,
    IAC_CLK,
    DDS_CS,
    SELIRNG0,
    RTD_SDI,
    ICE_IOT_221,
    ICE_IOT_197,
    DDS_MCLK,
    RTD_SCLK,
    RTD_CS,
    ICE_IOR_137,
    IAC_OSR1,
    VAC_FLT0,
    ICE_IOR_144,
    ICE_IOR_128,
    ICE_GPMO_1,
    IAC_SCLK,
    EIS_SYNCCLK,
    ICE_IOR_139,
    ICE_IOL_4A,
    VAC_SCLK,
    THERMOSTAT,
    ICE_IOR_164,
    ICE_IOB_103,
    AMPV_POW,
    VDC_SDO,
    ICE_IOT_174,
    ICE_IOR_140,
    ICE_IOB_96,
    CONT_SD,
    AC_ADC_SYNC,
    SELIRNG1,
    ICE_IOL_12B,
    ICE_IOR_160,
    ICE_IOR_136,
    DDS_MCLK1,
    ICE_IOT_198,
    ICE_IOT_173,
    IAC_DRDY,
    ICE_IOT_178,
    ICE_IOR_138,
    ICE_IOR_120,
    IAC_FLT0,
    DDS_SCK1);

    input VAC_DRDY;
    output IAC_FLT1;
    output DDS_SCK;
    input ICE_IOR_166;
    input ICE_IOR_119;
    output DDS_MOSI;
    input VAC_MISO;
    output DDS_MOSI1;
    input ICE_IOR_146;
    output VDC_CLK;
    input ICE_IOT_222;
    output IAC_CS;
    input ICE_IOL_18B;
    input ICE_IOL_13A;
    input ICE_IOB_81;
    output VAC_OSR1;
    output IAC_MOSI;
    output DDS_CS1;
    input ICE_IOL_4B;
    input ICE_IOB_94;
    output VAC_CS;
    output VAC_CLK;
    input ICE_SPI_CE0;
    input ICE_IOR_167;
    input ICE_IOR_118;
    input RTD_SDO;
    output IAC_OSR0;
    output VDC_SCLK;
    output VAC_FLT1;
    input ICE_SPI_MOSI;
    input ICE_IOR_165;
    input ICE_IOR_147;
    input ICE_IOL_14A;
    input ICE_IOL_13B;
    input ICE_IOB_91;
    input ICE_GPMO_0;
    output DDS_RNG_0;
    output VDC_RNG0;
    input ICE_SPI_SCLK;
    input ICE_IOR_152;
    input ICE_IOL_12A;
    input RTD_DRDY;
    output ICE_SPI_MISO;
    input ICE_IOT_177;
    input ICE_IOR_141;
    input ICE_IOB_80;
    input ICE_IOB_102;
    input ICE_GPMO_2;
    output ICE_GPMI_0;
    input IAC_MISO;
    output VAC_OSR0;
    output VAC_MOSI;
    output TEST_LED;
    input ICE_IOR_148;
    output STAT_COMM;
    input ICE_SYSCLK;
    input ICE_IOR_161;
    input ICE_IOB_95;
    input ICE_IOB_82;
    input ICE_IOB_104;
    output IAC_CLK;
    output DDS_CS;
    output SELIRNG0;
    output RTD_SDI;
    input ICE_IOT_221;
    input ICE_IOT_197;
    output DDS_MCLK;
    output RTD_SCLK;
    output RTD_CS;
    input ICE_IOR_137;
    output IAC_OSR1;
    output VAC_FLT0;
    input ICE_IOR_144;
    input ICE_IOR_128;
    input ICE_GPMO_1;
    output IAC_SCLK;
    input EIS_SYNCCLK;
    input ICE_IOR_139;
    input ICE_IOL_4A;
    output VAC_SCLK;
    input THERMOSTAT;
    input ICE_IOR_164;
    input ICE_IOB_103;
    output AMPV_POW;
    input VDC_SDO;
    input ICE_IOT_174;
    input ICE_IOR_140;
    input ICE_IOB_96;
    output CONT_SD;
    output AC_ADC_SYNC;
    output SELIRNG1;
    input ICE_IOL_12B;
    input ICE_IOR_160;
    input ICE_IOR_136;
    output DDS_MCLK1;
    input ICE_IOT_198;
    input ICE_IOT_173;
    input IAC_DRDY;
    input ICE_IOT_178;
    input ICE_IOR_138;
    input ICE_IOR_120;
    output IAC_FLT0;
    output DDS_SCK1;

    wire N__59563;
    wire N__59562;
    wire N__59561;
    wire N__59554;
    wire N__59553;
    wire N__59552;
    wire N__59545;
    wire N__59544;
    wire N__59543;
    wire N__59536;
    wire N__59535;
    wire N__59534;
    wire N__59527;
    wire N__59526;
    wire N__59525;
    wire N__59518;
    wire N__59517;
    wire N__59516;
    wire N__59509;
    wire N__59508;
    wire N__59507;
    wire N__59500;
    wire N__59499;
    wire N__59498;
    wire N__59491;
    wire N__59490;
    wire N__59489;
    wire N__59482;
    wire N__59481;
    wire N__59480;
    wire N__59473;
    wire N__59472;
    wire N__59471;
    wire N__59464;
    wire N__59463;
    wire N__59462;
    wire N__59455;
    wire N__59454;
    wire N__59453;
    wire N__59446;
    wire N__59445;
    wire N__59444;
    wire N__59437;
    wire N__59436;
    wire N__59435;
    wire N__59428;
    wire N__59427;
    wire N__59426;
    wire N__59419;
    wire N__59418;
    wire N__59417;
    wire N__59410;
    wire N__59409;
    wire N__59408;
    wire N__59401;
    wire N__59400;
    wire N__59399;
    wire N__59392;
    wire N__59391;
    wire N__59390;
    wire N__59383;
    wire N__59382;
    wire N__59381;
    wire N__59374;
    wire N__59373;
    wire N__59372;
    wire N__59365;
    wire N__59364;
    wire N__59363;
    wire N__59356;
    wire N__59355;
    wire N__59354;
    wire N__59347;
    wire N__59346;
    wire N__59345;
    wire N__59338;
    wire N__59337;
    wire N__59336;
    wire N__59329;
    wire N__59328;
    wire N__59327;
    wire N__59320;
    wire N__59319;
    wire N__59318;
    wire N__59311;
    wire N__59310;
    wire N__59309;
    wire N__59302;
    wire N__59301;
    wire N__59300;
    wire N__59293;
    wire N__59292;
    wire N__59291;
    wire N__59284;
    wire N__59283;
    wire N__59282;
    wire N__59275;
    wire N__59274;
    wire N__59273;
    wire N__59266;
    wire N__59265;
    wire N__59264;
    wire N__59257;
    wire N__59256;
    wire N__59255;
    wire N__59248;
    wire N__59247;
    wire N__59246;
    wire N__59239;
    wire N__59238;
    wire N__59237;
    wire N__59230;
    wire N__59229;
    wire N__59228;
    wire N__59221;
    wire N__59220;
    wire N__59219;
    wire N__59212;
    wire N__59211;
    wire N__59210;
    wire N__59203;
    wire N__59202;
    wire N__59201;
    wire N__59194;
    wire N__59193;
    wire N__59192;
    wire N__59185;
    wire N__59184;
    wire N__59183;
    wire N__59176;
    wire N__59175;
    wire N__59174;
    wire N__59167;
    wire N__59166;
    wire N__59165;
    wire N__59158;
    wire N__59157;
    wire N__59156;
    wire N__59149;
    wire N__59148;
    wire N__59147;
    wire N__59140;
    wire N__59139;
    wire N__59138;
    wire N__59131;
    wire N__59130;
    wire N__59129;
    wire N__59122;
    wire N__59121;
    wire N__59120;
    wire N__59113;
    wire N__59112;
    wire N__59111;
    wire N__59104;
    wire N__59103;
    wire N__59102;
    wire N__59095;
    wire N__59094;
    wire N__59093;
    wire N__59086;
    wire N__59085;
    wire N__59084;
    wire N__59077;
    wire N__59076;
    wire N__59075;
    wire N__59068;
    wire N__59067;
    wire N__59066;
    wire N__59059;
    wire N__59058;
    wire N__59057;
    wire N__59050;
    wire N__59049;
    wire N__59048;
    wire N__59041;
    wire N__59040;
    wire N__59039;
    wire N__59032;
    wire N__59031;
    wire N__59030;
    wire N__59023;
    wire N__59022;
    wire N__59021;
    wire N__59014;
    wire N__59013;
    wire N__59012;
    wire N__59005;
    wire N__59004;
    wire N__59003;
    wire N__58996;
    wire N__58995;
    wire N__58994;
    wire N__58987;
    wire N__58986;
    wire N__58985;
    wire N__58978;
    wire N__58977;
    wire N__58976;
    wire N__58969;
    wire N__58968;
    wire N__58967;
    wire N__58960;
    wire N__58959;
    wire N__58958;
    wire N__58951;
    wire N__58950;
    wire N__58949;
    wire N__58942;
    wire N__58941;
    wire N__58940;
    wire N__58933;
    wire N__58932;
    wire N__58931;
    wire N__58924;
    wire N__58923;
    wire N__58922;
    wire N__58915;
    wire N__58914;
    wire N__58913;
    wire N__58906;
    wire N__58905;
    wire N__58904;
    wire N__58897;
    wire N__58896;
    wire N__58895;
    wire N__58888;
    wire N__58887;
    wire N__58886;
    wire N__58879;
    wire N__58878;
    wire N__58877;
    wire N__58870;
    wire N__58869;
    wire N__58868;
    wire N__58861;
    wire N__58860;
    wire N__58859;
    wire N__58852;
    wire N__58851;
    wire N__58850;
    wire N__58843;
    wire N__58842;
    wire N__58841;
    wire N__58834;
    wire N__58833;
    wire N__58832;
    wire N__58825;
    wire N__58824;
    wire N__58823;
    wire N__58816;
    wire N__58815;
    wire N__58814;
    wire N__58807;
    wire N__58806;
    wire N__58805;
    wire N__58798;
    wire N__58797;
    wire N__58796;
    wire N__58789;
    wire N__58788;
    wire N__58787;
    wire N__58780;
    wire N__58779;
    wire N__58778;
    wire N__58771;
    wire N__58770;
    wire N__58769;
    wire N__58762;
    wire N__58761;
    wire N__58760;
    wire N__58753;
    wire N__58752;
    wire N__58751;
    wire N__58744;
    wire N__58743;
    wire N__58742;
    wire N__58735;
    wire N__58734;
    wire N__58733;
    wire N__58726;
    wire N__58725;
    wire N__58724;
    wire N__58717;
    wire N__58716;
    wire N__58715;
    wire N__58708;
    wire N__58707;
    wire N__58706;
    wire N__58699;
    wire N__58698;
    wire N__58697;
    wire N__58690;
    wire N__58689;
    wire N__58688;
    wire N__58681;
    wire N__58680;
    wire N__58679;
    wire N__58672;
    wire N__58671;
    wire N__58670;
    wire N__58663;
    wire N__58662;
    wire N__58661;
    wire N__58654;
    wire N__58653;
    wire N__58652;
    wire N__58645;
    wire N__58644;
    wire N__58643;
    wire N__58626;
    wire N__58623;
    wire N__58622;
    wire N__58621;
    wire N__58620;
    wire N__58617;
    wire N__58616;
    wire N__58613;
    wire N__58612;
    wire N__58609;
    wire N__58608;
    wire N__58607;
    wire N__58592;
    wire N__58589;
    wire N__58586;
    wire N__58585;
    wire N__58584;
    wire N__58581;
    wire N__58580;
    wire N__58579;
    wire N__58578;
    wire N__58577;
    wire N__58576;
    wire N__58575;
    wire N__58574;
    wire N__58573;
    wire N__58570;
    wire N__58567;
    wire N__58566;
    wire N__58565;
    wire N__58564;
    wire N__58561;
    wire N__58560;
    wire N__58557;
    wire N__58554;
    wire N__58553;
    wire N__58550;
    wire N__58549;
    wire N__58546;
    wire N__58545;
    wire N__58542;
    wire N__58541;
    wire N__58538;
    wire N__58537;
    wire N__58534;
    wire N__58533;
    wire N__58530;
    wire N__58529;
    wire N__58526;
    wire N__58525;
    wire N__58524;
    wire N__58523;
    wire N__58522;
    wire N__58519;
    wire N__58516;
    wire N__58513;
    wire N__58510;
    wire N__58509;
    wire N__58508;
    wire N__58507;
    wire N__58504;
    wire N__58503;
    wire N__58502;
    wire N__58501;
    wire N__58500;
    wire N__58497;
    wire N__58494;
    wire N__58491;
    wire N__58476;
    wire N__58459;
    wire N__58456;
    wire N__58455;
    wire N__58452;
    wire N__58451;
    wire N__58448;
    wire N__58447;
    wire N__58444;
    wire N__58435;
    wire N__58432;
    wire N__58429;
    wire N__58428;
    wire N__58425;
    wire N__58424;
    wire N__58421;
    wire N__58420;
    wire N__58417;
    wire N__58416;
    wire N__58413;
    wire N__58412;
    wire N__58409;
    wire N__58408;
    wire N__58405;
    wire N__58400;
    wire N__58397;
    wire N__58394;
    wire N__58391;
    wire N__58376;
    wire N__58369;
    wire N__58366;
    wire N__58363;
    wire N__58360;
    wire N__58359;
    wire N__58356;
    wire N__58339;
    wire N__58336;
    wire N__58335;
    wire N__58326;
    wire N__58317;
    wire N__58314;
    wire N__58311;
    wire N__58308;
    wire N__58305;
    wire N__58302;
    wire N__58299;
    wire N__58294;
    wire N__58293;
    wire N__58288;
    wire N__58283;
    wire N__58278;
    wire N__58275;
    wire N__58266;
    wire N__58263;
    wire N__58260;
    wire N__58259;
    wire N__58258;
    wire N__58255;
    wire N__58252;
    wire N__58249;
    wire N__58244;
    wire N__58243;
    wire N__58240;
    wire N__58237;
    wire N__58234;
    wire N__58231;
    wire N__58226;
    wire N__58221;
    wire N__58218;
    wire N__58217;
    wire N__58214;
    wire N__58211;
    wire N__58206;
    wire N__58205;
    wire N__58202;
    wire N__58199;
    wire N__58194;
    wire N__58193;
    wire N__58190;
    wire N__58187;
    wire N__58184;
    wire N__58181;
    wire N__58176;
    wire N__58175;
    wire N__58172;
    wire N__58169;
    wire N__58164;
    wire N__58161;
    wire N__58160;
    wire N__58157;
    wire N__58154;
    wire N__58151;
    wire N__58148;
    wire N__58145;
    wire N__58142;
    wire N__58139;
    wire N__58136;
    wire N__58131;
    wire N__58130;
    wire N__58127;
    wire N__58124;
    wire N__58119;
    wire N__58116;
    wire N__58115;
    wire N__58112;
    wire N__58109;
    wire N__58104;
    wire N__58103;
    wire N__58100;
    wire N__58097;
    wire N__58094;
    wire N__58089;
    wire N__58088;
    wire N__58085;
    wire N__58082;
    wire N__58077;
    wire N__58074;
    wire N__58071;
    wire N__58070;
    wire N__58067;
    wire N__58064;
    wire N__58059;
    wire N__58056;
    wire N__58055;
    wire N__58052;
    wire N__58049;
    wire N__58044;
    wire N__58043;
    wire N__58040;
    wire N__58037;
    wire N__58034;
    wire N__58029;
    wire N__58028;
    wire N__58025;
    wire N__58022;
    wire N__58017;
    wire N__58014;
    wire N__58011;
    wire N__58010;
    wire N__58007;
    wire N__58006;
    wire N__58005;
    wire N__58004;
    wire N__58003;
    wire N__58002;
    wire N__57999;
    wire N__57996;
    wire N__57993;
    wire N__57986;
    wire N__57983;
    wire N__57978;
    wire N__57975;
    wire N__57972;
    wire N__57963;
    wire N__57960;
    wire N__57959;
    wire N__57956;
    wire N__57953;
    wire N__57950;
    wire N__57947;
    wire N__57944;
    wire N__57941;
    wire N__57936;
    wire N__57935;
    wire N__57932;
    wire N__57929;
    wire N__57924;
    wire N__57921;
    wire N__57920;
    wire N__57917;
    wire N__57914;
    wire N__57909;
    wire N__57908;
    wire N__57905;
    wire N__57902;
    wire N__57899;
    wire N__57894;
    wire N__57891;
    wire N__57890;
    wire N__57887;
    wire N__57884;
    wire N__57879;
    wire N__57876;
    wire N__57873;
    wire N__57870;
    wire N__57867;
    wire N__57864;
    wire N__57861;
    wire N__57858;
    wire N__57855;
    wire N__57852;
    wire N__57849;
    wire N__57846;
    wire N__57843;
    wire N__57840;
    wire N__57837;
    wire N__57834;
    wire N__57831;
    wire N__57828;
    wire N__57825;
    wire N__57824;
    wire N__57823;
    wire N__57822;
    wire N__57821;
    wire N__57820;
    wire N__57819;
    wire N__57818;
    wire N__57817;
    wire N__57816;
    wire N__57815;
    wire N__57814;
    wire N__57813;
    wire N__57812;
    wire N__57809;
    wire N__57808;
    wire N__57807;
    wire N__57806;
    wire N__57805;
    wire N__57804;
    wire N__57803;
    wire N__57802;
    wire N__57801;
    wire N__57800;
    wire N__57797;
    wire N__57796;
    wire N__57795;
    wire N__57794;
    wire N__57793;
    wire N__57792;
    wire N__57789;
    wire N__57788;
    wire N__57787;
    wire N__57786;
    wire N__57785;
    wire N__57784;
    wire N__57783;
    wire N__57782;
    wire N__57781;
    wire N__57780;
    wire N__57779;
    wire N__57778;
    wire N__57777;
    wire N__57776;
    wire N__57773;
    wire N__57770;
    wire N__57767;
    wire N__57764;
    wire N__57763;
    wire N__57760;
    wire N__57759;
    wire N__57758;
    wire N__57757;
    wire N__57756;
    wire N__57755;
    wire N__57754;
    wire N__57751;
    wire N__57750;
    wire N__57749;
    wire N__57748;
    wire N__57747;
    wire N__57744;
    wire N__57741;
    wire N__57740;
    wire N__57739;
    wire N__57738;
    wire N__57737;
    wire N__57736;
    wire N__57729;
    wire N__57724;
    wire N__57717;
    wire N__57714;
    wire N__57705;
    wire N__57702;
    wire N__57701;
    wire N__57700;
    wire N__57699;
    wire N__57698;
    wire N__57695;
    wire N__57690;
    wire N__57685;
    wire N__57682;
    wire N__57675;
    wire N__57672;
    wire N__57669;
    wire N__57668;
    wire N__57667;
    wire N__57666;
    wire N__57665;
    wire N__57662;
    wire N__57661;
    wire N__57658;
    wire N__57655;
    wire N__57654;
    wire N__57653;
    wire N__57652;
    wire N__57651;
    wire N__57648;
    wire N__57643;
    wire N__57642;
    wire N__57641;
    wire N__57638;
    wire N__57635;
    wire N__57632;
    wire N__57627;
    wire N__57626;
    wire N__57625;
    wire N__57624;
    wire N__57619;
    wire N__57618;
    wire N__57617;
    wire N__57616;
    wire N__57615;
    wire N__57614;
    wire N__57611;
    wire N__57608;
    wire N__57605;
    wire N__57604;
    wire N__57603;
    wire N__57600;
    wire N__57597;
    wire N__57594;
    wire N__57593;
    wire N__57592;
    wire N__57591;
    wire N__57590;
    wire N__57589;
    wire N__57588;
    wire N__57585;
    wire N__57582;
    wire N__57579;
    wire N__57576;
    wire N__57573;
    wire N__57572;
    wire N__57569;
    wire N__57564;
    wire N__57561;
    wire N__57558;
    wire N__57555;
    wire N__57554;
    wire N__57553;
    wire N__57550;
    wire N__57547;
    wire N__57544;
    wire N__57539;
    wire N__57532;
    wire N__57527;
    wire N__57524;
    wire N__57521;
    wire N__57508;
    wire N__57505;
    wire N__57500;
    wire N__57499;
    wire N__57498;
    wire N__57493;
    wire N__57490;
    wire N__57487;
    wire N__57484;
    wire N__57481;
    wire N__57478;
    wire N__57477;
    wire N__57476;
    wire N__57475;
    wire N__57474;
    wire N__57467;
    wire N__57462;
    wire N__57459;
    wire N__57456;
    wire N__57451;
    wire N__57446;
    wire N__57443;
    wire N__57440;
    wire N__57437;
    wire N__57434;
    wire N__57423;
    wire N__57416;
    wire N__57411;
    wire N__57404;
    wire N__57399;
    wire N__57394;
    wire N__57389;
    wire N__57388;
    wire N__57387;
    wire N__57386;
    wire N__57385;
    wire N__57384;
    wire N__57383;
    wire N__57382;
    wire N__57381;
    wire N__57370;
    wire N__57367;
    wire N__57362;
    wire N__57355;
    wire N__57352;
    wire N__57349;
    wire N__57346;
    wire N__57335;
    wire N__57330;
    wire N__57323;
    wire N__57320;
    wire N__57317;
    wire N__57312;
    wire N__57303;
    wire N__57300;
    wire N__57293;
    wire N__57288;
    wire N__57281;
    wire N__57278;
    wire N__57263;
    wire N__57262;
    wire N__57261;
    wire N__57258;
    wire N__57251;
    wire N__57246;
    wire N__57241;
    wire N__57232;
    wire N__57225;
    wire N__57222;
    wire N__57215;
    wire N__57208;
    wire N__57199;
    wire N__57186;
    wire N__57181;
    wire N__57156;
    wire N__57153;
    wire N__57150;
    wire N__57147;
    wire N__57144;
    wire N__57143;
    wire N__57140;
    wire N__57139;
    wire N__57138;
    wire N__57135;
    wire N__57134;
    wire N__57133;
    wire N__57132;
    wire N__57127;
    wire N__57126;
    wire N__57125;
    wire N__57124;
    wire N__57123;
    wire N__57122;
    wire N__57119;
    wire N__57118;
    wire N__57115;
    wire N__57110;
    wire N__57109;
    wire N__57108;
    wire N__57105;
    wire N__57102;
    wire N__57099;
    wire N__57098;
    wire N__57097;
    wire N__57096;
    wire N__57095;
    wire N__57094;
    wire N__57093;
    wire N__57092;
    wire N__57091;
    wire N__57090;
    wire N__57089;
    wire N__57088;
    wire N__57087;
    wire N__57082;
    wire N__57079;
    wire N__57076;
    wire N__57073;
    wire N__57070;
    wire N__57069;
    wire N__57068;
    wire N__57067;
    wire N__57066;
    wire N__57065;
    wire N__57064;
    wire N__57063;
    wire N__57062;
    wire N__57061;
    wire N__57060;
    wire N__57059;
    wire N__57056;
    wire N__57053;
    wire N__57050;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57038;
    wire N__57035;
    wire N__57032;
    wire N__57029;
    wire N__57028;
    wire N__57025;
    wire N__57024;
    wire N__57023;
    wire N__57022;
    wire N__57021;
    wire N__57016;
    wire N__57015;
    wire N__57014;
    wire N__57013;
    wire N__57008;
    wire N__57005;
    wire N__57004;
    wire N__57001;
    wire N__57000;
    wire N__56999;
    wire N__56996;
    wire N__56993;
    wire N__56992;
    wire N__56983;
    wire N__56980;
    wire N__56973;
    wire N__56968;
    wire N__56959;
    wire N__56958;
    wire N__56957;
    wire N__56956;
    wire N__56955;
    wire N__56954;
    wire N__56953;
    wire N__56948;
    wire N__56947;
    wire N__56946;
    wire N__56945;
    wire N__56940;
    wire N__56937;
    wire N__56936;
    wire N__56935;
    wire N__56934;
    wire N__56933;
    wire N__56932;
    wire N__56931;
    wire N__56930;
    wire N__56929;
    wire N__56928;
    wire N__56927;
    wire N__56926;
    wire N__56925;
    wire N__56924;
    wire N__56923;
    wire N__56920;
    wire N__56917;
    wire N__56914;
    wire N__56905;
    wire N__56902;
    wire N__56901;
    wire N__56900;
    wire N__56899;
    wire N__56888;
    wire N__56885;
    wire N__56878;
    wire N__56875;
    wire N__56872;
    wire N__56869;
    wire N__56868;
    wire N__56867;
    wire N__56866;
    wire N__56865;
    wire N__56864;
    wire N__56863;
    wire N__56860;
    wire N__56857;
    wire N__56854;
    wire N__56853;
    wire N__56852;
    wire N__56845;
    wire N__56842;
    wire N__56835;
    wire N__56832;
    wire N__56831;
    wire N__56830;
    wire N__56827;
    wire N__56826;
    wire N__56825;
    wire N__56824;
    wire N__56823;
    wire N__56822;
    wire N__56811;
    wire N__56808;
    wire N__56801;
    wire N__56796;
    wire N__56787;
    wire N__56778;
    wire N__56773;
    wire N__56768;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56752;
    wire N__56743;
    wire N__56732;
    wire N__56727;
    wire N__56724;
    wire N__56715;
    wire N__56708;
    wire N__56703;
    wire N__56694;
    wire N__56693;
    wire N__56692;
    wire N__56689;
    wire N__56686;
    wire N__56683;
    wire N__56676;
    wire N__56671;
    wire N__56668;
    wire N__56651;
    wire N__56640;
    wire N__56629;
    wire N__56626;
    wire N__56621;
    wire N__56598;
    wire N__56595;
    wire N__56594;
    wire N__56591;
    wire N__56588;
    wire N__56585;
    wire N__56582;
    wire N__56579;
    wire N__56576;
    wire N__56571;
    wire N__56568;
    wire N__56567;
    wire N__56564;
    wire N__56563;
    wire N__56562;
    wire N__56561;
    wire N__56560;
    wire N__56559;
    wire N__56558;
    wire N__56557;
    wire N__56556;
    wire N__56555;
    wire N__56554;
    wire N__56553;
    wire N__56552;
    wire N__56551;
    wire N__56550;
    wire N__56549;
    wire N__56548;
    wire N__56547;
    wire N__56546;
    wire N__56545;
    wire N__56544;
    wire N__56541;
    wire N__56540;
    wire N__56539;
    wire N__56532;
    wire N__56527;
    wire N__56520;
    wire N__56519;
    wire N__56518;
    wire N__56517;
    wire N__56516;
    wire N__56513;
    wire N__56512;
    wire N__56509;
    wire N__56506;
    wire N__56505;
    wire N__56504;
    wire N__56501;
    wire N__56500;
    wire N__56499;
    wire N__56498;
    wire N__56497;
    wire N__56494;
    wire N__56489;
    wire N__56488;
    wire N__56485;
    wire N__56484;
    wire N__56483;
    wire N__56482;
    wire N__56481;
    wire N__56480;
    wire N__56479;
    wire N__56478;
    wire N__56477;
    wire N__56476;
    wire N__56475;
    wire N__56474;
    wire N__56473;
    wire N__56472;
    wire N__56471;
    wire N__56468;
    wire N__56467;
    wire N__56466;
    wire N__56459;
    wire N__56456;
    wire N__56453;
    wire N__56452;
    wire N__56451;
    wire N__56450;
    wire N__56447;
    wire N__56446;
    wire N__56445;
    wire N__56442;
    wire N__56441;
    wire N__56440;
    wire N__56433;
    wire N__56430;
    wire N__56427;
    wire N__56424;
    wire N__56421;
    wire N__56420;
    wire N__56419;
    wire N__56414;
    wire N__56409;
    wire N__56406;
    wire N__56401;
    wire N__56400;
    wire N__56395;
    wire N__56390;
    wire N__56387;
    wire N__56384;
    wire N__56379;
    wire N__56364;
    wire N__56361;
    wire N__56358;
    wire N__56357;
    wire N__56356;
    wire N__56351;
    wire N__56348;
    wire N__56345;
    wire N__56344;
    wire N__56343;
    wire N__56334;
    wire N__56331;
    wire N__56328;
    wire N__56325;
    wire N__56322;
    wire N__56321;
    wire N__56320;
    wire N__56317;
    wire N__56316;
    wire N__56315;
    wire N__56312;
    wire N__56305;
    wire N__56298;
    wire N__56293;
    wire N__56292;
    wire N__56291;
    wire N__56288;
    wire N__56281;
    wire N__56278;
    wire N__56275;
    wire N__56272;
    wire N__56267;
    wire N__56264;
    wire N__56253;
    wire N__56250;
    wire N__56247;
    wire N__56240;
    wire N__56237;
    wire N__56232;
    wire N__56229;
    wire N__56228;
    wire N__56227;
    wire N__56224;
    wire N__56223;
    wire N__56222;
    wire N__56221;
    wire N__56220;
    wire N__56215;
    wire N__56212;
    wire N__56207;
    wire N__56204;
    wire N__56203;
    wire N__56202;
    wire N__56199;
    wire N__56196;
    wire N__56191;
    wire N__56188;
    wire N__56181;
    wire N__56180;
    wire N__56179;
    wire N__56176;
    wire N__56175;
    wire N__56174;
    wire N__56171;
    wire N__56170;
    wire N__56169;
    wire N__56168;
    wire N__56165;
    wire N__56160;
    wire N__56157;
    wire N__56146;
    wire N__56143;
    wire N__56136;
    wire N__56129;
    wire N__56124;
    wire N__56121;
    wire N__56116;
    wire N__56109;
    wire N__56100;
    wire N__56091;
    wire N__56084;
    wire N__56075;
    wire N__56070;
    wire N__56065;
    wire N__56054;
    wire N__56031;
    wire N__56030;
    wire N__56027;
    wire N__56024;
    wire N__56021;
    wire N__56018;
    wire N__56015;
    wire N__56010;
    wire N__56007;
    wire N__56004;
    wire N__56001;
    wire N__55998;
    wire N__55995;
    wire N__55992;
    wire N__55989;
    wire N__55986;
    wire N__55983;
    wire N__55980;
    wire N__55977;
    wire N__55974;
    wire N__55971;
    wire N__55968;
    wire N__55967;
    wire N__55964;
    wire N__55961;
    wire N__55958;
    wire N__55955;
    wire N__55952;
    wire N__55949;
    wire N__55946;
    wire N__55943;
    wire N__55940;
    wire N__55937;
    wire N__55934;
    wire N__55931;
    wire N__55928;
    wire N__55925;
    wire N__55922;
    wire N__55917;
    wire N__55914;
    wire N__55911;
    wire N__55908;
    wire N__55905;
    wire N__55902;
    wire N__55901;
    wire N__55900;
    wire N__55897;
    wire N__55894;
    wire N__55891;
    wire N__55888;
    wire N__55885;
    wire N__55882;
    wire N__55875;
    wire N__55874;
    wire N__55873;
    wire N__55872;
    wire N__55871;
    wire N__55870;
    wire N__55869;
    wire N__55868;
    wire N__55867;
    wire N__55866;
    wire N__55865;
    wire N__55862;
    wire N__55859;
    wire N__55858;
    wire N__55857;
    wire N__55854;
    wire N__55851;
    wire N__55850;
    wire N__55849;
    wire N__55848;
    wire N__55847;
    wire N__55844;
    wire N__55843;
    wire N__55840;
    wire N__55837;
    wire N__55834;
    wire N__55833;
    wire N__55832;
    wire N__55831;
    wire N__55828;
    wire N__55827;
    wire N__55824;
    wire N__55821;
    wire N__55820;
    wire N__55819;
    wire N__55818;
    wire N__55817;
    wire N__55816;
    wire N__55811;
    wire N__55810;
    wire N__55795;
    wire N__55792;
    wire N__55787;
    wire N__55782;
    wire N__55779;
    wire N__55778;
    wire N__55777;
    wire N__55772;
    wire N__55769;
    wire N__55766;
    wire N__55765;
    wire N__55764;
    wire N__55763;
    wire N__55760;
    wire N__55759;
    wire N__55758;
    wire N__55757;
    wire N__55752;
    wire N__55749;
    wire N__55742;
    wire N__55739;
    wire N__55736;
    wire N__55733;
    wire N__55730;
    wire N__55725;
    wire N__55720;
    wire N__55717;
    wire N__55714;
    wire N__55709;
    wire N__55706;
    wire N__55699;
    wire N__55696;
    wire N__55689;
    wire N__55680;
    wire N__55677;
    wire N__55674;
    wire N__55667;
    wire N__55656;
    wire N__55649;
    wire N__55638;
    wire N__55637;
    wire N__55636;
    wire N__55633;
    wire N__55630;
    wire N__55627;
    wire N__55624;
    wire N__55621;
    wire N__55618;
    wire N__55615;
    wire N__55614;
    wire N__55611;
    wire N__55608;
    wire N__55605;
    wire N__55602;
    wire N__55601;
    wire N__55598;
    wire N__55595;
    wire N__55590;
    wire N__55587;
    wire N__55578;
    wire N__55575;
    wire N__55572;
    wire N__55569;
    wire N__55566;
    wire N__55563;
    wire N__55560;
    wire N__55557;
    wire N__55556;
    wire N__55553;
    wire N__55552;
    wire N__55551;
    wire N__55550;
    wire N__55549;
    wire N__55548;
    wire N__55547;
    wire N__55546;
    wire N__55545;
    wire N__55544;
    wire N__55543;
    wire N__55542;
    wire N__55541;
    wire N__55538;
    wire N__55535;
    wire N__55526;
    wire N__55525;
    wire N__55524;
    wire N__55523;
    wire N__55522;
    wire N__55519;
    wire N__55518;
    wire N__55517;
    wire N__55516;
    wire N__55515;
    wire N__55514;
    wire N__55513;
    wire N__55512;
    wire N__55511;
    wire N__55510;
    wire N__55507;
    wire N__55504;
    wire N__55501;
    wire N__55500;
    wire N__55499;
    wire N__55492;
    wire N__55489;
    wire N__55486;
    wire N__55481;
    wire N__55480;
    wire N__55473;
    wire N__55470;
    wire N__55467;
    wire N__55464;
    wire N__55459;
    wire N__55452;
    wire N__55451;
    wire N__55448;
    wire N__55447;
    wire N__55444;
    wire N__55441;
    wire N__55434;
    wire N__55431;
    wire N__55430;
    wire N__55429;
    wire N__55426;
    wire N__55423;
    wire N__55422;
    wire N__55421;
    wire N__55418;
    wire N__55415;
    wire N__55412;
    wire N__55409;
    wire N__55408;
    wire N__55407;
    wire N__55406;
    wire N__55405;
    wire N__55404;
    wire N__55397;
    wire N__55394;
    wire N__55391;
    wire N__55388;
    wire N__55385;
    wire N__55380;
    wire N__55375;
    wire N__55370;
    wire N__55365;
    wire N__55360;
    wire N__55357;
    wire N__55354;
    wire N__55353;
    wire N__55352;
    wire N__55351;
    wire N__55350;
    wire N__55349;
    wire N__55348;
    wire N__55339;
    wire N__55336;
    wire N__55331;
    wire N__55326;
    wire N__55317;
    wire N__55314;
    wire N__55309;
    wire N__55302;
    wire N__55299;
    wire N__55296;
    wire N__55287;
    wire N__55282;
    wire N__55277;
    wire N__55270;
    wire N__55263;
    wire N__55248;
    wire N__55245;
    wire N__55242;
    wire N__55239;
    wire N__55236;
    wire N__55235;
    wire N__55234;
    wire N__55233;
    wire N__55232;
    wire N__55231;
    wire N__55230;
    wire N__55225;
    wire N__55220;
    wire N__55219;
    wire N__55218;
    wire N__55217;
    wire N__55216;
    wire N__55215;
    wire N__55214;
    wire N__55213;
    wire N__55212;
    wire N__55211;
    wire N__55210;
    wire N__55209;
    wire N__55208;
    wire N__55205;
    wire N__55200;
    wire N__55195;
    wire N__55190;
    wire N__55189;
    wire N__55188;
    wire N__55187;
    wire N__55184;
    wire N__55177;
    wire N__55176;
    wire N__55175;
    wire N__55174;
    wire N__55173;
    wire N__55172;
    wire N__55171;
    wire N__55170;
    wire N__55169;
    wire N__55166;
    wire N__55165;
    wire N__55164;
    wire N__55163;
    wire N__55162;
    wire N__55161;
    wire N__55160;
    wire N__55159;
    wire N__55158;
    wire N__55157;
    wire N__55156;
    wire N__55155;
    wire N__55154;
    wire N__55153;
    wire N__55152;
    wire N__55151;
    wire N__55150;
    wire N__55149;
    wire N__55148;
    wire N__55147;
    wire N__55146;
    wire N__55145;
    wire N__55142;
    wire N__55141;
    wire N__55140;
    wire N__55137;
    wire N__55136;
    wire N__55133;
    wire N__55132;
    wire N__55129;
    wire N__55126;
    wire N__55125;
    wire N__55116;
    wire N__55109;
    wire N__55104;
    wire N__55101;
    wire N__55098;
    wire N__55095;
    wire N__55092;
    wire N__55085;
    wire N__55082;
    wire N__55071;
    wire N__55066;
    wire N__55063;
    wire N__55060;
    wire N__55059;
    wire N__55058;
    wire N__55057;
    wire N__55056;
    wire N__55053;
    wire N__55050;
    wire N__55047;
    wire N__55042;
    wire N__55037;
    wire N__55036;
    wire N__55035;
    wire N__55034;
    wire N__55029;
    wire N__55026;
    wire N__55023;
    wire N__55022;
    wire N__55019;
    wire N__55012;
    wire N__55009;
    wire N__55006;
    wire N__55003;
    wire N__54996;
    wire N__54993;
    wire N__54990;
    wire N__54985;
    wire N__54980;
    wire N__54979;
    wire N__54978;
    wire N__54975;
    wire N__54968;
    wire N__54965;
    wire N__54962;
    wire N__54959;
    wire N__54956;
    wire N__54953;
    wire N__54950;
    wire N__54947;
    wire N__54944;
    wire N__54941;
    wire N__54930;
    wire N__54925;
    wire N__54922;
    wire N__54917;
    wire N__54914;
    wire N__54913;
    wire N__54910;
    wire N__54907;
    wire N__54904;
    wire N__54895;
    wire N__54892;
    wire N__54885;
    wire N__54884;
    wire N__54879;
    wire N__54874;
    wire N__54869;
    wire N__54868;
    wire N__54865;
    wire N__54860;
    wire N__54857;
    wire N__54852;
    wire N__54849;
    wire N__54838;
    wire N__54837;
    wire N__54836;
    wire N__54835;
    wire N__54832;
    wire N__54827;
    wire N__54818;
    wire N__54815;
    wire N__54808;
    wire N__54805;
    wire N__54800;
    wire N__54791;
    wire N__54784;
    wire N__54765;
    wire N__54764;
    wire N__54763;
    wire N__54762;
    wire N__54761;
    wire N__54760;
    wire N__54759;
    wire N__54758;
    wire N__54757;
    wire N__54756;
    wire N__54755;
    wire N__54754;
    wire N__54753;
    wire N__54750;
    wire N__54749;
    wire N__54748;
    wire N__54747;
    wire N__54746;
    wire N__54745;
    wire N__54744;
    wire N__54741;
    wire N__54738;
    wire N__54733;
    wire N__54728;
    wire N__54723;
    wire N__54720;
    wire N__54719;
    wire N__54716;
    wire N__54713;
    wire N__54712;
    wire N__54711;
    wire N__54708;
    wire N__54707;
    wire N__54706;
    wire N__54703;
    wire N__54698;
    wire N__54697;
    wire N__54696;
    wire N__54695;
    wire N__54694;
    wire N__54693;
    wire N__54692;
    wire N__54691;
    wire N__54688;
    wire N__54687;
    wire N__54686;
    wire N__54683;
    wire N__54680;
    wire N__54677;
    wire N__54672;
    wire N__54665;
    wire N__54662;
    wire N__54659;
    wire N__54654;
    wire N__54653;
    wire N__54648;
    wire N__54645;
    wire N__54644;
    wire N__54641;
    wire N__54638;
    wire N__54635;
    wire N__54632;
    wire N__54631;
    wire N__54628;
    wire N__54625;
    wire N__54622;
    wire N__54619;
    wire N__54614;
    wire N__54611;
    wire N__54608;
    wire N__54603;
    wire N__54602;
    wire N__54601;
    wire N__54598;
    wire N__54595;
    wire N__54588;
    wire N__54585;
    wire N__54582;
    wire N__54579;
    wire N__54576;
    wire N__54573;
    wire N__54570;
    wire N__54569;
    wire N__54566;
    wire N__54563;
    wire N__54558;
    wire N__54555;
    wire N__54554;
    wire N__54551;
    wire N__54546;
    wire N__54539;
    wire N__54532;
    wire N__54529;
    wire N__54526;
    wire N__54517;
    wire N__54512;
    wire N__54505;
    wire N__54502;
    wire N__54493;
    wire N__54490;
    wire N__54481;
    wire N__54478;
    wire N__54459;
    wire N__54456;
    wire N__54453;
    wire N__54450;
    wire N__54449;
    wire N__54446;
    wire N__54443;
    wire N__54438;
    wire N__54437;
    wire N__54436;
    wire N__54435;
    wire N__54434;
    wire N__54433;
    wire N__54432;
    wire N__54431;
    wire N__54430;
    wire N__54429;
    wire N__54428;
    wire N__54427;
    wire N__54426;
    wire N__54425;
    wire N__54424;
    wire N__54423;
    wire N__54422;
    wire N__54421;
    wire N__54420;
    wire N__54419;
    wire N__54418;
    wire N__54417;
    wire N__54416;
    wire N__54415;
    wire N__54414;
    wire N__54413;
    wire N__54412;
    wire N__54411;
    wire N__54410;
    wire N__54409;
    wire N__54408;
    wire N__54407;
    wire N__54406;
    wire N__54405;
    wire N__54404;
    wire N__54403;
    wire N__54402;
    wire N__54401;
    wire N__54400;
    wire N__54399;
    wire N__54398;
    wire N__54397;
    wire N__54396;
    wire N__54395;
    wire N__54394;
    wire N__54393;
    wire N__54392;
    wire N__54391;
    wire N__54390;
    wire N__54389;
    wire N__54388;
    wire N__54387;
    wire N__54386;
    wire N__54385;
    wire N__54384;
    wire N__54383;
    wire N__54382;
    wire N__54381;
    wire N__54380;
    wire N__54379;
    wire N__54378;
    wire N__54377;
    wire N__54376;
    wire N__54375;
    wire N__54374;
    wire N__54373;
    wire N__54372;
    wire N__54371;
    wire N__54370;
    wire N__54369;
    wire N__54368;
    wire N__54367;
    wire N__54366;
    wire N__54365;
    wire N__54364;
    wire N__54363;
    wire N__54362;
    wire N__54361;
    wire N__54360;
    wire N__54359;
    wire N__54358;
    wire N__54357;
    wire N__54356;
    wire N__54355;
    wire N__54354;
    wire N__54353;
    wire N__54352;
    wire N__54351;
    wire N__54350;
    wire N__54349;
    wire N__54348;
    wire N__54347;
    wire N__54346;
    wire N__54345;
    wire N__54344;
    wire N__54343;
    wire N__54342;
    wire N__54341;
    wire N__54340;
    wire N__54339;
    wire N__54338;
    wire N__54337;
    wire N__54336;
    wire N__54335;
    wire N__54334;
    wire N__54333;
    wire N__54332;
    wire N__54331;
    wire N__54330;
    wire N__54329;
    wire N__54328;
    wire N__54327;
    wire N__54326;
    wire N__54325;
    wire N__54324;
    wire N__54323;
    wire N__54322;
    wire N__54321;
    wire N__54320;
    wire N__54319;
    wire N__54318;
    wire N__54317;
    wire N__54316;
    wire N__54315;
    wire N__54314;
    wire N__54313;
    wire N__54312;
    wire N__54311;
    wire N__54310;
    wire N__54309;
    wire N__54308;
    wire N__54307;
    wire N__54306;
    wire N__54305;
    wire N__54304;
    wire N__54303;
    wire N__54302;
    wire N__54301;
    wire N__54300;
    wire N__54299;
    wire N__54298;
    wire N__54297;
    wire N__54296;
    wire N__54295;
    wire N__54294;
    wire N__54293;
    wire N__54292;
    wire N__54291;
    wire N__54290;
    wire N__54289;
    wire N__54288;
    wire N__54287;
    wire N__54286;
    wire N__54285;
    wire N__54284;
    wire N__54283;
    wire N__54282;
    wire N__54281;
    wire N__54280;
    wire N__54279;
    wire N__54278;
    wire N__54277;
    wire N__54276;
    wire N__54275;
    wire N__54274;
    wire N__54273;
    wire N__54272;
    wire N__54271;
    wire N__54270;
    wire N__54269;
    wire N__53928;
    wire N__53925;
    wire N__53924;
    wire N__53921;
    wire N__53918;
    wire N__53917;
    wire N__53914;
    wire N__53911;
    wire N__53908;
    wire N__53901;
    wire N__53898;
    wire N__53895;
    wire N__53892;
    wire N__53889;
    wire N__53886;
    wire N__53883;
    wire N__53880;
    wire N__53877;
    wire N__53874;
    wire N__53871;
    wire N__53868;
    wire N__53865;
    wire N__53862;
    wire N__53859;
    wire N__53856;
    wire N__53853;
    wire N__53850;
    wire N__53847;
    wire N__53844;
    wire N__53841;
    wire N__53838;
    wire N__53835;
    wire N__53832;
    wire N__53831;
    wire N__53828;
    wire N__53825;
    wire N__53822;
    wire N__53819;
    wire N__53814;
    wire N__53813;
    wire N__53810;
    wire N__53807;
    wire N__53804;
    wire N__53799;
    wire N__53798;
    wire N__53797;
    wire N__53796;
    wire N__53795;
    wire N__53794;
    wire N__53793;
    wire N__53792;
    wire N__53791;
    wire N__53790;
    wire N__53789;
    wire N__53788;
    wire N__53787;
    wire N__53786;
    wire N__53785;
    wire N__53784;
    wire N__53783;
    wire N__53782;
    wire N__53781;
    wire N__53780;
    wire N__53779;
    wire N__53778;
    wire N__53777;
    wire N__53772;
    wire N__53771;
    wire N__53768;
    wire N__53767;
    wire N__53766;
    wire N__53765;
    wire N__53764;
    wire N__53763;
    wire N__53762;
    wire N__53761;
    wire N__53758;
    wire N__53757;
    wire N__53756;
    wire N__53755;
    wire N__53754;
    wire N__53751;
    wire N__53750;
    wire N__53749;
    wire N__53746;
    wire N__53739;
    wire N__53730;
    wire N__53729;
    wire N__53728;
    wire N__53727;
    wire N__53724;
    wire N__53723;
    wire N__53722;
    wire N__53721;
    wire N__53720;
    wire N__53717;
    wire N__53710;
    wire N__53707;
    wire N__53704;
    wire N__53699;
    wire N__53696;
    wire N__53693;
    wire N__53690;
    wire N__53687;
    wire N__53684;
    wire N__53683;
    wire N__53682;
    wire N__53681;
    wire N__53680;
    wire N__53679;
    wire N__53676;
    wire N__53673;
    wire N__53672;
    wire N__53671;
    wire N__53670;
    wire N__53669;
    wire N__53668;
    wire N__53667;
    wire N__53666;
    wire N__53659;
    wire N__53654;
    wire N__53645;
    wire N__53642;
    wire N__53637;
    wire N__53634;
    wire N__53631;
    wire N__53628;
    wire N__53621;
    wire N__53618;
    wire N__53615;
    wire N__53614;
    wire N__53613;
    wire N__53612;
    wire N__53611;
    wire N__53608;
    wire N__53605;
    wire N__53602;
    wire N__53597;
    wire N__53590;
    wire N__53585;
    wire N__53580;
    wire N__53577;
    wire N__53568;
    wire N__53565;
    wire N__53562;
    wire N__53559;
    wire N__53556;
    wire N__53555;
    wire N__53554;
    wire N__53553;
    wire N__53552;
    wire N__53549;
    wire N__53548;
    wire N__53545;
    wire N__53536;
    wire N__53529;
    wire N__53526;
    wire N__53523;
    wire N__53520;
    wire N__53513;
    wire N__53510;
    wire N__53507;
    wire N__53502;
    wire N__53499;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53489;
    wire N__53486;
    wire N__53483;
    wire N__53480;
    wire N__53475;
    wire N__53472;
    wire N__53469;
    wire N__53466;
    wire N__53459;
    wire N__53458;
    wire N__53457;
    wire N__53454;
    wire N__53447;
    wire N__53444;
    wire N__53441;
    wire N__53430;
    wire N__53423;
    wire N__53420;
    wire N__53409;
    wire N__53406;
    wire N__53397;
    wire N__53388;
    wire N__53383;
    wire N__53358;
    wire N__53355;
    wire N__53352;
    wire N__53351;
    wire N__53348;
    wire N__53345;
    wire N__53342;
    wire N__53339;
    wire N__53334;
    wire N__53331;
    wire N__53328;
    wire N__53325;
    wire N__53324;
    wire N__53321;
    wire N__53320;
    wire N__53319;
    wire N__53318;
    wire N__53315;
    wire N__53312;
    wire N__53309;
    wire N__53306;
    wire N__53303;
    wire N__53302;
    wire N__53301;
    wire N__53300;
    wire N__53299;
    wire N__53298;
    wire N__53295;
    wire N__53294;
    wire N__53293;
    wire N__53288;
    wire N__53285;
    wire N__53282;
    wire N__53279;
    wire N__53278;
    wire N__53277;
    wire N__53276;
    wire N__53275;
    wire N__53272;
    wire N__53269;
    wire N__53266;
    wire N__53265;
    wire N__53262;
    wire N__53261;
    wire N__53260;
    wire N__53257;
    wire N__53256;
    wire N__53255;
    wire N__53254;
    wire N__53253;
    wire N__53250;
    wire N__53247;
    wire N__53244;
    wire N__53237;
    wire N__53234;
    wire N__53231;
    wire N__53228;
    wire N__53225;
    wire N__53220;
    wire N__53217;
    wire N__53214;
    wire N__53211;
    wire N__53208;
    wire N__53207;
    wire N__53204;
    wire N__53201;
    wire N__53198;
    wire N__53195;
    wire N__53194;
    wire N__53191;
    wire N__53188;
    wire N__53183;
    wire N__53176;
    wire N__53173;
    wire N__53168;
    wire N__53163;
    wire N__53160;
    wire N__53155;
    wire N__53152;
    wire N__53149;
    wire N__53142;
    wire N__53139;
    wire N__53132;
    wire N__53129;
    wire N__53124;
    wire N__53119;
    wire N__53114;
    wire N__53109;
    wire N__53106;
    wire N__53103;
    wire N__53100;
    wire N__53093;
    wire N__53088;
    wire N__53085;
    wire N__53082;
    wire N__53079;
    wire N__53076;
    wire N__53067;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53052;
    wire N__53051;
    wire N__53050;
    wire N__53047;
    wire N__53044;
    wire N__53041;
    wire N__53040;
    wire N__53039;
    wire N__53038;
    wire N__53037;
    wire N__53036;
    wire N__53035;
    wire N__53030;
    wire N__53027;
    wire N__53022;
    wire N__53019;
    wire N__53016;
    wire N__53013;
    wire N__53010;
    wire N__53007;
    wire N__53000;
    wire N__52995;
    wire N__52992;
    wire N__52989;
    wire N__52986;
    wire N__52983;
    wire N__52980;
    wire N__52971;
    wire N__52970;
    wire N__52969;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52953;
    wire N__52950;
    wire N__52949;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52939;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52923;
    wire N__52920;
    wire N__52917;
    wire N__52914;
    wire N__52911;
    wire N__52908;
    wire N__52907;
    wire N__52906;
    wire N__52901;
    wire N__52898;
    wire N__52895;
    wire N__52894;
    wire N__52893;
    wire N__52890;
    wire N__52887;
    wire N__52882;
    wire N__52875;
    wire N__52874;
    wire N__52871;
    wire N__52868;
    wire N__52863;
    wire N__52862;
    wire N__52859;
    wire N__52856;
    wire N__52851;
    wire N__52848;
    wire N__52845;
    wire N__52844;
    wire N__52841;
    wire N__52840;
    wire N__52837;
    wire N__52834;
    wire N__52831;
    wire N__52824;
    wire N__52821;
    wire N__52818;
    wire N__52815;
    wire N__52812;
    wire N__52811;
    wire N__52810;
    wire N__52807;
    wire N__52802;
    wire N__52797;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52787;
    wire N__52784;
    wire N__52781;
    wire N__52778;
    wire N__52775;
    wire N__52774;
    wire N__52771;
    wire N__52768;
    wire N__52765;
    wire N__52762;
    wire N__52759;
    wire N__52752;
    wire N__52749;
    wire N__52746;
    wire N__52743;
    wire N__52740;
    wire N__52737;
    wire N__52734;
    wire N__52731;
    wire N__52728;
    wire N__52725;
    wire N__52722;
    wire N__52719;
    wire N__52716;
    wire N__52713;
    wire N__52710;
    wire N__52707;
    wire N__52704;
    wire N__52701;
    wire N__52698;
    wire N__52695;
    wire N__52692;
    wire N__52689;
    wire N__52686;
    wire N__52683;
    wire N__52680;
    wire N__52677;
    wire N__52674;
    wire N__52671;
    wire N__52668;
    wire N__52665;
    wire N__52662;
    wire N__52659;
    wire N__52656;
    wire N__52653;
    wire N__52650;
    wire N__52647;
    wire N__52644;
    wire N__52641;
    wire N__52640;
    wire N__52639;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52628;
    wire N__52627;
    wire N__52626;
    wire N__52623;
    wire N__52620;
    wire N__52617;
    wire N__52614;
    wire N__52611;
    wire N__52610;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52602;
    wire N__52601;
    wire N__52598;
    wire N__52589;
    wire N__52588;
    wire N__52587;
    wire N__52586;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52574;
    wire N__52571;
    wire N__52570;
    wire N__52567;
    wire N__52562;
    wire N__52559;
    wire N__52556;
    wire N__52553;
    wire N__52552;
    wire N__52549;
    wire N__52548;
    wire N__52547;
    wire N__52546;
    wire N__52543;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52531;
    wire N__52528;
    wire N__52523;
    wire N__52518;
    wire N__52515;
    wire N__52512;
    wire N__52509;
    wire N__52506;
    wire N__52503;
    wire N__52502;
    wire N__52499;
    wire N__52498;
    wire N__52495;
    wire N__52490;
    wire N__52487;
    wire N__52482;
    wire N__52473;
    wire N__52468;
    wire N__52465;
    wire N__52462;
    wire N__52459;
    wire N__52452;
    wire N__52449;
    wire N__52442;
    wire N__52437;
    wire N__52428;
    wire N__52425;
    wire N__52422;
    wire N__52419;
    wire N__52416;
    wire N__52413;
    wire N__52412;
    wire N__52411;
    wire N__52410;
    wire N__52409;
    wire N__52408;
    wire N__52407;
    wire N__52406;
    wire N__52405;
    wire N__52404;
    wire N__52401;
    wire N__52398;
    wire N__52395;
    wire N__52392;
    wire N__52389;
    wire N__52388;
    wire N__52387;
    wire N__52386;
    wire N__52383;
    wire N__52374;
    wire N__52371;
    wire N__52370;
    wire N__52367;
    wire N__52362;
    wire N__52359;
    wire N__52356;
    wire N__52355;
    wire N__52354;
    wire N__52351;
    wire N__52348;
    wire N__52347;
    wire N__52346;
    wire N__52345;
    wire N__52344;
    wire N__52339;
    wire N__52336;
    wire N__52333;
    wire N__52332;
    wire N__52331;
    wire N__52330;
    wire N__52321;
    wire N__52316;
    wire N__52311;
    wire N__52302;
    wire N__52299;
    wire N__52294;
    wire N__52287;
    wire N__52284;
    wire N__52269;
    wire N__52266;
    wire N__52265;
    wire N__52262;
    wire N__52259;
    wire N__52258;
    wire N__52255;
    wire N__52254;
    wire N__52251;
    wire N__52248;
    wire N__52245;
    wire N__52244;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52231;
    wire N__52228;
    wire N__52225;
    wire N__52212;
    wire N__52209;
    wire N__52206;
    wire N__52203;
    wire N__52200;
    wire N__52197;
    wire N__52194;
    wire N__52191;
    wire N__52188;
    wire N__52187;
    wire N__52184;
    wire N__52181;
    wire N__52178;
    wire N__52177;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52156;
    wire N__52153;
    wire N__52146;
    wire N__52143;
    wire N__52140;
    wire N__52137;
    wire N__52134;
    wire N__52131;
    wire N__52128;
    wire N__52125;
    wire N__52124;
    wire N__52121;
    wire N__52118;
    wire N__52117;
    wire N__52114;
    wire N__52113;
    wire N__52112;
    wire N__52111;
    wire N__52108;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52092;
    wire N__52087;
    wire N__52084;
    wire N__52079;
    wire N__52076;
    wire N__52073;
    wire N__52066;
    wire N__52063;
    wire N__52060;
    wire N__52059;
    wire N__52058;
    wire N__52055;
    wire N__52052;
    wire N__52049;
    wire N__52046;
    wire N__52043;
    wire N__52032;
    wire N__52029;
    wire N__52028;
    wire N__52027;
    wire N__52026;
    wire N__52023;
    wire N__52022;
    wire N__52021;
    wire N__52020;
    wire N__52019;
    wire N__52018;
    wire N__52017;
    wire N__52016;
    wire N__52015;
    wire N__52014;
    wire N__52013;
    wire N__52012;
    wire N__52011;
    wire N__52010;
    wire N__52009;
    wire N__52008;
    wire N__52007;
    wire N__52004;
    wire N__52001;
    wire N__52000;
    wire N__51999;
    wire N__51998;
    wire N__51997;
    wire N__51996;
    wire N__51995;
    wire N__51994;
    wire N__51993;
    wire N__51992;
    wire N__51989;
    wire N__51986;
    wire N__51983;
    wire N__51978;
    wire N__51961;
    wire N__51960;
    wire N__51959;
    wire N__51958;
    wire N__51951;
    wire N__51950;
    wire N__51949;
    wire N__51948;
    wire N__51947;
    wire N__51946;
    wire N__51945;
    wire N__51944;
    wire N__51943;
    wire N__51940;
    wire N__51937;
    wire N__51932;
    wire N__51929;
    wire N__51926;
    wire N__51925;
    wire N__51924;
    wire N__51921;
    wire N__51918;
    wire N__51917;
    wire N__51916;
    wire N__51913;
    wire N__51910;
    wire N__51909;
    wire N__51906;
    wire N__51905;
    wire N__51904;
    wire N__51901;
    wire N__51898;
    wire N__51887;
    wire N__51884;
    wire N__51881;
    wire N__51880;
    wire N__51879;
    wire N__51878;
    wire N__51877;
    wire N__51876;
    wire N__51873;
    wire N__51872;
    wire N__51871;
    wire N__51870;
    wire N__51869;
    wire N__51868;
    wire N__51867;
    wire N__51866;
    wire N__51865;
    wire N__51864;
    wire N__51863;
    wire N__51862;
    wire N__51861;
    wire N__51860;
    wire N__51859;
    wire N__51858;
    wire N__51855;
    wire N__51838;
    wire N__51827;
    wire N__51826;
    wire N__51825;
    wire N__51824;
    wire N__51821;
    wire N__51818;
    wire N__51813;
    wire N__51808;
    wire N__51801;
    wire N__51800;
    wire N__51799;
    wire N__51796;
    wire N__51793;
    wire N__51792;
    wire N__51789;
    wire N__51778;
    wire N__51775;
    wire N__51772;
    wire N__51769;
    wire N__51762;
    wire N__51761;
    wire N__51760;
    wire N__51759;
    wire N__51758;
    wire N__51755;
    wire N__51740;
    wire N__51731;
    wire N__51728;
    wire N__51727;
    wire N__51726;
    wire N__51725;
    wire N__51724;
    wire N__51723;
    wire N__51722;
    wire N__51721;
    wire N__51720;
    wire N__51719;
    wire N__51718;
    wire N__51715;
    wire N__51714;
    wire N__51711;
    wire N__51708;
    wire N__51703;
    wire N__51696;
    wire N__51685;
    wire N__51682;
    wire N__51679;
    wire N__51674;
    wire N__51671;
    wire N__51666;
    wire N__51657;
    wire N__51656;
    wire N__51655;
    wire N__51654;
    wire N__51653;
    wire N__51652;
    wire N__51651;
    wire N__51650;
    wire N__51649;
    wire N__51646;
    wire N__51645;
    wire N__51644;
    wire N__51643;
    wire N__51642;
    wire N__51641;
    wire N__51638;
    wire N__51637;
    wire N__51636;
    wire N__51633;
    wire N__51632;
    wire N__51629;
    wire N__51626;
    wire N__51623;
    wire N__51620;
    wire N__51617;
    wire N__51614;
    wire N__51611;
    wire N__51604;
    wire N__51599;
    wire N__51596;
    wire N__51587;
    wire N__51578;
    wire N__51575;
    wire N__51574;
    wire N__51573;
    wire N__51572;
    wire N__51569;
    wire N__51566;
    wire N__51563;
    wire N__51556;
    wire N__51539;
    wire N__51536;
    wire N__51533;
    wire N__51526;
    wire N__51519;
    wire N__51512;
    wire N__51503;
    wire N__51496;
    wire N__51491;
    wire N__51486;
    wire N__51481;
    wire N__51474;
    wire N__51465;
    wire N__51438;
    wire N__51437;
    wire N__51436;
    wire N__51435;
    wire N__51432;
    wire N__51429;
    wire N__51428;
    wire N__51425;
    wire N__51422;
    wire N__51419;
    wire N__51416;
    wire N__51413;
    wire N__51410;
    wire N__51407;
    wire N__51400;
    wire N__51397;
    wire N__51394;
    wire N__51389;
    wire N__51384;
    wire N__51383;
    wire N__51382;
    wire N__51381;
    wire N__51378;
    wire N__51375;
    wire N__51374;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51358;
    wire N__51357;
    wire N__51356;
    wire N__51353;
    wire N__51350;
    wire N__51347;
    wire N__51342;
    wire N__51339;
    wire N__51336;
    wire N__51333;
    wire N__51330;
    wire N__51327;
    wire N__51324;
    wire N__51321;
    wire N__51306;
    wire N__51303;
    wire N__51302;
    wire N__51301;
    wire N__51300;
    wire N__51299;
    wire N__51296;
    wire N__51293;
    wire N__51290;
    wire N__51287;
    wire N__51284;
    wire N__51283;
    wire N__51278;
    wire N__51277;
    wire N__51270;
    wire N__51267;
    wire N__51264;
    wire N__51261;
    wire N__51258;
    wire N__51257;
    wire N__51250;
    wire N__51247;
    wire N__51244;
    wire N__51241;
    wire N__51238;
    wire N__51233;
    wire N__51228;
    wire N__51225;
    wire N__51222;
    wire N__51219;
    wire N__51216;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51204;
    wire N__51201;
    wire N__51198;
    wire N__51195;
    wire N__51194;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51182;
    wire N__51177;
    wire N__51176;
    wire N__51173;
    wire N__51170;
    wire N__51167;
    wire N__51164;
    wire N__51161;
    wire N__51156;
    wire N__51155;
    wire N__51152;
    wire N__51151;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51120;
    wire N__51117;
    wire N__51114;
    wire N__51111;
    wire N__51110;
    wire N__51109;
    wire N__51108;
    wire N__51107;
    wire N__51106;
    wire N__51103;
    wire N__51100;
    wire N__51097;
    wire N__51094;
    wire N__51091;
    wire N__51088;
    wire N__51083;
    wire N__51078;
    wire N__51075;
    wire N__51072;
    wire N__51071;
    wire N__51068;
    wire N__51065;
    wire N__51062;
    wire N__51059;
    wire N__51056;
    wire N__51055;
    wire N__51054;
    wire N__51049;
    wire N__51046;
    wire N__51041;
    wire N__51038;
    wire N__51035;
    wire N__51024;
    wire N__51021;
    wire N__51020;
    wire N__51019;
    wire N__51016;
    wire N__51013;
    wire N__51012;
    wire N__51009;
    wire N__51006;
    wire N__51003;
    wire N__51000;
    wire N__50999;
    wire N__50996;
    wire N__50993;
    wire N__50990;
    wire N__50987;
    wire N__50984;
    wire N__50981;
    wire N__50978;
    wire N__50973;
    wire N__50970;
    wire N__50967;
    wire N__50962;
    wire N__50959;
    wire N__50956;
    wire N__50949;
    wire N__50946;
    wire N__50943;
    wire N__50940;
    wire N__50939;
    wire N__50936;
    wire N__50933;
    wire N__50930;
    wire N__50927;
    wire N__50922;
    wire N__50921;
    wire N__50920;
    wire N__50917;
    wire N__50914;
    wire N__50911;
    wire N__50908;
    wire N__50905;
    wire N__50902;
    wire N__50899;
    wire N__50896;
    wire N__50889;
    wire N__50886;
    wire N__50883;
    wire N__50882;
    wire N__50879;
    wire N__50876;
    wire N__50873;
    wire N__50870;
    wire N__50867;
    wire N__50862;
    wire N__50861;
    wire N__50858;
    wire N__50855;
    wire N__50854;
    wire N__50851;
    wire N__50848;
    wire N__50845;
    wire N__50840;
    wire N__50835;
    wire N__50832;
    wire N__50829;
    wire N__50826;
    wire N__50823;
    wire N__50820;
    wire N__50817;
    wire N__50814;
    wire N__50811;
    wire N__50808;
    wire N__50807;
    wire N__50802;
    wire N__50799;
    wire N__50798;
    wire N__50797;
    wire N__50796;
    wire N__50795;
    wire N__50794;
    wire N__50793;
    wire N__50792;
    wire N__50791;
    wire N__50790;
    wire N__50787;
    wire N__50786;
    wire N__50783;
    wire N__50782;
    wire N__50781;
    wire N__50780;
    wire N__50779;
    wire N__50778;
    wire N__50777;
    wire N__50768;
    wire N__50761;
    wire N__50758;
    wire N__50757;
    wire N__50756;
    wire N__50755;
    wire N__50754;
    wire N__50753;
    wire N__50752;
    wire N__50751;
    wire N__50748;
    wire N__50743;
    wire N__50740;
    wire N__50737;
    wire N__50734;
    wire N__50733;
    wire N__50732;
    wire N__50731;
    wire N__50730;
    wire N__50729;
    wire N__50726;
    wire N__50721;
    wire N__50714;
    wire N__50705;
    wire N__50702;
    wire N__50697;
    wire N__50694;
    wire N__50689;
    wire N__50688;
    wire N__50681;
    wire N__50672;
    wire N__50671;
    wire N__50670;
    wire N__50669;
    wire N__50668;
    wire N__50659;
    wire N__50658;
    wire N__50657;
    wire N__50654;
    wire N__50647;
    wire N__50644;
    wire N__50639;
    wire N__50630;
    wire N__50627;
    wire N__50622;
    wire N__50617;
    wire N__50604;
    wire N__50603;
    wire N__50602;
    wire N__50601;
    wire N__50600;
    wire N__50599;
    wire N__50598;
    wire N__50597;
    wire N__50596;
    wire N__50595;
    wire N__50594;
    wire N__50593;
    wire N__50588;
    wire N__50585;
    wire N__50584;
    wire N__50581;
    wire N__50580;
    wire N__50579;
    wire N__50578;
    wire N__50573;
    wire N__50572;
    wire N__50571;
    wire N__50566;
    wire N__50557;
    wire N__50552;
    wire N__50549;
    wire N__50546;
    wire N__50543;
    wire N__50540;
    wire N__50539;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50527;
    wire N__50522;
    wire N__50515;
    wire N__50510;
    wire N__50505;
    wire N__50498;
    wire N__50495;
    wire N__50490;
    wire N__50481;
    wire N__50478;
    wire N__50477;
    wire N__50474;
    wire N__50471;
    wire N__50468;
    wire N__50465;
    wire N__50462;
    wire N__50457;
    wire N__50454;
    wire N__50453;
    wire N__50452;
    wire N__50449;
    wire N__50446;
    wire N__50443;
    wire N__50440;
    wire N__50433;
    wire N__50430;
    wire N__50427;
    wire N__50424;
    wire N__50421;
    wire N__50418;
    wire N__50415;
    wire N__50412;
    wire N__50411;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50405;
    wire N__50402;
    wire N__50399;
    wire N__50396;
    wire N__50393;
    wire N__50390;
    wire N__50389;
    wire N__50384;
    wire N__50381;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50366;
    wire N__50363;
    wire N__50358;
    wire N__50355;
    wire N__50350;
    wire N__50349;
    wire N__50346;
    wire N__50343;
    wire N__50340;
    wire N__50337;
    wire N__50328;
    wire N__50325;
    wire N__50322;
    wire N__50321;
    wire N__50320;
    wire N__50319;
    wire N__50318;
    wire N__50315;
    wire N__50312;
    wire N__50309;
    wire N__50306;
    wire N__50303;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50272;
    wire N__50267;
    wire N__50264;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50238;
    wire N__50235;
    wire N__50232;
    wire N__50231;
    wire N__50228;
    wire N__50225;
    wire N__50220;
    wire N__50217;
    wire N__50216;
    wire N__50213;
    wire N__50210;
    wire N__50205;
    wire N__50202;
    wire N__50201;
    wire N__50198;
    wire N__50195;
    wire N__50192;
    wire N__50187;
    wire N__50184;
    wire N__50181;
    wire N__50178;
    wire N__50177;
    wire N__50174;
    wire N__50171;
    wire N__50168;
    wire N__50165;
    wire N__50160;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50148;
    wire N__50145;
    wire N__50142;
    wire N__50141;
    wire N__50138;
    wire N__50135;
    wire N__50132;
    wire N__50129;
    wire N__50124;
    wire N__50121;
    wire N__50118;
    wire N__50117;
    wire N__50114;
    wire N__50113;
    wire N__50110;
    wire N__50107;
    wire N__50104;
    wire N__50101;
    wire N__50098;
    wire N__50095;
    wire N__50088;
    wire N__50087;
    wire N__50084;
    wire N__50081;
    wire N__50080;
    wire N__50077;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50065;
    wire N__50058;
    wire N__50055;
    wire N__50052;
    wire N__50051;
    wire N__50048;
    wire N__50047;
    wire N__50046;
    wire N__50045;
    wire N__50042;
    wire N__50039;
    wire N__50038;
    wire N__50037;
    wire N__50036;
    wire N__50035;
    wire N__50032;
    wire N__50031;
    wire N__50030;
    wire N__50027;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50014;
    wire N__50013;
    wire N__50012;
    wire N__50009;
    wire N__50008;
    wire N__50001;
    wire N__49998;
    wire N__49995;
    wire N__49994;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49984;
    wire N__49981;
    wire N__49976;
    wire N__49973;
    wire N__49966;
    wire N__49965;
    wire N__49964;
    wire N__49961;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49941;
    wire N__49936;
    wire N__49933;
    wire N__49928;
    wire N__49921;
    wire N__49918;
    wire N__49913;
    wire N__49908;
    wire N__49905;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49886;
    wire N__49881;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49873;
    wire N__49872;
    wire N__49871;
    wire N__49868;
    wire N__49867;
    wire N__49864;
    wire N__49859;
    wire N__49850;
    wire N__49849;
    wire N__49848;
    wire N__49847;
    wire N__49846;
    wire N__49843;
    wire N__49840;
    wire N__49837;
    wire N__49832;
    wire N__49829;
    wire N__49826;
    wire N__49823;
    wire N__49820;
    wire N__49813;
    wire N__49800;
    wire N__49797;
    wire N__49794;
    wire N__49793;
    wire N__49790;
    wire N__49787;
    wire N__49786;
    wire N__49781;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49761;
    wire N__49756;
    wire N__49749;
    wire N__49748;
    wire N__49745;
    wire N__49742;
    wire N__49737;
    wire N__49734;
    wire N__49733;
    wire N__49732;
    wire N__49731;
    wire N__49728;
    wire N__49723;
    wire N__49720;
    wire N__49713;
    wire N__49712;
    wire N__49709;
    wire N__49706;
    wire N__49701;
    wire N__49700;
    wire N__49697;
    wire N__49696;
    wire N__49695;
    wire N__49692;
    wire N__49689;
    wire N__49686;
    wire N__49683;
    wire N__49674;
    wire N__49671;
    wire N__49668;
    wire N__49665;
    wire N__49662;
    wire N__49659;
    wire N__49656;
    wire N__49655;
    wire N__49654;
    wire N__49653;
    wire N__49650;
    wire N__49643;
    wire N__49640;
    wire N__49637;
    wire N__49634;
    wire N__49629;
    wire N__49626;
    wire N__49623;
    wire N__49620;
    wire N__49619;
    wire N__49616;
    wire N__49613;
    wire N__49610;
    wire N__49605;
    wire N__49602;
    wire N__49601;
    wire N__49598;
    wire N__49595;
    wire N__49592;
    wire N__49591;
    wire N__49590;
    wire N__49589;
    wire N__49588;
    wire N__49587;
    wire N__49586;
    wire N__49585;
    wire N__49582;
    wire N__49579;
    wire N__49576;
    wire N__49575;
    wire N__49574;
    wire N__49567;
    wire N__49566;
    wire N__49563;
    wire N__49562;
    wire N__49559;
    wire N__49556;
    wire N__49553;
    wire N__49550;
    wire N__49543;
    wire N__49540;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49526;
    wire N__49519;
    wire N__49512;
    wire N__49503;
    wire N__49500;
    wire N__49499;
    wire N__49498;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49493;
    wire N__49492;
    wire N__49491;
    wire N__49490;
    wire N__49489;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49485;
    wire N__49484;
    wire N__49483;
    wire N__49482;
    wire N__49481;
    wire N__49478;
    wire N__49471;
    wire N__49468;
    wire N__49465;
    wire N__49464;
    wire N__49463;
    wire N__49460;
    wire N__49457;
    wire N__49454;
    wire N__49449;
    wire N__49446;
    wire N__49439;
    wire N__49430;
    wire N__49427;
    wire N__49426;
    wire N__49425;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49409;
    wire N__49408;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49404;
    wire N__49403;
    wire N__49402;
    wire N__49401;
    wire N__49394;
    wire N__49391;
    wire N__49388;
    wire N__49385;
    wire N__49380;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49362;
    wire N__49353;
    wire N__49348;
    wire N__49339;
    wire N__49332;
    wire N__49327;
    wire N__49324;
    wire N__49317;
    wire N__49310;
    wire N__49293;
    wire N__49292;
    wire N__49289;
    wire N__49286;
    wire N__49281;
    wire N__49280;
    wire N__49279;
    wire N__49272;
    wire N__49271;
    wire N__49268;
    wire N__49265;
    wire N__49262;
    wire N__49259;
    wire N__49254;
    wire N__49251;
    wire N__49248;
    wire N__49245;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49230;
    wire N__49227;
    wire N__49224;
    wire N__49221;
    wire N__49218;
    wire N__49215;
    wire N__49212;
    wire N__49211;
    wire N__49208;
    wire N__49205;
    wire N__49202;
    wire N__49197;
    wire N__49196;
    wire N__49193;
    wire N__49190;
    wire N__49187;
    wire N__49184;
    wire N__49181;
    wire N__49176;
    wire N__49173;
    wire N__49172;
    wire N__49171;
    wire N__49168;
    wire N__49167;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49143;
    wire N__49140;
    wire N__49137;
    wire N__49134;
    wire N__49131;
    wire N__49128;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49104;
    wire N__49101;
    wire N__49098;
    wire N__49095;
    wire N__49092;
    wire N__49089;
    wire N__49088;
    wire N__49087;
    wire N__49086;
    wire N__49083;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49071;
    wire N__49068;
    wire N__49063;
    wire N__49058;
    wire N__49055;
    wire N__49050;
    wire N__49047;
    wire N__49044;
    wire N__49041;
    wire N__49038;
    wire N__49035;
    wire N__49032;
    wire N__49029;
    wire N__49026;
    wire N__49023;
    wire N__49020;
    wire N__49017;
    wire N__49014;
    wire N__49011;
    wire N__49008;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__48998;
    wire N__48993;
    wire N__48990;
    wire N__48989;
    wire N__48986;
    wire N__48983;
    wire N__48978;
    wire N__48975;
    wire N__48974;
    wire N__48971;
    wire N__48968;
    wire N__48965;
    wire N__48962;
    wire N__48957;
    wire N__48954;
    wire N__48953;
    wire N__48950;
    wire N__48947;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48935;
    wire N__48932;
    wire N__48929;
    wire N__48924;
    wire N__48921;
    wire N__48920;
    wire N__48917;
    wire N__48914;
    wire N__48909;
    wire N__48906;
    wire N__48903;
    wire N__48902;
    wire N__48899;
    wire N__48896;
    wire N__48891;
    wire N__48888;
    wire N__48887;
    wire N__48884;
    wire N__48881;
    wire N__48876;
    wire N__48873;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48869;
    wire N__48868;
    wire N__48867;
    wire N__48866;
    wire N__48865;
    wire N__48864;
    wire N__48863;
    wire N__48862;
    wire N__48859;
    wire N__48856;
    wire N__48855;
    wire N__48854;
    wire N__48853;
    wire N__48852;
    wire N__48851;
    wire N__48848;
    wire N__48847;
    wire N__48846;
    wire N__48845;
    wire N__48844;
    wire N__48843;
    wire N__48840;
    wire N__48837;
    wire N__48836;
    wire N__48835;
    wire N__48834;
    wire N__48833;
    wire N__48832;
    wire N__48817;
    wire N__48806;
    wire N__48805;
    wire N__48804;
    wire N__48801;
    wire N__48800;
    wire N__48799;
    wire N__48798;
    wire N__48797;
    wire N__48796;
    wire N__48793;
    wire N__48792;
    wire N__48787;
    wire N__48786;
    wire N__48785;
    wire N__48784;
    wire N__48779;
    wire N__48778;
    wire N__48775;
    wire N__48774;
    wire N__48773;
    wire N__48772;
    wire N__48769;
    wire N__48764;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48758;
    wire N__48755;
    wire N__48754;
    wire N__48747;
    wire N__48742;
    wire N__48735;
    wire N__48728;
    wire N__48721;
    wire N__48718;
    wire N__48715;
    wire N__48710;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48696;
    wire N__48693;
    wire N__48690;
    wire N__48689;
    wire N__48684;
    wire N__48681;
    wire N__48678;
    wire N__48675;
    wire N__48668;
    wire N__48657;
    wire N__48654;
    wire N__48651;
    wire N__48648;
    wire N__48645;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48629;
    wire N__48626;
    wire N__48613;
    wire N__48608;
    wire N__48591;
    wire N__48590;
    wire N__48589;
    wire N__48588;
    wire N__48587;
    wire N__48586;
    wire N__48585;
    wire N__48584;
    wire N__48583;
    wire N__48582;
    wire N__48581;
    wire N__48580;
    wire N__48579;
    wire N__48578;
    wire N__48577;
    wire N__48576;
    wire N__48575;
    wire N__48570;
    wire N__48569;
    wire N__48568;
    wire N__48567;
    wire N__48566;
    wire N__48565;
    wire N__48564;
    wire N__48563;
    wire N__48562;
    wire N__48561;
    wire N__48560;
    wire N__48559;
    wire N__48558;
    wire N__48557;
    wire N__48556;
    wire N__48539;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48531;
    wire N__48530;
    wire N__48529;
    wire N__48528;
    wire N__48517;
    wire N__48514;
    wire N__48509;
    wire N__48502;
    wire N__48497;
    wire N__48482;
    wire N__48481;
    wire N__48480;
    wire N__48479;
    wire N__48476;
    wire N__48473;
    wire N__48470;
    wire N__48467;
    wire N__48466;
    wire N__48465;
    wire N__48464;
    wire N__48461;
    wire N__48458;
    wire N__48457;
    wire N__48456;
    wire N__48455;
    wire N__48452;
    wire N__48449;
    wire N__48444;
    wire N__48441;
    wire N__48434;
    wire N__48431;
    wire N__48426;
    wire N__48419;
    wire N__48416;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48393;
    wire N__48384;
    wire N__48371;
    wire N__48360;
    wire N__48357;
    wire N__48356;
    wire N__48355;
    wire N__48354;
    wire N__48351;
    wire N__48350;
    wire N__48349;
    wire N__48348;
    wire N__48347;
    wire N__48346;
    wire N__48345;
    wire N__48340;
    wire N__48339;
    wire N__48338;
    wire N__48331;
    wire N__48328;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48314;
    wire N__48309;
    wire N__48306;
    wire N__48301;
    wire N__48300;
    wire N__48299;
    wire N__48298;
    wire N__48297;
    wire N__48292;
    wire N__48289;
    wire N__48288;
    wire N__48287;
    wire N__48280;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48276;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48263;
    wire N__48258;
    wire N__48253;
    wire N__48250;
    wire N__48245;
    wire N__48238;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48206;
    wire N__48203;
    wire N__48200;
    wire N__48195;
    wire N__48192;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48180;
    wire N__48177;
    wire N__48174;
    wire N__48173;
    wire N__48170;
    wire N__48167;
    wire N__48162;
    wire N__48159;
    wire N__48158;
    wire N__48155;
    wire N__48152;
    wire N__48147;
    wire N__48144;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48128;
    wire N__48123;
    wire N__48120;
    wire N__48119;
    wire N__48116;
    wire N__48113;
    wire N__48110;
    wire N__48105;
    wire N__48102;
    wire N__48099;
    wire N__48098;
    wire N__48095;
    wire N__48092;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48080;
    wire N__48077;
    wire N__48074;
    wire N__48069;
    wire N__48068;
    wire N__48067;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48048;
    wire N__48045;
    wire N__48042;
    wire N__48035;
    wire N__48030;
    wire N__48027;
    wire N__48026;
    wire N__48025;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48013;
    wire N__48012;
    wire N__48011;
    wire N__48010;
    wire N__48009;
    wire N__48006;
    wire N__48001;
    wire N__47998;
    wire N__47997;
    wire N__47996;
    wire N__47995;
    wire N__47992;
    wire N__47987;
    wire N__47986;
    wire N__47981;
    wire N__47978;
    wire N__47975;
    wire N__47970;
    wire N__47969;
    wire N__47968;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47951;
    wire N__47948;
    wire N__47941;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47915;
    wire N__47914;
    wire N__47911;
    wire N__47906;
    wire N__47901;
    wire N__47898;
    wire N__47897;
    wire N__47896;
    wire N__47895;
    wire N__47892;
    wire N__47891;
    wire N__47888;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47878;
    wire N__47875;
    wire N__47872;
    wire N__47869;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47839;
    wire N__47832;
    wire N__47829;
    wire N__47828;
    wire N__47825;
    wire N__47822;
    wire N__47819;
    wire N__47816;
    wire N__47813;
    wire N__47810;
    wire N__47805;
    wire N__47802;
    wire N__47801;
    wire N__47798;
    wire N__47795;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47784;
    wire N__47783;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47764;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47740;
    wire N__47737;
    wire N__47732;
    wire N__47727;
    wire N__47724;
    wire N__47723;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47713;
    wire N__47706;
    wire N__47703;
    wire N__47702;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47691;
    wire N__47690;
    wire N__47689;
    wire N__47684;
    wire N__47683;
    wire N__47682;
    wire N__47681;
    wire N__47680;
    wire N__47677;
    wire N__47674;
    wire N__47669;
    wire N__47666;
    wire N__47663;
    wire N__47656;
    wire N__47651;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47633;
    wire N__47630;
    wire N__47627;
    wire N__47622;
    wire N__47621;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47604;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47586;
    wire N__47583;
    wire N__47580;
    wire N__47577;
    wire N__47574;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47564;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47552;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47522;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47492;
    wire N__47491;
    wire N__47490;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47480;
    wire N__47477;
    wire N__47474;
    wire N__47473;
    wire N__47470;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47456;
    wire N__47453;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47427;
    wire N__47426;
    wire N__47419;
    wire N__47416;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47398;
    wire N__47395;
    wire N__47388;
    wire N__47385;
    wire N__47384;
    wire N__47383;
    wire N__47378;
    wire N__47377;
    wire N__47374;
    wire N__47371;
    wire N__47368;
    wire N__47367;
    wire N__47366;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47361;
    wire N__47360;
    wire N__47359;
    wire N__47358;
    wire N__47357;
    wire N__47352;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47344;
    wire N__47341;
    wire N__47336;
    wire N__47335;
    wire N__47334;
    wire N__47333;
    wire N__47332;
    wire N__47329;
    wire N__47322;
    wire N__47317;
    wire N__47314;
    wire N__47309;
    wire N__47304;
    wire N__47297;
    wire N__47290;
    wire N__47287;
    wire N__47284;
    wire N__47279;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47243;
    wire N__47240;
    wire N__47237;
    wire N__47236;
    wire N__47233;
    wire N__47232;
    wire N__47231;
    wire N__47228;
    wire N__47225;
    wire N__47224;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47214;
    wire N__47209;
    wire N__47206;
    wire N__47203;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47179;
    wire N__47176;
    wire N__47175;
    wire N__47174;
    wire N__47171;
    wire N__47166;
    wire N__47163;
    wire N__47160;
    wire N__47151;
    wire N__47148;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47135;
    wire N__47132;
    wire N__47127;
    wire N__47124;
    wire N__47123;
    wire N__47122;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47096;
    wire N__47093;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47083;
    wire N__47080;
    wire N__47077;
    wire N__47074;
    wire N__47071;
    wire N__47068;
    wire N__47063;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47032;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46997;
    wire N__46994;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46982;
    wire N__46977;
    wire N__46976;
    wire N__46973;
    wire N__46972;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46956;
    wire N__46953;
    wire N__46952;
    wire N__46949;
    wire N__46946;
    wire N__46945;
    wire N__46942;
    wire N__46939;
    wire N__46936;
    wire N__46933;
    wire N__46930;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46912;
    wire N__46909;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46882;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46868;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46838;
    wire N__46837;
    wire N__46834;
    wire N__46829;
    wire N__46824;
    wire N__46821;
    wire N__46818;
    wire N__46817;
    wire N__46814;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46802;
    wire N__46797;
    wire N__46794;
    wire N__46791;
    wire N__46788;
    wire N__46787;
    wire N__46786;
    wire N__46783;
    wire N__46780;
    wire N__46777;
    wire N__46776;
    wire N__46773;
    wire N__46772;
    wire N__46769;
    wire N__46766;
    wire N__46763;
    wire N__46762;
    wire N__46759;
    wire N__46756;
    wire N__46755;
    wire N__46748;
    wire N__46745;
    wire N__46740;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46730;
    wire N__46727;
    wire N__46724;
    wire N__46719;
    wire N__46716;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46700;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46665;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46655;
    wire N__46652;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46633;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46607;
    wire N__46604;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46580;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46557;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46535;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46515;
    wire N__46512;
    wire N__46511;
    wire N__46508;
    wire N__46507;
    wire N__46504;
    wire N__46501;
    wire N__46498;
    wire N__46495;
    wire N__46492;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46476;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46463;
    wire N__46462;
    wire N__46461;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46449;
    wire N__46448;
    wire N__46447;
    wire N__46446;
    wire N__46443;
    wire N__46436;
    wire N__46433;
    wire N__46430;
    wire N__46427;
    wire N__46424;
    wire N__46421;
    wire N__46418;
    wire N__46413;
    wire N__46406;
    wire N__46405;
    wire N__46404;
    wire N__46401;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46374;
    wire N__46371;
    wire N__46368;
    wire N__46365;
    wire N__46364;
    wire N__46361;
    wire N__46358;
    wire N__46353;
    wire N__46350;
    wire N__46349;
    wire N__46346;
    wire N__46343;
    wire N__46342;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46330;
    wire N__46327;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46268;
    wire N__46265;
    wire N__46262;
    wire N__46259;
    wire N__46256;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46240;
    wire N__46235;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46217;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46197;
    wire N__46194;
    wire N__46193;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46173;
    wire N__46170;
    wire N__46169;
    wire N__46168;
    wire N__46167;
    wire N__46166;
    wire N__46165;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46138;
    wire N__46135;
    wire N__46132;
    wire N__46127;
    wire N__46124;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46114;
    wire N__46109;
    wire N__46106;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46082;
    wire N__46081;
    wire N__46080;
    wire N__46079;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46071;
    wire N__46070;
    wire N__46067;
    wire N__46064;
    wire N__46061;
    wire N__46058;
    wire N__46055;
    wire N__46050;
    wire N__46047;
    wire N__46040;
    wire N__46037;
    wire N__46032;
    wire N__46025;
    wire N__46022;
    wire N__46019;
    wire N__46014;
    wire N__46013;
    wire N__46012;
    wire N__46009;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__46001;
    wire N__46000;
    wire N__45999;
    wire N__45998;
    wire N__45995;
    wire N__45992;
    wire N__45987;
    wire N__45984;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45970;
    wire N__45961;
    wire N__45954;
    wire N__45953;
    wire N__45952;
    wire N__45949;
    wire N__45944;
    wire N__45939;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45921;
    wire N__45920;
    wire N__45917;
    wire N__45916;
    wire N__45915;
    wire N__45914;
    wire N__45911;
    wire N__45910;
    wire N__45907;
    wire N__45904;
    wire N__45899;
    wire N__45894;
    wire N__45885;
    wire N__45882;
    wire N__45881;
    wire N__45880;
    wire N__45879;
    wire N__45878;
    wire N__45877;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45865;
    wire N__45862;
    wire N__45861;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45847;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45829;
    wire N__45826;
    wire N__45819;
    wire N__45810;
    wire N__45807;
    wire N__45806;
    wire N__45803;
    wire N__45800;
    wire N__45795;
    wire N__45794;
    wire N__45793;
    wire N__45792;
    wire N__45791;
    wire N__45788;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45775;
    wire N__45772;
    wire N__45769;
    wire N__45768;
    wire N__45765;
    wire N__45760;
    wire N__45757;
    wire N__45754;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45740;
    wire N__45737;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45725;
    wire N__45724;
    wire N__45721;
    wire N__45716;
    wire N__45713;
    wire N__45710;
    wire N__45707;
    wire N__45696;
    wire N__45693;
    wire N__45690;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45669;
    wire N__45666;
    wire N__45663;
    wire N__45660;
    wire N__45657;
    wire N__45654;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45632;
    wire N__45631;
    wire N__45628;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45614;
    wire N__45611;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45543;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45483;
    wire N__45480;
    wire N__45477;
    wire N__45474;
    wire N__45471;
    wire N__45468;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45447;
    wire N__45444;
    wire N__45441;
    wire N__45438;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45426;
    wire N__45423;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45381;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45362;
    wire N__45359;
    wire N__45358;
    wire N__45357;
    wire N__45354;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45340;
    wire N__45339;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45308;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45280;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45261;
    wire N__45260;
    wire N__45259;
    wire N__45256;
    wire N__45253;
    wire N__45250;
    wire N__45243;
    wire N__45240;
    wire N__45237;
    wire N__45236;
    wire N__45235;
    wire N__45234;
    wire N__45233;
    wire N__45230;
    wire N__45227;
    wire N__45226;
    wire N__45223;
    wire N__45220;
    wire N__45217;
    wire N__45212;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45187;
    wire N__45184;
    wire N__45177;
    wire N__45174;
    wire N__45173;
    wire N__45172;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45164;
    wire N__45161;
    wire N__45158;
    wire N__45157;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45092;
    wire N__45089;
    wire N__45086;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45035;
    wire N__45032;
    wire N__45029;
    wire N__45026;
    wire N__45023;
    wire N__45020;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45008;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44996;
    wire N__44993;
    wire N__44990;
    wire N__44987;
    wire N__44984;
    wire N__44979;
    wire N__44978;
    wire N__44977;
    wire N__44976;
    wire N__44975;
    wire N__44972;
    wire N__44971;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44957;
    wire N__44954;
    wire N__44951;
    wire N__44948;
    wire N__44947;
    wire N__44942;
    wire N__44939;
    wire N__44936;
    wire N__44935;
    wire N__44934;
    wire N__44933;
    wire N__44932;
    wire N__44931;
    wire N__44928;
    wire N__44923;
    wire N__44920;
    wire N__44917;
    wire N__44910;
    wire N__44909;
    wire N__44908;
    wire N__44907;
    wire N__44902;
    wire N__44895;
    wire N__44890;
    wire N__44887;
    wire N__44882;
    wire N__44875;
    wire N__44862;
    wire N__44861;
    wire N__44860;
    wire N__44857;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44838;
    wire N__44835;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44821;
    wire N__44820;
    wire N__44819;
    wire N__44816;
    wire N__44813;
    wire N__44810;
    wire N__44807;
    wire N__44804;
    wire N__44793;
    wire N__44792;
    wire N__44789;
    wire N__44788;
    wire N__44787;
    wire N__44786;
    wire N__44783;
    wire N__44780;
    wire N__44779;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44759;
    wire N__44756;
    wire N__44753;
    wire N__44750;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44734;
    wire N__44729;
    wire N__44726;
    wire N__44723;
    wire N__44720;
    wire N__44713;
    wire N__44710;
    wire N__44703;
    wire N__44700;
    wire N__44695;
    wire N__44692;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44678;
    wire N__44675;
    wire N__44672;
    wire N__44669;
    wire N__44668;
    wire N__44665;
    wire N__44662;
    wire N__44659;
    wire N__44656;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44640;
    wire N__44637;
    wire N__44634;
    wire N__44633;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44623;
    wire N__44616;
    wire N__44613;
    wire N__44612;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44592;
    wire N__44589;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44562;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44550;
    wire N__44547;
    wire N__44546;
    wire N__44543;
    wire N__44540;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44528;
    wire N__44525;
    wire N__44522;
    wire N__44517;
    wire N__44516;
    wire N__44513;
    wire N__44510;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44486;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44469;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44457;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44445;
    wire N__44442;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44430;
    wire N__44427;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44330;
    wire N__44329;
    wire N__44328;
    wire N__44327;
    wire N__44326;
    wire N__44325;
    wire N__44324;
    wire N__44323;
    wire N__44322;
    wire N__44321;
    wire N__44318;
    wire N__44317;
    wire N__44316;
    wire N__44311;
    wire N__44308;
    wire N__44303;
    wire N__44300;
    wire N__44299;
    wire N__44298;
    wire N__44297;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44271;
    wire N__44268;
    wire N__44261;
    wire N__44258;
    wire N__44253;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44229;
    wire N__44228;
    wire N__44227;
    wire N__44226;
    wire N__44223;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44204;
    wire N__44201;
    wire N__44198;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44177;
    wire N__44174;
    wire N__44171;
    wire N__44168;
    wire N__44165;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44143;
    wire N__44140;
    wire N__44133;
    wire N__44128;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44108;
    wire N__44105;
    wire N__44104;
    wire N__44101;
    wire N__44098;
    wire N__44095;
    wire N__44092;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44059;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44044;
    wire N__44041;
    wire N__44038;
    wire N__44033;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44017;
    wire N__44014;
    wire N__44011;
    wire N__44008;
    wire N__44001;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43974;
    wire N__43971;
    wire N__43970;
    wire N__43967;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43946;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43910;
    wire N__43907;
    wire N__43906;
    wire N__43905;
    wire N__43904;
    wire N__43901;
    wire N__43898;
    wire N__43895;
    wire N__43890;
    wire N__43881;
    wire N__43878;
    wire N__43877;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43861;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43835;
    wire N__43832;
    wire N__43831;
    wire N__43830;
    wire N__43829;
    wire N__43826;
    wire N__43825;
    wire N__43824;
    wire N__43819;
    wire N__43816;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43808;
    wire N__43805;
    wire N__43802;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43783;
    wire N__43780;
    wire N__43775;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43750;
    wire N__43745;
    wire N__43740;
    wire N__43735;
    wire N__43730;
    wire N__43725;
    wire N__43724;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43700;
    wire N__43699;
    wire N__43698;
    wire N__43695;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43601;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43593;
    wire N__43590;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43569;
    wire N__43568;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43539;
    wire N__43536;
    wire N__43531;
    wire N__43528;
    wire N__43521;
    wire N__43518;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43504;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43487;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43470;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43443;
    wire N__43440;
    wire N__43439;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43392;
    wire N__43391;
    wire N__43388;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43373;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43361;
    wire N__43358;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43334;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43316;
    wire N__43311;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43292;
    wire N__43291;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43283;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43243;
    wire N__43240;
    wire N__43235;
    wire N__43230;
    wire N__43229;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43201;
    wire N__43194;
    wire N__43191;
    wire N__43188;
    wire N__43185;
    wire N__43184;
    wire N__43181;
    wire N__43178;
    wire N__43175;
    wire N__43170;
    wire N__43169;
    wire N__43168;
    wire N__43161;
    wire N__43158;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43127;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43116;
    wire N__43113;
    wire N__43106;
    wire N__43103;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43091;
    wire N__43090;
    wire N__43087;
    wire N__43082;
    wire N__43079;
    wire N__43074;
    wire N__43071;
    wire N__43070;
    wire N__43069;
    wire N__43068;
    wire N__43067;
    wire N__43066;
    wire N__43065;
    wire N__43064;
    wire N__43063;
    wire N__43062;
    wire N__43061;
    wire N__43060;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43052;
    wire N__43051;
    wire N__43050;
    wire N__43049;
    wire N__43048;
    wire N__43047;
    wire N__43046;
    wire N__43045;
    wire N__43044;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43006;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42983;
    wire N__42980;
    wire N__42977;
    wire N__42976;
    wire N__42973;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42958;
    wire N__42957;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42933;
    wire N__42930;
    wire N__42925;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42905;
    wire N__42900;
    wire N__42885;
    wire N__42882;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42815;
    wire N__42814;
    wire N__42811;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42803;
    wire N__42802;
    wire N__42799;
    wire N__42794;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42777;
    wire N__42774;
    wire N__42771;
    wire N__42770;
    wire N__42767;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42735;
    wire N__42734;
    wire N__42729;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42437;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42386;
    wire N__42383;
    wire N__42380;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42308;
    wire N__42305;
    wire N__42302;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42287;
    wire N__42286;
    wire N__42285;
    wire N__42284;
    wire N__42283;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42275;
    wire N__42274;
    wire N__42273;
    wire N__42272;
    wire N__42271;
    wire N__42270;
    wire N__42269;
    wire N__42268;
    wire N__42267;
    wire N__42266;
    wire N__42263;
    wire N__42262;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42201;
    wire N__42198;
    wire N__42197;
    wire N__42196;
    wire N__42191;
    wire N__42190;
    wire N__42189;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42179;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42165;
    wire N__42158;
    wire N__42153;
    wire N__42150;
    wire N__42147;
    wire N__42132;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42124;
    wire N__42121;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42108;
    wire N__42105;
    wire N__42100;
    wire N__42097;
    wire N__42090;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42074;
    wire N__42071;
    wire N__42068;
    wire N__42063;
    wire N__42062;
    wire N__42059;
    wire N__42058;
    wire N__42055;
    wire N__42052;
    wire N__42049;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42035;
    wire N__42032;
    wire N__42029;
    wire N__42024;
    wire N__42023;
    wire N__42020;
    wire N__42017;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41991;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41979;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41969;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41954;
    wire N__41953;
    wire N__41950;
    wire N__41947;
    wire N__41944;
    wire N__41939;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41927;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41911;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41891;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41875;
    wire N__41874;
    wire N__41871;
    wire N__41866;
    wire N__41863;
    wire N__41862;
    wire N__41861;
    wire N__41858;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41789;
    wire N__41786;
    wire N__41783;
    wire N__41778;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41764;
    wire N__41763;
    wire N__41762;
    wire N__41757;
    wire N__41754;
    wire N__41749;
    wire N__41742;
    wire N__41741;
    wire N__41740;
    wire N__41739;
    wire N__41736;
    wire N__41731;
    wire N__41730;
    wire N__41729;
    wire N__41726;
    wire N__41725;
    wire N__41724;
    wire N__41723;
    wire N__41718;
    wire N__41713;
    wire N__41708;
    wire N__41705;
    wire N__41704;
    wire N__41703;
    wire N__41702;
    wire N__41701;
    wire N__41700;
    wire N__41699;
    wire N__41698;
    wire N__41695;
    wire N__41688;
    wire N__41679;
    wire N__41672;
    wire N__41669;
    wire N__41666;
    wire N__41663;
    wire N__41660;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41634;
    wire N__41631;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41617;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41601;
    wire N__41598;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41583;
    wire N__41580;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41570;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41541;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41533;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41503;
    wire N__41496;
    wire N__41495;
    wire N__41494;
    wire N__41493;
    wire N__41492;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41456;
    wire N__41453;
    wire N__41450;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41433;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41417;
    wire N__41412;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41377;
    wire N__41374;
    wire N__41371;
    wire N__41368;
    wire N__41365;
    wire N__41358;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41350;
    wire N__41345;
    wire N__41342;
    wire N__41337;
    wire N__41336;
    wire N__41335;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41327;
    wire N__41324;
    wire N__41323;
    wire N__41320;
    wire N__41317;
    wire N__41312;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41301;
    wire N__41296;
    wire N__41293;
    wire N__41288;
    wire N__41285;
    wire N__41284;
    wire N__41281;
    wire N__41276;
    wire N__41273;
    wire N__41270;
    wire N__41267;
    wire N__41264;
    wire N__41261;
    wire N__41258;
    wire N__41255;
    wire N__41244;
    wire N__41241;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41229;
    wire N__41226;
    wire N__41225;
    wire N__41222;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41175;
    wire N__41172;
    wire N__41171;
    wire N__41168;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41151;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41124;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41100;
    wire N__41099;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41070;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41054;
    wire N__41049;
    wire N__41046;
    wire N__41045;
    wire N__41042;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41025;
    wire N__41022;
    wire N__41021;
    wire N__41020;
    wire N__41017;
    wire N__41012;
    wire N__41007;
    wire N__41004;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40996;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40980;
    wire N__40977;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40969;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40953;
    wire N__40950;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40938;
    wire N__40937;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40898;
    wire N__40895;
    wire N__40892;
    wire N__40891;
    wire N__40890;
    wire N__40889;
    wire N__40886;
    wire N__40885;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40863;
    wire N__40862;
    wire N__40859;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40841;
    wire N__40834;
    wire N__40821;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40782;
    wire N__40781;
    wire N__40778;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40754;
    wire N__40751;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40734;
    wire N__40731;
    wire N__40730;
    wire N__40729;
    wire N__40726;
    wire N__40721;
    wire N__40716;
    wire N__40715;
    wire N__40712;
    wire N__40709;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40696;
    wire N__40691;
    wire N__40688;
    wire N__40685;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40670;
    wire N__40669;
    wire N__40668;
    wire N__40667;
    wire N__40666;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40656;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40638;
    wire N__40637;
    wire N__40636;
    wire N__40635;
    wire N__40632;
    wire N__40631;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40586;
    wire N__40569;
    wire N__40568;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40452;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40434;
    wire N__40433;
    wire N__40430;
    wire N__40429;
    wire N__40426;
    wire N__40423;
    wire N__40420;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40357;
    wire N__40354;
    wire N__40347;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40327;
    wire N__40320;
    wire N__40317;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40241;
    wire N__40238;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40160;
    wire N__40157;
    wire N__40156;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40146;
    wire N__40145;
    wire N__40142;
    wire N__40139;
    wire N__40136;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40122;
    wire N__40121;
    wire N__40120;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40071;
    wire N__40068;
    wire N__40065;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40029;
    wire N__40026;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39787;
    wire N__39784;
    wire N__39781;
    wire N__39778;
    wire N__39773;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39754;
    wire N__39749;
    wire N__39746;
    wire N__39743;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39728;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39659;
    wire N__39658;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39638;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39605;
    wire N__39604;
    wire N__39597;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39476;
    wire N__39475;
    wire N__39472;
    wire N__39467;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39344;
    wire N__39341;
    wire N__39338;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39287;
    wire N__39284;
    wire N__39281;
    wire N__39276;
    wire N__39275;
    wire N__39272;
    wire N__39269;
    wire N__39264;
    wire N__39261;
    wire N__39260;
    wire N__39259;
    wire N__39256;
    wire N__39251;
    wire N__39246;
    wire N__39245;
    wire N__39242;
    wire N__39241;
    wire N__39240;
    wire N__39237;
    wire N__39230;
    wire N__39225;
    wire N__39224;
    wire N__39223;
    wire N__39222;
    wire N__39219;
    wire N__39212;
    wire N__39207;
    wire N__39206;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39147;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39135;
    wire N__39132;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39122;
    wire N__39119;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39095;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39078;
    wire N__39077;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38966;
    wire N__38963;
    wire N__38960;
    wire N__38955;
    wire N__38952;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38813;
    wire N__38810;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38798;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38769;
    wire N__38766;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38755;
    wire N__38754;
    wire N__38753;
    wire N__38752;
    wire N__38751;
    wire N__38750;
    wire N__38749;
    wire N__38748;
    wire N__38747;
    wire N__38746;
    wire N__38745;
    wire N__38742;
    wire N__38741;
    wire N__38740;
    wire N__38739;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38679;
    wire N__38676;
    wire N__38675;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38607;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38595;
    wire N__38592;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38562;
    wire N__38559;
    wire N__38558;
    wire N__38557;
    wire N__38556;
    wire N__38553;
    wire N__38552;
    wire N__38549;
    wire N__38546;
    wire N__38543;
    wire N__38540;
    wire N__38537;
    wire N__38534;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38508;
    wire N__38501;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38482;
    wire N__38481;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38451;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38426;
    wire N__38423;
    wire N__38420;
    wire N__38417;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38393;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38186;
    wire N__38183;
    wire N__38180;
    wire N__38177;
    wire N__38174;
    wire N__38171;
    wire N__38168;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38109;
    wire N__38106;
    wire N__38105;
    wire N__38102;
    wire N__38099;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38075;
    wire N__38070;
    wire N__38069;
    wire N__38066;
    wire N__38063;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37986;
    wire N__37983;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37958;
    wire N__37955;
    wire N__37954;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37923;
    wire N__37920;
    wire N__37919;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37877;
    wire N__37874;
    wire N__37871;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37857;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37805;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37749;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37731;
    wire N__37728;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37698;
    wire N__37695;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37652;
    wire N__37649;
    wire N__37646;
    wire N__37645;
    wire N__37644;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37580;
    wire N__37575;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37500;
    wire N__37497;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37470;
    wire N__37467;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37448;
    wire N__37447;
    wire N__37444;
    wire N__37441;
    wire N__37440;
    wire N__37437;
    wire N__37432;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37413;
    wire N__37410;
    wire N__37405;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37389;
    wire N__37386;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37344;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37332;
    wire N__37329;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37317;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37309;
    wire N__37308;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37300;
    wire N__37299;
    wire N__37298;
    wire N__37297;
    wire N__37294;
    wire N__37293;
    wire N__37292;
    wire N__37291;
    wire N__37288;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37276;
    wire N__37273;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37258;
    wire N__37255;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37235;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37145;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37115;
    wire N__37112;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37085;
    wire N__37082;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37029;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36968;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36920;
    wire N__36919;
    wire N__36914;
    wire N__36913;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36885;
    wire N__36882;
    wire N__36881;
    wire N__36880;
    wire N__36879;
    wire N__36876;
    wire N__36873;
    wire N__36868;
    wire N__36865;
    wire N__36858;
    wire N__36855;
    wire N__36854;
    wire N__36853;
    wire N__36852;
    wire N__36849;
    wire N__36844;
    wire N__36841;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36827;
    wire N__36826;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36741;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36707;
    wire N__36706;
    wire N__36705;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36681;
    wire N__36672;
    wire N__36669;
    wire N__36668;
    wire N__36667;
    wire N__36666;
    wire N__36663;
    wire N__36658;
    wire N__36655;
    wire N__36648;
    wire N__36645;
    wire N__36644;
    wire N__36641;
    wire N__36640;
    wire N__36639;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36624;
    wire N__36615;
    wire N__36612;
    wire N__36611;
    wire N__36610;
    wire N__36605;
    wire N__36604;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36566;
    wire N__36563;
    wire N__36562;
    wire N__36561;
    wire N__36560;
    wire N__36559;
    wire N__36558;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36539;
    wire N__36538;
    wire N__36537;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36496;
    wire N__36487;
    wire N__36480;
    wire N__36477;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36366;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36303;
    wire N__36302;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36287;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36231;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36209;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36195;
    wire N__36192;
    wire N__36189;
    wire N__36186;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36159;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36056;
    wire N__36055;
    wire N__36052;
    wire N__36047;
    wire N__36044;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35894;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35885;
    wire N__35884;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35846;
    wire N__35845;
    wire N__35844;
    wire N__35843;
    wire N__35842;
    wire N__35841;
    wire N__35840;
    wire N__35837;
    wire N__35822;
    wire N__35817;
    wire N__35816;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35808;
    wire N__35807;
    wire N__35806;
    wire N__35805;
    wire N__35804;
    wire N__35803;
    wire N__35802;
    wire N__35799;
    wire N__35798;
    wire N__35797;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35779;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35760;
    wire N__35759;
    wire N__35758;
    wire N__35757;
    wire N__35756;
    wire N__35751;
    wire N__35748;
    wire N__35743;
    wire N__35742;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35719;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35703;
    wire N__35702;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35688;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35668;
    wire N__35663;
    wire N__35660;
    wire N__35653;
    wire N__35646;
    wire N__35637;
    wire N__35636;
    wire N__35635;
    wire N__35634;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35630;
    wire N__35629;
    wire N__35628;
    wire N__35627;
    wire N__35626;
    wire N__35625;
    wire N__35624;
    wire N__35623;
    wire N__35622;
    wire N__35621;
    wire N__35620;
    wire N__35619;
    wire N__35618;
    wire N__35617;
    wire N__35616;
    wire N__35613;
    wire N__35608;
    wire N__35599;
    wire N__35598;
    wire N__35595;
    wire N__35586;
    wire N__35585;
    wire N__35580;
    wire N__35579;
    wire N__35574;
    wire N__35571;
    wire N__35570;
    wire N__35569;
    wire N__35560;
    wire N__35559;
    wire N__35558;
    wire N__35557;
    wire N__35556;
    wire N__35555;
    wire N__35554;
    wire N__35553;
    wire N__35552;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35538;
    wire N__35537;
    wire N__35536;
    wire N__35535;
    wire N__35532;
    wire N__35531;
    wire N__35530;
    wire N__35529;
    wire N__35528;
    wire N__35527;
    wire N__35526;
    wire N__35521;
    wire N__35520;
    wire N__35517;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35496;
    wire N__35495;
    wire N__35494;
    wire N__35493;
    wire N__35492;
    wire N__35487;
    wire N__35478;
    wire N__35473;
    wire N__35470;
    wire N__35465;
    wire N__35460;
    wire N__35459;
    wire N__35458;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35412;
    wire N__35411;
    wire N__35410;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35405;
    wire N__35404;
    wire N__35403;
    wire N__35402;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35394;
    wire N__35383;
    wire N__35380;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35353;
    wire N__35350;
    wire N__35339;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35304;
    wire N__35301;
    wire N__35294;
    wire N__35281;
    wire N__35278;
    wire N__35273;
    wire N__35250;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35233;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35219;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35199;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35177;
    wire N__35176;
    wire N__35173;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35120;
    wire N__35109;
    wire N__35108;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35072;
    wire N__35067;
    wire N__35066;
    wire N__35065;
    wire N__35062;
    wire N__35057;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35045;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35004;
    wire N__35003;
    wire N__34998;
    wire N__34997;
    wire N__34996;
    wire N__34995;
    wire N__34994;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34980;
    wire N__34977;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34941;
    wire N__34938;
    wire N__34937;
    wire N__34934;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34902;
    wire N__34901;
    wire N__34898;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34794;
    wire N__34793;
    wire N__34792;
    wire N__34791;
    wire N__34790;
    wire N__34789;
    wire N__34788;
    wire N__34787;
    wire N__34786;
    wire N__34785;
    wire N__34784;
    wire N__34783;
    wire N__34782;
    wire N__34781;
    wire N__34780;
    wire N__34777;
    wire N__34776;
    wire N__34773;
    wire N__34772;
    wire N__34771;
    wire N__34768;
    wire N__34753;
    wire N__34752;
    wire N__34751;
    wire N__34750;
    wire N__34749;
    wire N__34732;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34711;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34692;
    wire N__34687;
    wire N__34684;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34656;
    wire N__34651;
    wire N__34646;
    wire N__34643;
    wire N__34638;
    wire N__34629;
    wire N__34620;
    wire N__34619;
    wire N__34618;
    wire N__34617;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34602;
    wire N__34601;
    wire N__34600;
    wire N__34599;
    wire N__34598;
    wire N__34597;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34567;
    wire N__34564;
    wire N__34549;
    wire N__34548;
    wire N__34547;
    wire N__34542;
    wire N__34537;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34529;
    wire N__34526;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34492;
    wire N__34489;
    wire N__34484;
    wire N__34477;
    wire N__34464;
    wire N__34463;
    wire N__34460;
    wire N__34459;
    wire N__34458;
    wire N__34457;
    wire N__34454;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34426;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34407;
    wire N__34404;
    wire N__34399;
    wire N__34386;
    wire N__34383;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34285;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34273;
    wire N__34266;
    wire N__34265;
    wire N__34262;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34112;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34094;
    wire N__34089;
    wire N__34088;
    wire N__34087;
    wire N__34084;
    wire N__34079;
    wire N__34074;
    wire N__34073;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34030;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33992;
    wire N__33989;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33972;
    wire N__33969;
    wire N__33968;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33953;
    wire N__33948;
    wire N__33945;
    wire N__33944;
    wire N__33941;
    wire N__33940;
    wire N__33937;
    wire N__33934;
    wire N__33931;
    wire N__33924;
    wire N__33923;
    wire N__33920;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33903;
    wire N__33900;
    wire N__33897;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33884;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33863;
    wire N__33860;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33848;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33833;
    wire N__33828;
    wire N__33825;
    wire N__33822;
    wire N__33821;
    wire N__33820;
    wire N__33817;
    wire N__33812;
    wire N__33807;
    wire N__33806;
    wire N__33803;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33780;
    wire N__33777;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33762;
    wire N__33759;
    wire N__33758;
    wire N__33755;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33738;
    wire N__33735;
    wire N__33734;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33717;
    wire N__33714;
    wire N__33713;
    wire N__33710;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33686;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33677;
    wire N__33676;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33663;
    wire N__33662;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33652;
    wire N__33651;
    wire N__33650;
    wire N__33649;
    wire N__33648;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33621;
    wire N__33620;
    wire N__33615;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33603;
    wire N__33598;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33571;
    wire N__33566;
    wire N__33563;
    wire N__33556;
    wire N__33553;
    wire N__33544;
    wire N__33535;
    wire N__33530;
    wire N__33527;
    wire N__33522;
    wire N__33519;
    wire N__33514;
    wire N__33507;
    wire N__33506;
    wire N__33505;
    wire N__33504;
    wire N__33503;
    wire N__33502;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33494;
    wire N__33493;
    wire N__33492;
    wire N__33491;
    wire N__33490;
    wire N__33489;
    wire N__33488;
    wire N__33487;
    wire N__33486;
    wire N__33485;
    wire N__33484;
    wire N__33483;
    wire N__33482;
    wire N__33481;
    wire N__33480;
    wire N__33479;
    wire N__33478;
    wire N__33477;
    wire N__33476;
    wire N__33475;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33451;
    wire N__33450;
    wire N__33439;
    wire N__33432;
    wire N__33421;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33399;
    wire N__33394;
    wire N__33391;
    wire N__33390;
    wire N__33389;
    wire N__33388;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33378;
    wire N__33377;
    wire N__33376;
    wire N__33375;
    wire N__33374;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33347;
    wire N__33346;
    wire N__33345;
    wire N__33344;
    wire N__33343;
    wire N__33340;
    wire N__33335;
    wire N__33332;
    wire N__33329;
    wire N__33324;
    wire N__33313;
    wire N__33310;
    wire N__33309;
    wire N__33308;
    wire N__33307;
    wire N__33306;
    wire N__33301;
    wire N__33292;
    wire N__33285;
    wire N__33278;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33266;
    wire N__33265;
    wire N__33264;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33254;
    wire N__33251;
    wire N__33246;
    wire N__33245;
    wire N__33234;
    wire N__33227;
    wire N__33222;
    wire N__33221;
    wire N__33220;
    wire N__33219;
    wire N__33218;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33202;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33178;
    wire N__33175;
    wire N__33168;
    wire N__33161;
    wire N__33158;
    wire N__33129;
    wire N__33128;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33116;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33075;
    wire N__33072;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33051;
    wire N__33048;
    wire N__33047;
    wire N__33044;
    wire N__33041;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32847;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32828;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32715;
    wire N__32712;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32697;
    wire N__32694;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32646;
    wire N__32643;
    wire N__32638;
    wire N__32635;
    wire N__32630;
    wire N__32627;
    wire N__32622;
    wire N__32619;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32556;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32499;
    wire N__32496;
    wire N__32495;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32460;
    wire N__32457;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32421;
    wire N__32418;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32360;
    wire N__32359;
    wire N__32356;
    wire N__32351;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32321;
    wire N__32318;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32308;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32274;
    wire N__32273;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32252;
    wire N__32247;
    wire N__32244;
    wire N__32243;
    wire N__32240;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32213;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32207;
    wire N__32206;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32190;
    wire N__32187;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32175;
    wire N__32174;
    wire N__32173;
    wire N__32170;
    wire N__32165;
    wire N__32158;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32134;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32078;
    wire N__32075;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32065;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32036;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31994;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31968;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31943;
    wire N__31938;
    wire N__31937;
    wire N__31934;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31802;
    wire N__31799;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31711;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31692;
    wire N__31691;
    wire N__31690;
    wire N__31689;
    wire N__31688;
    wire N__31687;
    wire N__31686;
    wire N__31685;
    wire N__31684;
    wire N__31683;
    wire N__31678;
    wire N__31673;
    wire N__31672;
    wire N__31671;
    wire N__31670;
    wire N__31669;
    wire N__31668;
    wire N__31661;
    wire N__31660;
    wire N__31659;
    wire N__31658;
    wire N__31657;
    wire N__31656;
    wire N__31655;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31637;
    wire N__31630;
    wire N__31629;
    wire N__31628;
    wire N__31625;
    wire N__31620;
    wire N__31619;
    wire N__31610;
    wire N__31607;
    wire N__31598;
    wire N__31593;
    wire N__31592;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31574;
    wire N__31571;
    wire N__31566;
    wire N__31565;
    wire N__31564;
    wire N__31563;
    wire N__31562;
    wire N__31561;
    wire N__31560;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31542;
    wire N__31537;
    wire N__31530;
    wire N__31515;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31482;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31470;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31458;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31443;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31407;
    wire N__31404;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31386;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31332;
    wire N__31323;
    wire N__31320;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31302;
    wire N__31301;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31249;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31215;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31203;
    wire N__31200;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31188;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31146;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31138;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31117;
    wire N__31114;
    wire N__31107;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31095;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31083;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31068;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31040;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30996;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30942;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30930;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30915;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30903;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30891;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30879;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30864;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30852;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30840;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30830;
    wire N__30825;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30813;
    wire N__30812;
    wire N__30809;
    wire N__30806;
    wire N__30801;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30789;
    wire N__30786;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30750;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30729;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30721;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30713;
    wire N__30710;
    wire N__30709;
    wire N__30708;
    wire N__30707;
    wire N__30706;
    wire N__30703;
    wire N__30702;
    wire N__30701;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30666;
    wire N__30661;
    wire N__30654;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30594;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30582;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30570;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30558;
    wire N__30555;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30527;
    wire N__30526;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30518;
    wire N__30517;
    wire N__30514;
    wire N__30513;
    wire N__30510;
    wire N__30509;
    wire N__30508;
    wire N__30507;
    wire N__30506;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30493;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30476;
    wire N__30473;
    wire N__30472;
    wire N__30469;
    wire N__30468;
    wire N__30467;
    wire N__30460;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30403;
    wire N__30400;
    wire N__30395;
    wire N__30392;
    wire N__30387;
    wire N__30382;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30362;
    wire N__30359;
    wire N__30354;
    wire N__30347;
    wire N__30346;
    wire N__30341;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30321;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30309;
    wire N__30308;
    wire N__30307;
    wire N__30306;
    wire N__30303;
    wire N__30302;
    wire N__30299;
    wire N__30298;
    wire N__30297;
    wire N__30296;
    wire N__30295;
    wire N__30290;
    wire N__30287;
    wire N__30286;
    wire N__30285;
    wire N__30282;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30274;
    wire N__30273;
    wire N__30272;
    wire N__30267;
    wire N__30264;
    wire N__30259;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30226;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30140;
    wire N__30139;
    wire N__30136;
    wire N__30135;
    wire N__30128;
    wire N__30127;
    wire N__30126;
    wire N__30123;
    wire N__30122;
    wire N__30119;
    wire N__30118;
    wire N__30117;
    wire N__30116;
    wire N__30115;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30103;
    wire N__30100;
    wire N__30089;
    wire N__30078;
    wire N__30075;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30051;
    wire N__30050;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30006;
    wire N__30003;
    wire N__30002;
    wire N__30001;
    wire N__30000;
    wire N__29997;
    wire N__29996;
    wire N__29995;
    wire N__29994;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29974;
    wire N__29973;
    wire N__29968;
    wire N__29967;
    wire N__29960;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29916;
    wire N__29913;
    wire N__29912;
    wire N__29911;
    wire N__29910;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29902;
    wire N__29901;
    wire N__29900;
    wire N__29899;
    wire N__29896;
    wire N__29891;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29883;
    wire N__29882;
    wire N__29879;
    wire N__29874;
    wire N__29871;
    wire N__29866;
    wire N__29863;
    wire N__29858;
    wire N__29853;
    wire N__29850;
    wire N__29843;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29798;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29687;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29579;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29468;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29453;
    wire N__29450;
    wire N__29449;
    wire N__29446;
    wire N__29441;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29429;
    wire N__29428;
    wire N__29425;
    wire N__29420;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29293;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29270;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29165;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28898;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28733;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28607;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28457;
    wire N__28456;
    wire N__28455;
    wire N__28448;
    wire N__28445;
    wire N__28440;
    wire N__28439;
    wire N__28438;
    wire N__28435;
    wire N__28430;
    wire N__28427;
    wire N__28422;
    wire N__28419;
    wire N__28418;
    wire N__28417;
    wire N__28416;
    wire N__28415;
    wire N__28406;
    wire N__28403;
    wire N__28398;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28361;
    wire N__28360;
    wire N__28357;
    wire N__28352;
    wire N__28347;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28333;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28314;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28306;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28172;
    wire N__28171;
    wire N__28168;
    wire N__28163;
    wire N__28160;
    wire N__28155;
    wire N__28154;
    wire N__28153;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28139;
    wire N__28138;
    wire N__28135;
    wire N__28128;
    wire N__28125;
    wire N__28124;
    wire N__28123;
    wire N__28122;
    wire N__28119;
    wire N__28118;
    wire N__28117;
    wire N__28116;
    wire N__28115;
    wire N__28114;
    wire N__28113;
    wire N__28112;
    wire N__28109;
    wire N__28108;
    wire N__28105;
    wire N__28104;
    wire N__28103;
    wire N__28100;
    wire N__28099;
    wire N__28098;
    wire N__28097;
    wire N__28094;
    wire N__28093;
    wire N__28092;
    wire N__28091;
    wire N__28088;
    wire N__28083;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28066;
    wire N__28065;
    wire N__28064;
    wire N__28063;
    wire N__28056;
    wire N__28051;
    wire N__28048;
    wire N__28047;
    wire N__28046;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28035;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28009;
    wire N__28006;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27991;
    wire N__27984;
    wire N__27979;
    wire N__27976;
    wire N__27975;
    wire N__27970;
    wire N__27959;
    wire N__27954;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27938;
    wire N__27931;
    wire N__27928;
    wire N__27923;
    wire N__27920;
    wire N__27911;
    wire N__27908;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27887;
    wire N__27886;
    wire N__27883;
    wire N__27878;
    wire N__27875;
    wire N__27870;
    wire N__27867;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27824;
    wire N__27823;
    wire N__27822;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27810;
    wire N__27803;
    wire N__27800;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27758;
    wire N__27757;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27749;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27730;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27709;
    wire N__27708;
    wire N__27707;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27668;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27590;
    wire N__27587;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27551;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27479;
    wire N__27476;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27449;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27441;
    wire N__27440;
    wire N__27439;
    wire N__27438;
    wire N__27435;
    wire N__27434;
    wire N__27433;
    wire N__27432;
    wire N__27431;
    wire N__27430;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27405;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27375;
    wire N__27374;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27348;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27321;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27313;
    wire N__27310;
    wire N__27305;
    wire N__27300;
    wire N__27299;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27295;
    wire N__27294;
    wire N__27291;
    wire N__27284;
    wire N__27281;
    wire N__27276;
    wire N__27273;
    wire N__27268;
    wire N__27265;
    wire N__27264;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27200;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27180;
    wire N__27177;
    wire N__27176;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27102;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27084;
    wire N__27081;
    wire N__27080;
    wire N__27077;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27015;
    wire N__27014;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26885;
    wire N__26880;
    wire N__26879;
    wire N__26876;
    wire N__26871;
    wire N__26868;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26856;
    wire N__26853;
    wire N__26852;
    wire N__26851;
    wire N__26850;
    wire N__26849;
    wire N__26848;
    wire N__26847;
    wire N__26846;
    wire N__26845;
    wire N__26844;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26840;
    wire N__26839;
    wire N__26838;
    wire N__26837;
    wire N__26836;
    wire N__26835;
    wire N__26834;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26830;
    wire N__26829;
    wire N__26826;
    wire N__26821;
    wire N__26820;
    wire N__26819;
    wire N__26816;
    wire N__26815;
    wire N__26798;
    wire N__26789;
    wire N__26786;
    wire N__26785;
    wire N__26784;
    wire N__26783;
    wire N__26782;
    wire N__26779;
    wire N__26778;
    wire N__26773;
    wire N__26768;
    wire N__26767;
    wire N__26766;
    wire N__26765;
    wire N__26764;
    wire N__26763;
    wire N__26762;
    wire N__26761;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26744;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26732;
    wire N__26727;
    wire N__26726;
    wire N__26725;
    wire N__26724;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26700;
    wire N__26693;
    wire N__26686;
    wire N__26681;
    wire N__26674;
    wire N__26669;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26637;
    wire N__26622;
    wire N__26615;
    wire N__26598;
    wire N__26597;
    wire N__26596;
    wire N__26595;
    wire N__26594;
    wire N__26593;
    wire N__26592;
    wire N__26591;
    wire N__26590;
    wire N__26589;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26581;
    wire N__26580;
    wire N__26577;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26565;
    wire N__26562;
    wire N__26561;
    wire N__26560;
    wire N__26559;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26544;
    wire N__26543;
    wire N__26542;
    wire N__26541;
    wire N__26536;
    wire N__26535;
    wire N__26534;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26522;
    wire N__26513;
    wire N__26510;
    wire N__26505;
    wire N__26498;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26482;
    wire N__26479;
    wire N__26470;
    wire N__26463;
    wire N__26448;
    wire N__26447;
    wire N__26444;
    wire N__26443;
    wire N__26442;
    wire N__26441;
    wire N__26438;
    wire N__26437;
    wire N__26436;
    wire N__26435;
    wire N__26434;
    wire N__26433;
    wire N__26432;
    wire N__26431;
    wire N__26428;
    wire N__26427;
    wire N__26426;
    wire N__26425;
    wire N__26422;
    wire N__26421;
    wire N__26420;
    wire N__26419;
    wire N__26416;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26404;
    wire N__26401;
    wire N__26392;
    wire N__26391;
    wire N__26390;
    wire N__26389;
    wire N__26386;
    wire N__26385;
    wire N__26382;
    wire N__26381;
    wire N__26380;
    wire N__26373;
    wire N__26370;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26311;
    wire N__26306;
    wire N__26303;
    wire N__26298;
    wire N__26277;
    wire N__26274;
    wire N__26273;
    wire N__26272;
    wire N__26271;
    wire N__26270;
    wire N__26269;
    wire N__26268;
    wire N__26267;
    wire N__26266;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26262;
    wire N__26261;
    wire N__26260;
    wire N__26259;
    wire N__26258;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26252;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26235;
    wire N__26234;
    wire N__26233;
    wire N__26232;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26214;
    wire N__26207;
    wire N__26206;
    wire N__26205;
    wire N__26204;
    wire N__26203;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26189;
    wire N__26188;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26174;
    wire N__26171;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26151;
    wire N__26134;
    wire N__26131;
    wire N__26126;
    wire N__26119;
    wire N__26112;
    wire N__26101;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26055;
    wire N__26052;
    wire N__26051;
    wire N__26048;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26028;
    wire N__26025;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25940;
    wire N__25937;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25922;
    wire N__25919;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25891;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25752;
    wire N__25751;
    wire N__25750;
    wire N__25749;
    wire N__25748;
    wire N__25747;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25743;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25737;
    wire N__25736;
    wire N__25735;
    wire N__25720;
    wire N__25709;
    wire N__25702;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25688;
    wire N__25687;
    wire N__25686;
    wire N__25685;
    wire N__25684;
    wire N__25683;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25665;
    wire N__25660;
    wire N__25653;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25611;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25599;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25584;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25572;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25560;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25524;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25512;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25497;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25485;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25473;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25461;
    wire N__25458;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25422;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25403;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25352;
    wire N__25351;
    wire N__25348;
    wire N__25343;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25286;
    wire N__25283;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25218;
    wire N__25217;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25205;
    wire N__25202;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25190;
    wire N__25185;
    wire N__25184;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25172;
    wire N__25169;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25131;
    wire N__25128;
    wire N__25127;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25091;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25062;
    wire N__25059;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25041;
    wire N__25038;
    wire N__25037;
    wire N__25036;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24998;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24969;
    wire N__24966;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24948;
    wire N__24947;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24932;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24917;
    wire N__24916;
    wire N__24913;
    wire N__24908;
    wire N__24903;
    wire N__24902;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24879;
    wire N__24878;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24866;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24854;
    wire N__24851;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24834;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24776;
    wire N__24775;
    wire N__24774;
    wire N__24767;
    wire N__24764;
    wire N__24763;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24747;
    wire N__24744;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24696;
    wire N__24693;
    wire N__24692;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24651;
    wire N__24646;
    wire N__24641;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24612;
    wire N__24609;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24573;
    wire N__24570;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24552;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24540;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24528;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24509;
    wire N__24506;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24494;
    wire N__24489;
    wire N__24486;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24453;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24416;
    wire N__24413;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24379;
    wire N__24376;
    wire N__24371;
    wire N__24366;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24354;
    wire N__24351;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24321;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24309;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24297;
    wire N__24294;
    wire N__24293;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24270;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24258;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24246;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24234;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24212;
    wire N__24207;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24192;
    wire N__24189;
    wire N__24186;
    wire N__24185;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24162;
    wire N__24161;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24135;
    wire N__24132;
    wire N__24131;
    wire N__24128;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24108;
    wire N__24107;
    wire N__24106;
    wire N__24101;
    wire N__24098;
    wire N__24093;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24081;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24063;
    wire N__24062;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24039;
    wire N__24038;
    wire N__24037;
    wire N__24034;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24012;
    wire N__24011;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23988;
    wire N__23987;
    wire N__23984;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23964;
    wire N__23961;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23949;
    wire N__23948;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23925;
    wire N__23922;
    wire N__23921;
    wire N__23918;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23903;
    wire N__23900;
    wire N__23895;
    wire N__23894;
    wire N__23893;
    wire N__23892;
    wire N__23891;
    wire N__23890;
    wire N__23889;
    wire N__23888;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23880;
    wire N__23877;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23862;
    wire N__23861;
    wire N__23860;
    wire N__23857;
    wire N__23852;
    wire N__23841;
    wire N__23840;
    wire N__23839;
    wire N__23838;
    wire N__23837;
    wire N__23820;
    wire N__23815;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23787;
    wire N__23784;
    wire N__23777;
    wire N__23766;
    wire N__23763;
    wire N__23762;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23739;
    wire N__23736;
    wire N__23735;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23709;
    wire N__23706;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23694;
    wire N__23691;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23655;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23643;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23631;
    wire N__23630;
    wire N__23627;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23580;
    wire N__23579;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23559;
    wire N__23558;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23538;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23487;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23475;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23460;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23430;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23418;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23403;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23367;
    wire N__23364;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23335;
    wire N__23330;
    wire N__23327;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23262;
    wire N__23261;
    wire N__23258;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23220;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23205;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23174;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23157;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23127;
    wire N__23124;
    wire N__23123;
    wire N__23122;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23103;
    wire N__23102;
    wire N__23101;
    wire N__23100;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23051;
    wire N__23048;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22946;
    wire N__22945;
    wire N__22942;
    wire N__22937;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22895;
    wire N__22892;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22880;
    wire N__22875;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22852;
    wire N__22847;
    wire N__22844;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22781;
    wire N__22778;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22760;
    wire N__22757;
    wire N__22756;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22744;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22683;
    wire N__22680;
    wire N__22679;
    wire N__22676;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22659;
    wire N__22656;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22638;
    wire N__22637;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22614;
    wire N__22613;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22601;
    wire N__22596;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22520;
    wire N__22519;
    wire N__22516;
    wire N__22515;
    wire N__22514;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22467;
    wire N__22462;
    wire N__22455;
    wire N__22454;
    wire N__22453;
    wire N__22452;
    wire N__22451;
    wire N__22448;
    wire N__22447;
    wire N__22444;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22408;
    wire N__22401;
    wire N__22398;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22376;
    wire N__22375;
    wire N__22372;
    wire N__22367;
    wire N__22364;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22349;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22321;
    wire N__22318;
    wire N__22313;
    wire N__22310;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22271;
    wire N__22268;
    wire N__22267;
    wire N__22264;
    wire N__22259;
    wire N__22256;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22211;
    wire N__22210;
    wire N__22207;
    wire N__22202;
    wire N__22199;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22184;
    wire N__22183;
    wire N__22180;
    wire N__22175;
    wire N__22172;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22073;
    wire N__22072;
    wire N__22069;
    wire N__22064;
    wire N__22061;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22017;
    wire N__22014;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21930;
    wire N__21927;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21915;
    wire N__21914;
    wire N__21911;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21881;
    wire N__21878;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21844;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21822;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21797;
    wire N__21794;
    wire N__21793;
    wire N__21790;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21772;
    wire N__21765;
    wire N__21764;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21746;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21734;
    wire N__21733;
    wire N__21730;
    wire N__21725;
    wire N__21720;
    wire N__21719;
    wire N__21718;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21705;
    wire N__21704;
    wire N__21703;
    wire N__21702;
    wire N__21701;
    wire N__21698;
    wire N__21693;
    wire N__21688;
    wire N__21685;
    wire N__21684;
    wire N__21683;
    wire N__21680;
    wire N__21671;
    wire N__21670;
    wire N__21663;
    wire N__21660;
    wire N__21655;
    wire N__21650;
    wire N__21647;
    wire N__21640;
    wire N__21639;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21612;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21546;
    wire N__21543;
    wire N__21542;
    wire N__21539;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21513;
    wire N__21512;
    wire N__21509;
    wire N__21508;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21494;
    wire N__21489;
    wire N__21486;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21474;
    wire N__21473;
    wire N__21470;
    wire N__21469;
    wire N__21466;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21420;
    wire N__21417;
    wire N__21410;
    wire N__21407;
    wire N__21402;
    wire N__21399;
    wire N__21398;
    wire N__21397;
    wire N__21392;
    wire N__21389;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21320;
    wire N__21315;
    wire N__21312;
    wire N__21311;
    wire N__21308;
    wire N__21303;
    wire N__21300;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21246;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21179;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21152;
    wire N__21151;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21099;
    wire N__21096;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21069;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21051;
    wire N__21050;
    wire N__21047;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21032;
    wire N__21031;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21015;
    wire N__21012;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20994;
    wire N__20993;
    wire N__20992;
    wire N__20991;
    wire N__20990;
    wire N__20989;
    wire N__20988;
    wire N__20987;
    wire N__20986;
    wire N__20985;
    wire N__20984;
    wire N__20983;
    wire N__20980;
    wire N__20975;
    wire N__20968;
    wire N__20961;
    wire N__20958;
    wire N__20953;
    wire N__20952;
    wire N__20951;
    wire N__20950;
    wire N__20941;
    wire N__20936;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20913;
    wire N__20912;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20904;
    wire N__20903;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20897;
    wire N__20896;
    wire N__20895;
    wire N__20894;
    wire N__20893;
    wire N__20888;
    wire N__20883;
    wire N__20880;
    wire N__20871;
    wire N__20864;
    wire N__20863;
    wire N__20862;
    wire N__20861;
    wire N__20860;
    wire N__20855;
    wire N__20852;
    wire N__20847;
    wire N__20842;
    wire N__20837;
    wire N__20834;
    wire N__20829;
    wire N__20820;
    wire N__20817;
    wire N__20816;
    wire N__20815;
    wire N__20812;
    wire N__20807;
    wire N__20802;
    wire N__20801;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20781;
    wire N__20780;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20768;
    wire N__20763;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20745;
    wire N__20744;
    wire N__20741;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20729;
    wire N__20724;
    wire N__20721;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20709;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20701;
    wire N__20700;
    wire N__20699;
    wire N__20690;
    wire N__20687;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20649;
    wire N__20648;
    wire N__20645;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20618;
    wire N__20617;
    wire N__20610;
    wire N__20607;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20599;
    wire N__20596;
    wire N__20591;
    wire N__20586;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20578;
    wire N__20575;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20546;
    wire N__20545;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20529;
    wire N__20524;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20514;
    wire N__20507;
    wire N__20504;
    wire N__20499;
    wire N__20498;
    wire N__20497;
    wire N__20492;
    wire N__20489;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20477;
    wire N__20476;
    wire N__20473;
    wire N__20468;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20456;
    wire N__20455;
    wire N__20452;
    wire N__20447;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20429;
    wire N__20426;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20399;
    wire N__20398;
    wire N__20395;
    wire N__20390;
    wire N__20385;
    wire N__20384;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20372;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20362;
    wire N__20359;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20316;
    wire N__20315;
    wire N__20312;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20262;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20250;
    wire N__20249;
    wire N__20246;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20234;
    wire N__20229;
    wire N__20228;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20208;
    wire N__20207;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20195;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20076;
    wire N__20073;
    wire N__20072;
    wire N__20069;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20057;
    wire N__20056;
    wire N__20051;
    wire N__20048;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19991;
    wire N__19990;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19982;
    wire N__19981;
    wire N__19976;
    wire N__19971;
    wire N__19966;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19862;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19843;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19818;
    wire N__19817;
    wire N__19816;
    wire N__19813;
    wire N__19812;
    wire N__19809;
    wire N__19808;
    wire N__19805;
    wire N__19796;
    wire N__19791;
    wire N__19788;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19769;
    wire N__19768;
    wire N__19767;
    wire N__19766;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19750;
    wire N__19743;
    wire N__19740;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19718;
    wire N__19713;
    wire N__19710;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19635;
    wire N__19634;
    wire N__19631;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19619;
    wire N__19614;
    wire N__19613;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19601;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19548;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19455;
    wire N__19452;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19422;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19389;
    wire N__19386;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19337;
    wire N__19336;
    wire N__19335;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19319;
    wire N__19316;
    wire N__19311;
    wire N__19310;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19302;
    wire N__19301;
    wire N__19298;
    wire N__19297;
    wire N__19296;
    wire N__19295;
    wire N__19282;
    wire N__19277;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire ICE_GPMO_2;
    wire VCCG0;
    wire INViac_raw_buf_vac_raw_buf_merged11WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged3WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged10WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged8WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged4WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged9WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged5WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged0WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged6WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged1WCLKN_net;
    wire ICE_SYSCLK;
    wire INViac_raw_buf_vac_raw_buf_merged7WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged2WCLKN_net;
    wire RTD_SCLK;
    wire \RTD.n8 ;
    wire RTD_SDI;
    wire \RTD.n11718 ;
    wire \RTD.n21_cascade_ ;
    wire n13176_cascade_;
    wire n18755;
    wire n13176;
    wire n18755_cascade_;
    wire \RTD.n16 ;
    wire \RTD.cfg_buf_6 ;
    wire cfg_buf_0;
    wire \RTD.n9_cascade_ ;
    wire \RTD.adress_7_N_1339_7_cascade_ ;
    wire \RTD.cfg_buf_5 ;
    wire \RTD.cfg_buf_3 ;
    wire \RTD.n11_adj_1405 ;
    wire \RTD.cfg_buf_4 ;
    wire \RTD.cfg_buf_2 ;
    wire \RTD.n10 ;
    wire \RTD.adress_7 ;
    wire \RTD.n7318 ;
    wire \RTD.n7318_cascade_ ;
    wire \RTD.n4_cascade_ ;
    wire \RTD.cfg_buf_7 ;
    wire cfg_buf_1;
    wire \RTD.n12 ;
    wire \RTD.n11 ;
    wire \RTD.n11_adj_1403 ;
    wire \RTD.n32 ;
    wire \RTD.n32_cascade_ ;
    wire \RTD.n21555 ;
    wire \RTD.n6 ;
    wire RTD_SDO;
    wire n1_adj_1606_cascade_;
    wire \RTD.n20160 ;
    wire read_buf_3;
    wire read_buf_2;
    wire DDS_MCLK1;
    wire RTD_CS;
    wire \RTD.n11687 ;
    wire adress_5;
    wire adress_6;
    wire \RTD.n19_cascade_ ;
    wire adress_0;
    wire n13165_cascade_;
    wire adress_1;
    wire n14479_cascade_;
    wire adress_4;
    wire \RTD.n21362_cascade_ ;
    wire \RTD.n1 ;
    wire n14479;
    wire adress_2;
    wire n13165;
    wire adress_3;
    wire \RTD.mode ;
    wire RTD_DRDY;
    wire \RTD.adress_7_N_1339_7 ;
    wire \RTD.n16638 ;
    wire \RTD.n16638_cascade_ ;
    wire \RTD.n20787 ;
    wire \RTD.n17835 ;
    wire \RTD.n7 ;
    wire \RTD.n11726 ;
    wire \RTD.n19787 ;
    wire \RTD.n14_cascade_ ;
    wire \RTD.n20832 ;
    wire \RTD.n11704_cascade_ ;
    wire \RTD.cfg_tmp_1 ;
    wire \RTD.cfg_tmp_2 ;
    wire \RTD.cfg_tmp_3 ;
    wire \RTD.cfg_tmp_4 ;
    wire \RTD.cfg_tmp_5 ;
    wire \RTD.cfg_tmp_6 ;
    wire \RTD.cfg_tmp_7 ;
    wire \RTD.cfg_tmp_0 ;
    wire \RTD.n11704 ;
    wire \RTD.n14999 ;
    wire read_buf_4;
    wire read_buf_0;
    wire read_buf_1;
    wire read_buf_5;
    wire read_buf_6;
    wire read_buf_12;
    wire read_buf_14;
    wire VAC_MISO;
    wire cmd_rdadctmp_0_adj_1450;
    wire cmd_rdadctmp_1_adj_1449;
    wire DDS_CS1;
    wire \CLK_DDS.n9_adj_1394 ;
    wire buf_adcdata_vac_5;
    wire buf_adcdata_iac_5;
    wire n19_adj_1629_cascade_;
    wire buf_data_iac_6;
    wire buf_adcdata_vac_4;
    wire n19_adj_1632_cascade_;
    wire buf_adcdata_iac_4;
    wire buf_adcdata_iac_6;
    wire n22_adj_1627;
    wire cmd_rdadctmp_12;
    wire cmd_rdadctmp_13;
    wire \RTD.n17799 ;
    wire \RTD.bit_cnt_3 ;
    wire \RTD.bit_cnt_1 ;
    wire \RTD.bit_cnt_2 ;
    wire \RTD.bit_cnt_0 ;
    wire \RTD.n11740 ;
    wire \CLK_DDS.n16894 ;
    wire read_buf_15;
    wire read_buf_7;
    wire buf_readRTD_10;
    wire n1_adj_1606;
    wire n13293;
    wire read_buf_10;
    wire read_buf_11;
    wire read_buf_13;
    wire buf_readRTD_13;
    wire read_buf_9;
    wire buf_readRTD_9;
    wire buf_cfgRTD_1;
    wire n14_adj_1610_cascade_;
    wire VAC_CS;
    wire cmd_rdadctmp_14;
    wire cmd_rdadctmp_2_adj_1448;
    wire cmd_rdadctmp_3_adj_1447;
    wire cmd_rdadctmp_4_adj_1446;
    wire n20864;
    wire n20864_cascade_;
    wire \ADC_VAC.n17_cascade_ ;
    wire \ADC_VAC.n12 ;
    wire IAC_CS;
    wire n14_adj_1612;
    wire n20867;
    wire n20867_cascade_;
    wire IAC_MISO;
    wire n12498_cascade_;
    wire cmd_rdadctmp_0;
    wire cmd_rdadctmp_1;
    wire cmd_rdadctmp_2;
    wire AC_ADC_SYNC;
    wire buf_adcdata_vdc_5;
    wire n19_adj_1626;
    wire cmd_rdadctmp_16_adj_1434;
    wire buf_data_iac_4;
    wire n22_adj_1633;
    wire bit_cnt_3;
    wire n21456;
    wire bit_cnt_1;
    wire bit_cnt_2;
    wire n8_adj_1602;
    wire \CLK_DDS.n9 ;
    wire cmd_rdadctmp_13_adj_1437;
    wire buf_adcdata_vac_8;
    wire buf_adcdata_vac_6;
    wire cmd_rdadctmp_14_adj_1436;
    wire cmd_rdadctmp_15_adj_1435;
    wire buf_cfgRTD_2;
    wire buf_cfgRTD_5;
    wire cmd_rdadctmp_24_adj_1426;
    wire n22321_cascade_;
    wire read_buf_8;
    wire n11714;
    wire VAC_SCLK;
    wire cmd_rdadctmp_5_adj_1445;
    wire cmd_rdadctmp_6_adj_1444;
    wire \ADC_VAC.n21312 ;
    wire \ADC_VAC.n20958_cascade_ ;
    wire \ADC_VAC.n20959 ;
    wire \ADC_VDC.n19_cascade_ ;
    wire \ADC_VDC.n18563_cascade_ ;
    wire \ADC_VDC.n18563 ;
    wire \ADC_VDC.n21384_cascade_ ;
    wire \ADC_VDC.n13034 ;
    wire \ADC_VDC.avg_cnt_0 ;
    wire bfn_8_3_0_;
    wire \ADC_VDC.n19698 ;
    wire \ADC_VDC.n19699 ;
    wire \ADC_VDC.n19700 ;
    wire \ADC_VDC.n19701 ;
    wire \ADC_VDC.n19702 ;
    wire \ADC_VDC.n19703 ;
    wire \ADC_VDC.n19704 ;
    wire \ADC_VDC.n19705 ;
    wire \ADC_VDC.avg_cnt_8 ;
    wire bfn_8_4_0_;
    wire \ADC_VDC.avg_cnt_9 ;
    wire \ADC_VDC.n19706 ;
    wire \ADC_VDC.avg_cnt_10 ;
    wire \ADC_VDC.n19707 ;
    wire \ADC_VDC.n19708 ;
    wire \ADC_VDC.n13010_cascade_ ;
    wire n12871_cascade_;
    wire cmd_rdadctmp_0_adj_1479;
    wire \ADC_VDC.cmd_rdadcbuf_0 ;
    wire bfn_8_6_0_;
    wire cmd_rdadctmp_1_adj_1478;
    wire \ADC_VDC.cmd_rdadcbuf_1 ;
    wire \ADC_VDC.n19663 ;
    wire cmd_rdadctmp_2_adj_1477;
    wire \ADC_VDC.cmd_rdadcbuf_2 ;
    wire \ADC_VDC.n19664 ;
    wire \ADC_VDC.cmd_rdadcbuf_3 ;
    wire \ADC_VDC.n19665 ;
    wire \ADC_VDC.cmd_rdadcbuf_4 ;
    wire \ADC_VDC.n19666 ;
    wire \ADC_VDC.cmd_rdadcbuf_5 ;
    wire \ADC_VDC.n19667 ;
    wire \ADC_VDC.cmd_rdadcbuf_6 ;
    wire \ADC_VDC.n19668 ;
    wire \ADC_VDC.cmd_rdadcbuf_7 ;
    wire \ADC_VDC.n19669 ;
    wire \ADC_VDC.n19670 ;
    wire \ADC_VDC.cmd_rdadcbuf_8 ;
    wire bfn_8_7_0_;
    wire \ADC_VDC.cmd_rdadcbuf_9 ;
    wire \ADC_VDC.n19671 ;
    wire \ADC_VDC.cmd_rdadcbuf_10 ;
    wire \ADC_VDC.n19672 ;
    wire cmd_rdadctmp_11_adj_1468;
    wire \ADC_VDC.n19673 ;
    wire \ADC_VDC.n19674 ;
    wire \ADC_VDC.n19675 ;
    wire \ADC_VDC.n19676 ;
    wire \ADC_VDC.n19677 ;
    wire \ADC_VDC.n19678 ;
    wire cmd_rdadcbuf_16;
    wire bfn_8_8_0_;
    wire cmd_rdadctmp_17_adj_1462;
    wire \ADC_VDC.n19679 ;
    wire \ADC_VDC.n19680 ;
    wire \ADC_VDC.n19681 ;
    wire cmd_rdadctmp_20_adj_1459;
    wire \ADC_VDC.n19682 ;
    wire cmd_rdadctmp_21_adj_1458;
    wire \ADC_VDC.n19683 ;
    wire \ADC_VDC.n19684 ;
    wire \ADC_VDC.n19685 ;
    wire \ADC_VDC.n19686 ;
    wire bfn_8_9_0_;
    wire \ADC_VDC.n19687 ;
    wire \ADC_VDC.n19688 ;
    wire \ADC_VDC.n19689 ;
    wire \ADC_VDC.n19690 ;
    wire \ADC_VDC.n19691 ;
    wire \ADC_VDC.n19692 ;
    wire \ADC_VDC.n19693 ;
    wire \ADC_VDC.n19694 ;
    wire bfn_8_10_0_;
    wire \ADC_VDC.n19695 ;
    wire \ADC_VDC.n13010 ;
    wire \ADC_VDC.n14915 ;
    wire \ADC_VDC.n19696 ;
    wire \ADC_VDC.cmd_rdadcbuf_35_N_1138_34 ;
    wire buf_adcdata_vac_16;
    wire cmd_rdadctmp_3;
    wire cmd_rdadctmp_27_adj_1423;
    wire cmd_rdadctmp_28_adj_1422;
    wire cmd_rdadctmp_29_adj_1421;
    wire cmd_rdadctmp_7_adj_1443;
    wire cmd_rdadctmp_31_adj_1419;
    wire cmd_rdadctmp_30_adj_1420;
    wire n22405;
    wire buf_adcdata_vac_21;
    wire n21097;
    wire buf_cfgRTD_4;
    wire buf_readRTD_12;
    wire buf_readRTD_4;
    wire AMPV_POW;
    wire n23_adj_1540_cascade_;
    wire n21123;
    wire EIS_SYNCCLK;
    wire IAC_CLK;
    wire cmd_rdadctmp_15;
    wire n21082;
    wire n21201;
    wire n22315_cascade_;
    wire n22318;
    wire cmd_rdadctmp_22;
    wire buf_readRTD_8;
    wire buf_cfgRTD_0;
    wire n21202;
    wire VAC_OSR1;
    wire cmd_rdadctmp_16;
    wire cmd_rdadctmp_17;
    wire VAC_DRDY;
    wire cmd_rdadctmp_18;
    wire IAC_SCLK;
    wire bfn_8_17_0_;
    wire \ADC_IAC.n19649 ;
    wire \ADC_IAC.n19650 ;
    wire \ADC_IAC.n19651 ;
    wire \ADC_IAC.n19652 ;
    wire \ADC_IAC.n19653 ;
    wire \ADC_IAC.n19654 ;
    wire \ADC_IAC.n19655 ;
    wire \ADC_IAC.n14806 ;
    wire \ADC_IAC.n17_cascade_ ;
    wire \ADC_IAC.n12 ;
    wire \ADC_VDC.avg_cnt_4 ;
    wire \ADC_VDC.avg_cnt_7 ;
    wire \ADC_VDC.avg_cnt_3 ;
    wire \ADC_VDC.avg_cnt_5 ;
    wire \ADC_VDC.n20 ;
    wire \ADC_VDC.avg_cnt_11 ;
    wire \ADC_VDC.avg_cnt_2 ;
    wire \ADC_VDC.avg_cnt_1 ;
    wire \ADC_VDC.avg_cnt_6 ;
    wire \ADC_VDC.n21 ;
    wire cmd_rdadcbuf_27;
    wire buf_adcdata_vdc_16;
    wire cmd_rdadcbuf_19;
    wire buf_adcdata_vdc_8;
    wire cmd_rdadcbuf_12;
    wire cmd_rdadcbuf_13;
    wire cmd_rdadctmp_14_adj_1465;
    wire cmd_rdadctmp_3_adj_1476;
    wire cmd_rdadctmp_4_adj_1475;
    wire cmd_rdadctmp_8_adj_1471;
    wire cmd_rdadcbuf_18;
    wire cmd_rdadctmp_5_adj_1474;
    wire cmd_rdadctmp_6_adj_1473;
    wire cmd_rdadctmp_7_adj_1472;
    wire cmd_rdadcbuf_15;
    wire buf_adcdata_vdc_4;
    wire cmd_rdadctmp_12_adj_1467;
    wire cmd_rdadctmp_13_adj_1466;
    wire cmd_rdadctmp_9_adj_1470;
    wire cmd_rdadctmp_10_adj_1469;
    wire cmd_rdadcbuf_14;
    wire cmd_rdadctmp_15_adj_1464;
    wire cmd_rdadctmp_16_adj_1463;
    wire n12871;
    wire cmd_rdadctmp_18_adj_1461;
    wire cmd_rdadctmp_19_adj_1460;
    wire cmd_rdadcbuf_25;
    wire cmd_rdadcbuf_24;
    wire cmd_rdadcbuf_17;
    wire buf_adcdata_vdc_6;
    wire cmd_rdadcbuf_23;
    wire buf_adcdata_vdc_7;
    wire buf_adcdata_vac_7;
    wire cmd_rdadcbuf_20;
    wire cmd_rdadcbuf_22;
    wire cmd_rdadcbuf_28;
    wire cmd_rdadcbuf_34;
    wire buf_adcdata_vdc_23;
    wire buf_adcdata_vac_23;
    wire cmd_rdadcbuf_32;
    wire buf_adcdata_vdc_21;
    wire cmd_rdadcbuf_31;
    wire cmd_rdadcbuf_30;
    wire cmd_rdadcbuf_29;
    wire cmd_rdadctmp_23_adj_1427;
    wire cmd_rdadctmp_26_adj_1424;
    wire buf_adcdata_vdc_17;
    wire n22441;
    wire cmd_rdadctmp_25_adj_1425;
    wire buf_adcdata_vac_17;
    wire buf_adcdata_iac_7;
    wire n19_adj_1623;
    wire buf_data_iac_7;
    wire n22_adj_1624_cascade_;
    wire bit_cnt_0_adj_1456;
    wire cmd_rdadctmp_7;
    wire DDS_MOSI1;
    wire buf_cfgRTD_3;
    wire buf_readRTD_11;
    wire buf_adcdata_vdc_12;
    wire n19_adj_1511;
    wire buf_adcdata_vdc_13;
    wire cmd_rdadctmp_21_adj_1429;
    wire buf_adcdata_vac_13;
    wire cmd_rdadctmp_22_adj_1428;
    wire cmd_rdadctmp_20_adj_1430;
    wire buf_adcdata_vac_12;
    wire cmd_rdadctmp_23;
    wire n22417;
    wire buf_adcdata_vac_20;
    wire buf_adcdata_vdc_20;
    wire cmd_rdadctmp_20;
    wire n21139;
    wire n22291;
    wire n21138_cascade_;
    wire buf_adcdata_iac_21;
    wire buf_adcdata_vac_19;
    wire n22435;
    wire buf_adcdata_vdc_19;
    wire cmd_rdadctmp_31;
    wire cmd_rdadctmp_29;
    wire cmd_rdadctmp_30;
    wire buf_adcdata_iac_23;
    wire VAC_FLT1;
    wire bfn_9_16_0_;
    wire \ADC_VAC.n19656 ;
    wire \ADC_VAC.n19657 ;
    wire \ADC_VAC.n19658 ;
    wire \ADC_VAC.n19659 ;
    wire \ADC_VAC.bit_cnt_5 ;
    wire \ADC_VAC.n19660 ;
    wire \ADC_VAC.n19661 ;
    wire \ADC_VAC.n19662 ;
    wire \ADC_IAC.n20960_cascade_ ;
    wire \ADC_IAC.n20961 ;
    wire \ADC_IAC.bit_cnt_2 ;
    wire \ADC_IAC.bit_cnt_5 ;
    wire \ADC_IAC.bit_cnt_3 ;
    wire \ADC_IAC.bit_cnt_4 ;
    wire \ADC_IAC.bit_cnt_1 ;
    wire \ADC_IAC.bit_cnt_7 ;
    wire \ADC_IAC.n21295_cascade_ ;
    wire \ADC_IAC.n21294 ;
    wire \ADC_VAC.bit_cnt_4 ;
    wire \ADC_VAC.bit_cnt_3 ;
    wire \ADC_VAC.bit_cnt_1 ;
    wire \ADC_VAC.bit_cnt_2 ;
    wire \ADC_VAC.bit_cnt_0 ;
    wire \ADC_VAC.bit_cnt_6 ;
    wire \ADC_VAC.n21029_cascade_ ;
    wire \ADC_VAC.bit_cnt_7 ;
    wire \ADC_VAC.n21043 ;
    wire \ADC_IAC.bit_cnt_6 ;
    wire \ADC_IAC.bit_cnt_0 ;
    wire \ADC_IAC.n16 ;
    wire acadc_trig;
    wire INVacadc_trig_300C_net;
    wire IAC_DRDY;
    wire \ADC_IAC.n12473 ;
    wire \ADC_VDC.n11676_cascade_ ;
    wire VDC_SCLK;
    wire \comm_spi.iclk_N_763 ;
    wire cmd_rdadcbuf_33;
    wire cmd_rdadcbuf_11;
    wire cmd_rdadcbuf_21;
    wire n13087;
    wire n13087_cascade_;
    wire cmd_rdadcbuf_26;
    wire cmd_rdadctmp_22_adj_1457;
    wire \ADC_VDC.cmd_rdadctmp_23 ;
    wire \ADC_VDC.n12899 ;
    wire \ADC_VDC.n20656 ;
    wire \comm_spi.n22860 ;
    wire \comm_spi.n22860_cascade_ ;
    wire \comm_spi.n14597 ;
    wire buf_adcdata_vdc_0;
    wire n19_adj_1484_cascade_;
    wire n22_adj_1483_cascade_;
    wire buf_data_iac_0;
    wire buf_adcdata_iac_0;
    wire cmd_rdadctmp_8_adj_1442;
    wire buf_adcdata_vac_0;
    wire cmd_rdadctmp_8;
    wire \INVcomm_spi.bit_cnt_3767__i3C_net ;
    wire adc_state_2_adj_1481;
    wire \RTD.adc_state_1 ;
    wire \RTD.adc_state_3 ;
    wire \RTD.adc_state_0 ;
    wire \RTD.n15065 ;
    wire DDS_SCK1;
    wire buf_adcdata_vdc_18;
    wire buf_adcdata_vac_18;
    wire n21081;
    wire cmd_rdadctmp_6;
    wire cmd_rdadctmp_4;
    wire cmd_rdadctmp_5;
    wire THERMOSTAT;
    wire n11347_cascade_;
    wire n11919;
    wire buf_control_7;
    wire \CLK_DDS.tmp_buf_10 ;
    wire \CLK_DDS.tmp_buf_11 ;
    wire \CLK_DDS.tmp_buf_12 ;
    wire tmp_buf_15_adj_1455;
    wire \CLK_DDS.tmp_buf_7 ;
    wire buf_dds1_8;
    wire buf_dds1_13;
    wire cmd_rdadctmp_24;
    wire buf_adcdata_iac_16;
    wire cmd_rdadctmp_26;
    wire n12395;
    wire cmd_rdadctmp_27;
    wire cmd_rdadctmp_28;
    wire n19_adj_1527;
    wire n22279_cascade_;
    wire n17_adj_1526;
    wire n23_adj_1529;
    wire n22363_cascade_;
    wire n21285;
    wire n22282;
    wire n22366_cascade_;
    wire buf_dds1_15;
    wire n16_adj_1525;
    wire adc_state_1_adj_1417;
    wire IAC_OSR0;
    wire n12367_cascade_;
    wire n16563_cascade_;
    wire n22255;
    wire iac_raw_buf_N_734;
    wire INVeis_state_i0C_net;
    wire \ADC_VDC.n21952 ;
    wire \INVcomm_spi.MISO_48_12186_12187_resetC_net ;
    wire bfn_11_5_0_;
    wire n19746;
    wire n19747;
    wire n19748;
    wire n19749;
    wire ICE_SPI_SCLK;
    wire \comm_spi.n14596 ;
    wire \comm_spi.iclk_N_762 ;
    wire buf_adcdata_vdc_2;
    wire n19_adj_1639_cascade_;
    wire buf_data_iac_5;
    wire n22_adj_1630;
    wire buf_adcdata_iac_2;
    wire cmd_rdadctmp_9;
    wire cmd_rdadctmp_10;
    wire n12498;
    wire buf_adcdata_vac_2;
    wire buf_adcdata_vdc_3;
    wire \comm_spi.bit_cnt_1 ;
    wire \comm_spi.bit_cnt_2 ;
    wire \comm_spi.bit_cnt_0 ;
    wire cmd_rdadctmp_11;
    wire buf_adcdata_vac_3;
    wire cmd_rdadctmp_10_adj_1440;
    wire cmd_rdadctmp_11_adj_1439;
    wire cmd_rdadctmp_12_adj_1438;
    wire n22_adj_1640;
    wire buf_data_iac_2;
    wire bfn_11_9_0_;
    wire n19750;
    wire n19751;
    wire n19752;
    wire n19753;
    wire n19754;
    wire n19755;
    wire n19756;
    wire n19757;
    wire bfn_11_10_0_;
    wire n19758;
    wire n19759;
    wire n19760;
    wire n19761;
    wire n19762;
    wire n19763;
    wire n19764;
    wire n19765;
    wire bfn_11_11_0_;
    wire n19766;
    wire n19767;
    wire n19768;
    wire n19769;
    wire n19770;
    wire n19771;
    wire buf_dds1_14;
    wire \CLK_DDS.tmp_buf_13 ;
    wire \CLK_DDS.tmp_buf_14 ;
    wire \CLK_DDS.tmp_buf_0 ;
    wire \CLK_DDS.tmp_buf_1 ;
    wire \CLK_DDS.tmp_buf_2 ;
    wire \CLK_DDS.tmp_buf_3 ;
    wire \CLK_DDS.tmp_buf_4 ;
    wire \CLK_DDS.tmp_buf_5 ;
    wire \CLK_DDS.tmp_buf_6 ;
    wire \CLK_DDS.tmp_buf_8 ;
    wire \CLK_DDS.tmp_buf_9 ;
    wire data_count_0;
    wire bfn_11_13_0_;
    wire data_count_1;
    wire n19586;
    wire data_count_2;
    wire n19587;
    wire data_count_3;
    wire n19588;
    wire data_count_4;
    wire n19589;
    wire data_count_5;
    wire n19590;
    wire data_count_6;
    wire n19591;
    wire data_count_7;
    wire n19592;
    wire n19593;
    wire INVdata_count_i0_i0C_net;
    wire data_count_8;
    wire bfn_11_14_0_;
    wire n19594;
    wire data_count_9;
    wire INVdata_count_i0_i8C_net;
    wire \SIG_DDS.tmp_buf_10 ;
    wire buf_dds0_5;
    wire buf_dds0_14;
    wire \SIG_DDS.tmp_buf_13 ;
    wire \SIG_DDS.tmp_buf_11 ;
    wire \SIG_DDS.tmp_buf_12 ;
    wire \SIG_DDS.tmp_buf_9 ;
    wire \SIG_DDS.tmp_buf_5 ;
    wire n16554;
    wire iac_raw_buf_N_736_cascade_;
    wire n17_adj_1622;
    wire n20826_cascade_;
    wire INVeis_end_299C_net;
    wire eis_end;
    wire n26_adj_1530;
    wire n21234;
    wire n21;
    wire n30_adj_1604_cascade_;
    wire n31;
    wire DTRIG_N_918;
    wire adc_state_1;
    wire n14_adj_1509_cascade_;
    wire n26_adj_1508;
    wire n18_adj_1609;
    wire n20915;
    wire n20985;
    wire n16571;
    wire n13_cascade_;
    wire n21337;
    wire INVeis_state_i2C_net;
    wire n17507;
    wire eis_state_0;
    wire n11_adj_1621_cascade_;
    wire n11744;
    wire eis_end_N_724;
    wire \ADC_VDC.n10119_cascade_ ;
    wire \ADC_VDC.n12807 ;
    wire bfn_12_4_0_;
    wire n19739;
    wire n19740;
    wire n19741;
    wire n19742;
    wire n19743;
    wire n19744;
    wire n19745;
    wire INVdds0_mclkcnt_i7_3772__i0C_net;
    wire clk_cnt_0;
    wire clk_cnt_4;
    wire clk_cnt_2;
    wire clk_cnt_1;
    wire n6_cascade_;
    wire clk_cnt_3;
    wire n14714;
    wire n14714_cascade_;
    wire clk_RTD;
    wire dds0_mclkcnt_3;
    wire dds0_mclkcnt_5;
    wire dds0_mclkcnt_1;
    wire dds0_mclkcnt_4;
    wire dds0_mclkcnt_2;
    wire dds0_mclkcnt_0;
    wire n12_adj_1480_cascade_;
    wire dds0_mclkcnt_7;
    wire n20799_cascade_;
    wire n10;
    wire \INVcomm_spi.imiso_83_12192_12193_resetC_net ;
    wire \comm_spi.n14611 ;
    wire \INVcomm_spi.MISO_48_12186_12187_setC_net ;
    wire \ADC_VAC.n12594 ;
    wire DTRIG_N_918_adj_1451;
    wire \ADC_VAC.n14844 ;
    wire dds0_mclkcnt_6;
    wire n20799;
    wire INVdds0_mclk_294C_net;
    wire secclk_cnt_6;
    wire secclk_cnt_14;
    wire secclk_cnt_10;
    wire secclk_cnt_3;
    wire secclk_cnt_15;
    wire secclk_cnt_8;
    wire secclk_cnt_1;
    wire secclk_cnt_5;
    wire secclk_cnt_16;
    wire secclk_cnt_2;
    wire secclk_cnt_7;
    wire secclk_cnt_13;
    wire n27_adj_1597;
    wire n26_adj_1575_cascade_;
    wire n25_adj_1574;
    wire n19856_cascade_;
    wire secclk_cnt_20;
    wire n14715;
    wire secclk_cnt_0;
    wire secclk_cnt_18;
    wire secclk_cnt_11;
    wire secclk_cnt_4;
    wire n28_adj_1505;
    wire buf_adcdata_iac_3;
    wire n19_adj_1636;
    wire secclk_cnt_17;
    wire secclk_cnt_9;
    wire n10_adj_1601;
    wire buf_data_iac_3;
    wire n22_adj_1637;
    wire cmd_rdadctmp_17_adj_1433;
    wire n12653;
    wire cmd_rdadctmp_19_adj_1431;
    wire secclk_cnt_21;
    wire secclk_cnt_19;
    wire secclk_cnt_12;
    wire secclk_cnt_22;
    wire n14_adj_1599;
    wire \comm_spi.n14610 ;
    wire \INVcomm_spi.imiso_83_12192_12193_setC_net ;
    wire buf_readRTD_14;
    wire buf_cfgRTD_6;
    wire buf_readRTD_15;
    wire buf_cfgRTD_7;
    wire n20_adj_1528;
    wire cmd_rdadctmp_19;
    wire cmd_rdadctmp_25;
    wire buf_adcdata_iac_22;
    wire VAC_FLT0;
    wire VDC_RNG0;
    wire \SIG_DDS.n10 ;
    wire buf_dds1_10;
    wire SELIRNG0;
    wire buf_dds0_1;
    wire \SIG_DDS.tmp_buf_0 ;
    wire \SIG_DDS.tmp_buf_1 ;
    wire \SIG_DDS.tmp_buf_2 ;
    wire \SIG_DDS.tmp_buf_14 ;
    wire buf_dds0_15;
    wire \SIG_DDS.tmp_buf_3 ;
    wire \SIG_DDS.tmp_buf_4 ;
    wire buf_dds0_8;
    wire \SIG_DDS.tmp_buf_8 ;
    wire \SIG_DDS.tmp_buf_6 ;
    wire buf_dds0_7;
    wire \SIG_DDS.tmp_buf_7 ;
    wire acadc_skipCount_12;
    wire acadc_skipCount_10;
    wire acadc_skipCount_13;
    wire n20;
    wire acadc_dtrig_v;
    wire acadc_dtrig_i;
    wire n4_adj_1546;
    wire n23_adj_1501;
    wire n24_adj_1642;
    wire acadc_skipCount_15;
    wire bfn_12_18_0_;
    wire INVacadc_skipcnt_i0_i0C_net;
    wire n21037;
    wire n19610;
    wire n19610_THRU_CRY_0_THRU_CO;
    wire n19610_THRU_CRY_1_THRU_CO;
    wire n19610_THRU_CRY_2_THRU_CO;
    wire n19610_THRU_CRY_3_THRU_CO;
    wire n19610_THRU_CRY_4_THRU_CO;
    wire GNDG0;
    wire n19610_THRU_CRY_5_THRU_CO;
    wire n19610_THRU_CRY_6_THRU_CO;
    wire acadc_skipcnt_1;
    wire bfn_12_19_0_;
    wire n19611;
    wire acadc_skipcnt_3;
    wire n19612;
    wire acadc_skipcnt_4;
    wire n19613;
    wire acadc_skipcnt_5;
    wire n19614;
    wire n19615;
    wire n19616;
    wire acadc_skipcnt_8;
    wire n19617;
    wire n19618;
    wire INVacadc_skipcnt_i0_i1C_net;
    wire acadc_skipcnt_9;
    wire bfn_12_20_0_;
    wire acadc_skipcnt_10;
    wire n19619;
    wire acadc_skipcnt_11;
    wire n19620;
    wire acadc_skipcnt_12;
    wire n19621;
    wire acadc_skipcnt_13;
    wire n19622;
    wire acadc_skipcnt_14;
    wire n19623;
    wire n19624;
    wire acadc_skipcnt_15;
    wire INVacadc_skipcnt_i0_i9C_net;
    wire n11654;
    wire n14671;
    wire \ADC_VDC.n17 ;
    wire \ADC_VDC.n4 ;
    wire \ADC_VDC.n7_adj_1398 ;
    wire \ADC_VDC.n7_adj_1398_cascade_ ;
    wire \ADC_VDC.n77 ;
    wire \ADC_VDC.n77_cascade_ ;
    wire \ADC_VDC.n12 ;
    wire \ADC_VDC.n20899 ;
    wire \ADC_VDC.n72_cascade_ ;
    wire \ADC_VDC.n31_cascade_ ;
    wire \ADC_VDC.n22195_cascade_ ;
    wire \ADC_VDC.n22198_cascade_ ;
    wire \ADC_VDC.n18566 ;
    wire \ADC_VDC.n20811 ;
    wire \ADC_VDC.n6_adj_1399_cascade_ ;
    wire \ADC_VDC.n10536 ;
    wire \ADC_VDC.n21229 ;
    wire \ADC_VDC.n47 ;
    wire \comm_spi.n14608 ;
    wire buf_adcdata_vdc_1;
    wire buf_adcdata_iac_1;
    wire n19_adj_1491_cascade_;
    wire buf_data_iac_1;
    wire n22_adj_1488_cascade_;
    wire n30_adj_1506;
    wire comm_buf_2_1;
    wire n22249_cascade_;
    wire n30_adj_1482;
    wire n30_adj_1625;
    wire comm_buf_2_7;
    wire n30_adj_1628;
    wire n30_adj_1631;
    wire n30_adj_1634;
    wire n30_adj_1638;
    wire n30_adj_1641;
    wire n4_adj_1594_cascade_;
    wire comm_buf_2_3;
    wire n22387_cascade_;
    wire n21193;
    wire n22390_cascade_;
    wire n4_adj_1587_cascade_;
    wire n21175_cascade_;
    wire n2358_cascade_;
    wire n20850_cascade_;
    wire n31_adj_1613_cascade_;
    wire n12085;
    wire n12085_cascade_;
    wire n14764;
    wire n12228_cascade_;
    wire comm_buf_6_7;
    wire n20850;
    wire n20852;
    wire comm_buf_6_3;
    wire buf_dds1_1;
    wire cmd_rdadctmp_9_adj_1441;
    wire buf_adcdata_vac_1;
    wire n20853;
    wire adc_state_0_adj_1418;
    wire cmd_rdadctmp_18_adj_1432;
    wire n9_adj_1416;
    wire buf_dds1_0;
    wire n22_adj_1615;
    wire n10717_cascade_;
    wire n21344;
    wire buf_dds1_5;
    wire buf_dds1_7;
    wire acadc_skipCount_14;
    wire buf_dds0_4;
    wire buf_dds1_4;
    wire buf_dds0_0;
    wire req_data_cnt_13;
    wire n19_adj_1607;
    wire n29_cascade_;
    wire n16_adj_1603;
    wire n24;
    wire n21_adj_1492_cascade_;
    wire n30_adj_1618;
    wire n20_adj_1617;
    wire n10717;
    wire req_data_cnt_12;
    wire acadc_skipCount_9;
    wire n8_adj_1573_cascade_;
    wire eis_stop;
    wire req_data_cnt_9;
    wire n22375;
    wire n22381;
    wire n22384;
    wire n11396;
    wire DDS_SCK;
    wire \comm_spi.n14605 ;
    wire \comm_spi.n14604 ;
    wire ICE_SPI_MISO;
    wire \ADC_VDC.n19_adj_1401 ;
    wire \ADC_VDC.n21323_cascade_ ;
    wire \ADC_VDC.n21320 ;
    wire \ADC_VDC.n20965 ;
    wire \ADC_VDC.n10_cascade_ ;
    wire \ADC_VDC.n20812 ;
    wire \ADC_VDC.n20784 ;
    wire \ADC_VDC.n17509 ;
    wire \ADC_VDC.n11265 ;
    wire \ADC_VDC.n6 ;
    wire \ADC_VDC.n11265_cascade_ ;
    wire \ADC_VDC.n15 ;
    wire \ADC_VDC.n15_cascade_ ;
    wire \ADC_VDC.n20996 ;
    wire dds_state_1_adj_1453;
    wire dds_state_2_adj_1452;
    wire dds_state_0_adj_1454;
    wire \CLK_DDS.n12784 ;
    wire \comm_spi.n14607 ;
    wire n21122_cascade_;
    wire n21120;
    wire n11361;
    wire n7_adj_1616_cascade_;
    wire \comm_spi.bit_cnt_3 ;
    wire \comm_spi.n17036 ;
    wire \INVcomm_spi.data_valid_85C_net ;
    wire n20858;
    wire adc_state_0;
    wire cmd_rdadctmp_21;
    wire buf_data_iac_21;
    wire n21124;
    wire \comm_spi.n14603 ;
    wire \comm_spi.data_tx_7__N_774 ;
    wire comm_tx_buf_7;
    wire \comm_spi.data_tx_7__N_766 ;
    wire n12228;
    wire buf_adcdata_vdc_9;
    wire buf_adcdata_vac_9;
    wire comm_tx_buf_3;
    wire n16891_cascade_;
    wire \SIG_DDS.n21571 ;
    wire buf_adcdata_vdc_10;
    wire buf_adcdata_vac_10;
    wire ICE_GPMI_0;
    wire n11385;
    wire n10_adj_1554_cascade_;
    wire n11850;
    wire n20914_cascade_;
    wire n21014;
    wire n17_adj_1489;
    wire \SIG_DDS.n9 ;
    wire n22_adj_1499;
    wire n18;
    wire req_data_cnt_14;
    wire n23_adj_1614;
    wire n10520;
    wire req_data_cnt_15;
    wire n8_adj_1532_cascade_;
    wire data_index_9_N_216_0;
    wire n8_adj_1532;
    wire n11338;
    wire n11338_cascade_;
    wire n8813_cascade_;
    wire data_index_0;
    wire n7;
    wire bfn_14_18_0_;
    wire data_index_1;
    wire n19625;
    wire n19626;
    wire n19627;
    wire n19628;
    wire n19629;
    wire n19630;
    wire n19631;
    wire n19632;
    wire bfn_14_19_0_;
    wire n10598;
    wire n19633;
    wire n7_adj_1572;
    wire n8_adj_1573;
    wire data_index_9_N_216_1;
    wire DDS_RNG_0;
    wire tmp_buf_15;
    wire DDS_MOSI;
    wire DDS_CS;
    wire \SIG_DDS.n9_adj_1393 ;
    wire \comm_spi.data_tx_7__N_795 ;
    wire \ADC_VDC.bit_cnt_0 ;
    wire bfn_15_4_0_;
    wire \ADC_VDC.bit_cnt_1 ;
    wire \ADC_VDC.n19772 ;
    wire \ADC_VDC.bit_cnt_2 ;
    wire \ADC_VDC.n19773 ;
    wire \ADC_VDC.bit_cnt_3 ;
    wire \ADC_VDC.n19774 ;
    wire \ADC_VDC.bit_cnt_4 ;
    wire \ADC_VDC.n19775 ;
    wire \ADC_VDC.bit_cnt_5 ;
    wire \ADC_VDC.n19776 ;
    wire \ADC_VDC.bit_cnt_6 ;
    wire \ADC_VDC.n19777 ;
    wire \ADC_VDC.n19778 ;
    wire \ADC_VDC.bit_cnt_7 ;
    wire \ADC_VDC.n18550 ;
    wire \comm_spi.data_tx_7__N_786 ;
    wire n20944_cascade_;
    wire n20964;
    wire n20962;
    wire n3;
    wire n20801;
    wire n4_adj_1586;
    wire n20801_cascade_;
    wire n19902;
    wire n22423;
    wire n2_adj_1581_cascade_;
    wire n21370_cascade_;
    wire n21369;
    wire n22426;
    wire n14;
    wire n1264_cascade_;
    wire n4_adj_1643;
    wire n1264;
    wire n8_adj_1582;
    wire comm_state_3_N_420_3;
    wire comm_state_3_N_420_3_cascade_;
    wire n21435_cascade_;
    wire n20829;
    wire n20937_cascade_;
    wire n20939;
    wire n19_adj_1522;
    wire buf_readRTD_1;
    wire buf_adcdata_iac_9;
    wire n22261_cascade_;
    wire n16_adj_1521;
    wire n26_adj_1523_cascade_;
    wire acadc_skipCount_1;
    wire n22411_cascade_;
    wire req_data_cnt_1;
    wire n22264;
    wire n22414_cascade_;
    wire n30_adj_1524_cascade_;
    wire comm_buf_1_1;
    wire \comm_spi.n14623 ;
    wire \comm_spi.data_tx_7__N_770 ;
    wire \comm_spi.n14622 ;
    wire \comm_spi.n22857 ;
    wire eis_state_1;
    wire n26_adj_1644;
    wire n20893;
    wire n21521;
    wire n14_adj_1533;
    wire bfn_15_14_0_;
    wire n14_adj_1556;
    wire data_idxvec_1;
    wire n19634;
    wire n14_adj_1555;
    wire n19635;
    wire n19636;
    wire n14_adj_1553;
    wire n19637;
    wire n14_adj_1584;
    wire n19638;
    wire n19639;
    wire n14_adj_1551;
    wire n19640;
    wire n19641;
    wire n14_adj_1550;
    wire bfn_15_15_0_;
    wire n14_adj_1580;
    wire n19642;
    wire n14_adj_1579;
    wire n19643;
    wire n19644;
    wire n14_adj_1577;
    wire data_idxvec_12;
    wire n19645;
    wire n14_adj_1583;
    wire data_idxvec_13;
    wire n19646;
    wire n14_adj_1576;
    wire data_idxvec_14;
    wire n19647;
    wire n14_adj_1549;
    wire n19648;
    wire data_idxvec_15;
    wire n12280;
    wire iac_raw_buf_N_736;
    wire bfn_15_16_0_;
    wire data_cntvec_1;
    wire n19595;
    wire n19596;
    wire n19597;
    wire n19598;
    wire n19599;
    wire n19600;
    wire n19601;
    wire n19602;
    wire INVdata_cntvec_i0_i0C_net;
    wire bfn_15_17_0_;
    wire n19603;
    wire n19604;
    wire n19605;
    wire data_cntvec_12;
    wire n19606;
    wire data_cntvec_13;
    wire n19607;
    wire data_cntvec_14;
    wire n19608;
    wire n19609;
    wire data_cntvec_15;
    wire INVdata_cntvec_i0_i8C_net;
    wire n13457;
    wire n14647;
    wire acadc_skipcnt_0;
    wire acadc_skipcnt_6;
    wire n17;
    wire n8_adj_1565_cascade_;
    wire data_index_6;
    wire data_index_9_N_216_3;
    wire n8_adj_1565;
    wire n7_adj_1564;
    wire data_index_9_N_216_6;
    wire data_index_9;
    wire n8_adj_1559;
    wire n7_adj_1558;
    wire n8_adj_1559_cascade_;
    wire data_index_9_N_216_9;
    wire n7_adj_1560;
    wire data_index_9_N_216_8;
    wire data_index_9_N_216_7;
    wire clk_16MHz;
    wire dds0_mclk;
    wire buf_control_6;
    wire DDS_MCLK;
    wire \comm_spi.n14619 ;
    wire \comm_spi.n22884 ;
    wire \comm_spi.n22884_cascade_ ;
    wire \comm_spi.n14593 ;
    wire \comm_spi.n14618 ;
    wire \comm_spi.data_tx_7__N_772 ;
    wire \comm_spi.data_tx_7__N_792 ;
    wire \comm_spi.n22881 ;
    wire \comm_spi.data_tx_7__N_789 ;
    wire \comm_spi.data_tx_7__N_771 ;
    wire \comm_spi.n22878 ;
    wire wdtick_cnt_2;
    wire wdtick_cnt_0;
    wire wdtick_cnt_1;
    wire TEST_LED;
    wire \comm_spi.n14627 ;
    wire \comm_spi.n22875 ;
    wire \comm_spi.n14626 ;
    wire n11741;
    wire n20992;
    wire n9255_cascade_;
    wire n14737;
    wire flagcntwd;
    wire n11390;
    wire n12336_cascade_;
    wire n20378;
    wire comm_buf_2_4;
    wire comm_buf_6_4;
    wire n21538_cascade_;
    wire n1_adj_1591;
    wire n22369_cascade_;
    wire n2_adj_1592;
    wire n4_adj_1593;
    wire \comm_spi.data_tx_7__N_783 ;
    wire comm_tx_buf_4;
    wire \comm_spi.data_tx_7__N_769 ;
    wire comm_buf_2_2;
    wire n22393_cascade_;
    wire comm_buf_6_2;
    wire n4_adj_1595_cascade_;
    wire n22396;
    wire n21196_cascade_;
    wire comm_tx_buf_2;
    wire comm_buf_6_1;
    wire n4_adj_1596_cascade_;
    wire n22252;
    wire n21052_cascade_;
    wire comm_tx_buf_1;
    wire buf_data_vac_0;
    wire buf_data_vac_7;
    wire comm_buf_5_7;
    wire buf_data_vac_6;
    wire buf_data_vac_5;
    wire buf_data_vac_4;
    wire comm_buf_5_4;
    wire buf_data_vac_3;
    wire comm_buf_5_3;
    wire buf_data_vac_2;
    wire comm_buf_5_2;
    wire buf_data_vac_1;
    wire comm_buf_5_1;
    wire IAC_OSR1;
    wire buf_adcdata_iac_17;
    wire buf_dds0_9;
    wire n22237_cascade_;
    wire buf_dds1_9;
    wire buf_data_iac_17;
    wire n22378;
    wire n21062_cascade_;
    wire n22240;
    wire n22444;
    wire n22447_cascade_;
    wire n22450_cascade_;
    wire comm_buf_0_1;
    wire n30;
    wire n21272;
    wire n23_adj_1538;
    wire n22273_cascade_;
    wire n21286;
    wire n17_adj_1535;
    wire n16_adj_1534;
    wire n22288_cascade_;
    wire n22276;
    wire n30_adj_1539_cascade_;
    wire buf_adcdata_vdc_22;
    wire buf_adcdata_vac_22;
    wire n20_adj_1537;
    wire n19_adj_1536_cascade_;
    wire n22285;
    wire buf_adcdata_iac_20;
    wire buf_dds0_12;
    wire n22303_cascade_;
    wire buf_dds1_12;
    wire n21309;
    wire n23_adj_1541;
    wire n21568;
    wire n22243;
    wire n22306;
    wire n22420;
    wire n22246;
    wire n21092_cascade_;
    wire n30_adj_1542_cascade_;
    wire n21087;
    wire n22357_cascade_;
    wire n22360_cascade_;
    wire n21137_cascade_;
    wire n21072;
    wire n22327;
    wire n22330;
    wire data_idxvec_11;
    wire data_cntvec_11;
    wire buf_data_iac_19;
    wire n26_adj_1544_cascade_;
    wire acadc_rst;
    wire req_data_cnt_10;
    wire n21088;
    wire req_data_cnt_6;
    wire buf_dds1_6;
    wire buf_dds0_6;
    wire buf_adcdata_iac_18;
    wire n21073;
    wire n16891;
    wire data_index_5;
    wire data_idxvec_10;
    wire data_cntvec_10;
    wire n21150;
    wire data_idxvec_9;
    wire data_cntvec_9;
    wire n21060;
    wire n8_adj_1569;
    wire n7_adj_1568;
    wire data_index_3;
    wire data_idxvec_8;
    wire data_cntvec_8;
    wire req_data_cnt_11;
    wire n8_adj_1571_cascade_;
    wire data_index_2;
    wire buf_dds0_10;
    wire n20907;
    wire n12429;
    wire n9306_cascade_;
    wire buf_dds0_13;
    wire acadc_skipcnt_7;
    wire acadc_skipcnt_2;
    wire n22;
    wire n9;
    wire n20912;
    wire comm_buf_0_4;
    wire n12381_cascade_;
    wire VAC_OSR0;
    wire acadc_skipCount_6;
    wire dds_state_0;
    wire dds_state_2;
    wire trig_dds0;
    wire \SIG_DDS.n12722 ;
    wire data_index_8;
    wire n8_adj_1561;
    wire n8_adj_1563;
    wire n7_adj_1562;
    wire data_index_7;
    wire SELIRNG1;
    wire acadc_skipCount_11;
    wire n23_adj_1543;
    wire n11915;
    wire buf_data_iac_22;
    wire n21273;
    wire buf_data_iac_20;
    wire n21569;
    wire \comm_spi.n14592 ;
    wire \comm_spi.n14639 ;
    wire \comm_spi.data_tx_7__N_777 ;
    wire \comm_spi.data_tx_7__N_780 ;
    wire comm_buf_5_6;
    wire n22183_cascade_;
    wire comm_buf_5_0;
    wire n4;
    wire comm_buf_6_0;
    wire n21211;
    wire n1;
    wire comm_buf_2_0;
    wire n2;
    wire comm_tx_buf_0;
    wire \comm_spi.data_tx_7__N_773 ;
    wire n17479_cascade_;
    wire comm_buf_6_5;
    wire comm_buf_2_5;
    wire n17480;
    wire comm_buf_5_5;
    wire n21212;
    wire n17482_cascade_;
    wire n22189;
    wire comm_tx_buf_5;
    wire buf_data_vac_8;
    wire comm_buf_4_0;
    wire buf_data_vac_15;
    wire comm_buf_4_7;
    wire buf_data_vac_14;
    wire comm_buf_4_6;
    wire buf_data_vac_13;
    wire comm_buf_4_5;
    wire buf_data_vac_12;
    wire comm_buf_4_4;
    wire buf_data_vac_11;
    wire comm_buf_4_3;
    wire buf_data_vac_10;
    wire comm_buf_4_2;
    wire buf_data_vac_9;
    wire comm_buf_4_1;
    wire \SIG_DDS.bit_cnt_3 ;
    wire bit_cnt_0;
    wire \SIG_DDS.bit_cnt_1 ;
    wire \SIG_DDS.bit_cnt_2 ;
    wire dds_state_1;
    wire n14884;
    wire n12220;
    wire n12220_cascade_;
    wire n14785;
    wire n14778;
    wire n30_adj_1531;
    wire comm_buf_0_7;
    wire n22324;
    wire comm_buf_0_5;
    wire buf_adcdata_iac_8;
    wire n16_adj_1487;
    wire n19_adj_1486;
    wire buf_readRTD_0;
    wire n22213;
    wire data_idxvec_0;
    wire data_cntvec_0;
    wire n26_cascade_;
    wire acadc_skipCount_0;
    wire n22201_cascade_;
    wire req_data_cnt_0;
    wire n22216;
    wire n22204_cascade_;
    wire n30_adj_1485_cascade_;
    wire comm_buf_1_0;
    wire buf_adcdata_iac_19;
    wire buf_dds0_11;
    wire n22297_cascade_;
    wire buf_dds1_11;
    wire n21076;
    wire n22300;
    wire n22312_cascade_;
    wire eis_start;
    wire req_data_cnt_8;
    wire n22294;
    wire n21071_cascade_;
    wire comm_buf_0_0;
    wire n14750;
    wire n22219;
    wire acadc_skipCount_8;
    wire n14_adj_1578;
    wire n9_adj_1415;
    wire buf_data_iac_16;
    wire n21165;
    wire n21167_cascade_;
    wire n22222;
    wire n21070;
    wire n21084;
    wire n21085;
    wire n22309;
    wire n12399;
    wire comm_buf_0_3;
    wire IAC_FLT1;
    wire n20914;
    wire trig_dds1;
    wire n8_adj_1571;
    wire n7_adj_1570;
    wire data_index_9_N_216_2;
    wire n11819;
    wire n12381;
    wire comm_buf_0_2;
    wire IAC_FLT0;
    wire wdtick_flag;
    wire buf_control_0;
    wire CONT_SD;
    wire \comm_spi.imosi_N_753 ;
    wire \comm_spi.n22872 ;
    wire \comm_spi.n14630 ;
    wire \comm_spi.n14631 ;
    wire \comm_spi.data_tx_7__N_768 ;
    wire \comm_spi.n22869 ;
    wire \comm_spi.n14634 ;
    wire \comm_spi.n14635 ;
    wire \comm_spi.n14638 ;
    wire \ADC_VDC.genclk.n21446_cascade_ ;
    wire \ADC_VDC.genclk.n26 ;
    wire \ADC_VDC.genclk.n27 ;
    wire \ADC_VDC.genclk.n28_adj_1397 ;
    wire \comm_spi.data_tx_7__N_767 ;
    wire comm_buf_0_6;
    wire n1_adj_1588_cascade_;
    wire comm_tx_buf_6;
    wire n12336;
    wire n14799;
    wire comm_buf_2_6;
    wire n2_adj_1589;
    wire comm_buf_6_6;
    wire n4_adj_1590;
    wire n21539_cascade_;
    wire n22339;
    wire buf_data_vac_16;
    wire comm_buf_3_0;
    wire buf_data_vac_20;
    wire comm_buf_3_4;
    wire buf_data_vac_23;
    wire comm_buf_3_7;
    wire buf_data_vac_22;
    wire comm_buf_3_6;
    wire buf_data_vac_21;
    wire comm_buf_3_5;
    wire buf_data_vac_19;
    wire comm_buf_3_3;
    wire buf_data_vac_18;
    wire comm_buf_3_2;
    wire comm_rx_buf_1;
    wire buf_data_vac_17;
    wire comm_buf_3_1;
    wire n20878;
    wire n21352_cascade_;
    wire n12_cascade_;
    wire n12136;
    wire n12136_cascade_;
    wire n14771;
    wire n19783;
    wire n18991_cascade_;
    wire n4_adj_1545_cascade_;
    wire n11961;
    wire n18993_cascade_;
    wire n12_adj_1605;
    wire n11991_cascade_;
    wire n14506;
    wire n11896;
    wire n10697;
    wire n18993;
    wire n20843;
    wire n12_adj_1635_cascade_;
    wire n20917;
    wire n12178;
    wire n21177;
    wire n22225_cascade_;
    wire data_idxvec_6;
    wire data_cntvec_6;
    wire buf_data_iac_14;
    wire n26_adj_1507_cascade_;
    wire n21178;
    wire comm_rx_buf_6;
    wire n22228;
    wire buf_adcdata_vdc_14;
    wire buf_adcdata_vac_14;
    wire n19_cascade_;
    wire buf_readRTD_6;
    wire n21046;
    wire n16_adj_1510;
    wire buf_adcdata_iac_12;
    wire n22231;
    wire data_idxvec_4;
    wire data_cntvec_4;
    wire n26_adj_1512_cascade_;
    wire acadc_skipCount_4;
    wire n22351_cascade_;
    wire req_data_cnt_4;
    wire n22234;
    wire n22354_cascade_;
    wire comm_rx_buf_4;
    wire n30_adj_1513_cascade_;
    wire n19_adj_1518;
    wire buf_readRTD_2;
    wire buf_adcdata_iac_10;
    wire n22207_cascade_;
    wire req_data_cnt_2;
    wire n22429_cascade_;
    wire acadc_skipCount_2;
    wire n22210;
    wire n22432_cascade_;
    wire comm_rx_buf_2;
    wire n30_adj_1520_cascade_;
    wire data_idxvec_2;
    wire data_cntvec_2;
    wire n26_adj_1519;
    wire n14_adj_1585;
    wire n8;
    wire buf_adcdata_iac_14;
    wire n16;
    wire n21045;
    wire req_data_cnt_7;
    wire acadc_skipCount_7;
    wire buf_dds1_3;
    wire buf_dds0_3;
    wire buf_dds1_2;
    wire n16_adj_1517;
    wire comm_buf_1_2;
    wire n12367;
    wire buf_dds0_2;
    wire comm_buf_1_6;
    wire n14_adj_1552;
    wire comm_buf_1_4;
    wire data_index_4;
    wire n8813;
    wire n8_adj_1567;
    wire n7_adj_1566;
    wire data_index_9_N_216_4;
    wire \ADC_VDC.n11750 ;
    wire VDC_SDO;
    wire \ADC_VDC.adc_state_0 ;
    wire \ADC_VDC.n62 ;
    wire adc_state_2;
    wire adc_state_3;
    wire \ADC_VDC.n62_cascade_ ;
    wire \ADC_VDC.adc_state_1 ;
    wire \ADC_VDC.n11 ;
    wire \ADC_VDC.genclk.t0off_0 ;
    wire bfn_19_7_0_;
    wire \ADC_VDC.genclk.t0off_1 ;
    wire \ADC_VDC.genclk.n19709 ;
    wire \ADC_VDC.genclk.t0off_2 ;
    wire \ADC_VDC.genclk.n19710 ;
    wire \ADC_VDC.genclk.t0off_3 ;
    wire \ADC_VDC.genclk.n19711 ;
    wire \ADC_VDC.genclk.t0off_4 ;
    wire \ADC_VDC.genclk.n19712 ;
    wire \ADC_VDC.genclk.t0off_5 ;
    wire \ADC_VDC.genclk.n19713 ;
    wire \ADC_VDC.genclk.t0off_6 ;
    wire \ADC_VDC.genclk.n19714 ;
    wire \ADC_VDC.genclk.t0off_7 ;
    wire \ADC_VDC.genclk.n19715 ;
    wire \ADC_VDC.genclk.n19716 ;
    wire \INVADC_VDC.genclk.t0off_i0C_net ;
    wire \ADC_VDC.genclk.t0off_8 ;
    wire bfn_19_8_0_;
    wire \ADC_VDC.genclk.t0off_9 ;
    wire \ADC_VDC.genclk.n19717 ;
    wire \ADC_VDC.genclk.t0off_10 ;
    wire \ADC_VDC.genclk.n19718 ;
    wire \ADC_VDC.genclk.t0off_11 ;
    wire \ADC_VDC.genclk.n19719 ;
    wire \ADC_VDC.genclk.t0off_12 ;
    wire \ADC_VDC.genclk.n19720 ;
    wire \ADC_VDC.genclk.t0off_13 ;
    wire \ADC_VDC.genclk.n19721 ;
    wire \ADC_VDC.genclk.t0off_14 ;
    wire \ADC_VDC.genclk.n19722 ;
    wire \ADC_VDC.genclk.n19723 ;
    wire \ADC_VDC.genclk.t0off_15 ;
    wire \INVADC_VDC.genclk.t0off_i8C_net ;
    wire \ADC_VDC.genclk.n11735 ;
    wire n14529;
    wire n17815;
    wire n23_adj_1620;
    wire n21_adj_1598_cascade_;
    wire n17564;
    wire n2358;
    wire n20856;
    wire n15_cascade_;
    wire n18_adj_1619;
    wire n14130;
    wire n20880;
    wire n20880_cascade_;
    wire n12_adj_1548;
    wire ICE_SPI_CE0;
    wire comm_data_vld;
    wire n18984;
    wire comm_cmd_4;
    wire comm_cmd_6;
    wire comm_cmd_5;
    wire n21546;
    wire n12092;
    wire n12219;
    wire n9255;
    wire n11853_cascade_;
    wire n12226;
    wire comm_state_0;
    wire n18991;
    wire n20804;
    wire n21341;
    wire n21339_cascade_;
    wire n38_adj_1608;
    wire n21054;
    wire n22267_cascade_;
    wire data_idxvec_7;
    wire data_cntvec_7;
    wire buf_data_iac_15;
    wire n26_adj_1502_cascade_;
    wire n21055;
    wire comm_rx_buf_7;
    wire n22270;
    wire comm_buf_1_7;
    wire buf_adcdata_vdc_15;
    wire buf_adcdata_vac_15;
    wire n19_adj_1503_cascade_;
    wire buf_readRTD_7;
    wire n21049;
    wire buf_readRTD_3;
    wire req_data_cnt_3;
    wire acadc_skipCount_3;
    wire n21132_cascade_;
    wire n21127;
    wire n22333_cascade_;
    wire comm_rx_buf_3;
    wire n22336_cascade_;
    wire comm_buf_1_3;
    wire buf_adcdata_vdc_11;
    wire buf_adcdata_vac_11;
    wire n19_adj_1515;
    wire data_idxvec_3;
    wire data_cntvec_3;
    wire buf_data_iac_11;
    wire n26_adj_1516_cascade_;
    wire n21133;
    wire n21316_cascade_;
    wire comm_length_2;
    wire comm_index_0;
    wire comm_index_2;
    wire n4_adj_1600;
    wire n4_adj_1600_cascade_;
    wire comm_index_1;
    wire n5_cascade_;
    wire comm_cmd_7;
    wire n21888;
    wire n21317;
    wire buf_adcdata_iac_15;
    wire n16_adj_1504;
    wire n21048;
    wire comm_rx_buf_5;
    wire comm_state_1;
    wire comm_buf_1_5;
    wire n11991;
    wire n14757;
    wire n19_adj_1497;
    wire buf_readRTD_5;
    wire data_idxvec_5;
    wire data_cntvec_5;
    wire n26_adj_1498_cascade_;
    wire req_data_cnt_5;
    wire n22345_cascade_;
    wire acadc_skipCount_5;
    wire n22348_cascade_;
    wire n30_adj_1500;
    wire buf_adcdata_iac_11;
    wire n16_adj_1514;
    wire n21126;
    wire buf_data_iac_10;
    wire n21564;
    wire buf_data_iac_8;
    wire n21218;
    wire buf_data_iac_23;
    wire n21364;
    wire \INVADC_VDC.genclk.div_state_i1C_net ;
    wire \ADC_VDC.genclk.n6 ;
    wire \comm_spi.iclk ;
    wire \ADC_VDC.genclk.n21444 ;
    wire \comm_spi.DOUT_7__N_747 ;
    wire VDC_CLK;
    wire \INVADC_VDC.genclk.div_state_i0C_net ;
    wire \comm_spi.n14614 ;
    wire \comm_spi.n14615 ;
    wire comm_rx_buf_0;
    wire \comm_spi.n22866 ;
    wire \comm_spi.n22866_cascade_ ;
    wire \comm_spi.n14601 ;
    wire \comm_spi.imosi_cascade_ ;
    wire \comm_spi.DOUT_7__N_746 ;
    wire \ADC_VDC.genclk.div_state_0 ;
    wire \comm_spi.imosi ;
    wire \comm_spi.n22863 ;
    wire \comm_spi.n14600 ;
    wire comm_clear;
    wire ICE_SPI_MOSI;
    wire \comm_spi.imosi_N_752 ;
    wire comm_state_2;
    wire comm_length_0;
    wire comm_cmd_1;
    wire comm_cmd_3;
    wire comm_length_1;
    wire clk_32MHz;
    wire n11860;
    wire n14655;
    wire buf_data_iac_12;
    wire n21451;
    wire buf_data_iac_18;
    wire n21151;
    wire n16_adj_1496;
    wire n22399;
    wire buf_adcdata_iac_13;
    wire comm_cmd_2;
    wire n22402;
    wire buf_data_iac_13;
    wire n21350;
    wire buf_data_iac_9;
    wire comm_cmd_0;
    wire n21529;
    wire comm_state_3;
    wire n17489;
    wire n9306;
    wire n17487;
    wire data_index_9_N_216_5;
    wire bfn_22_7_0_;
    wire \ADC_VDC.genclk.n19724 ;
    wire \ADC_VDC.genclk.n19725 ;
    wire \ADC_VDC.genclk.n19726 ;
    wire \ADC_VDC.genclk.n19727 ;
    wire \ADC_VDC.genclk.n19728 ;
    wire \ADC_VDC.genclk.n19729 ;
    wire \ADC_VDC.genclk.n19730 ;
    wire \ADC_VDC.genclk.n19731 ;
    wire \INVADC_VDC.genclk.t0on_i0C_net ;
    wire bfn_22_8_0_;
    wire \ADC_VDC.genclk.n19732 ;
    wire \ADC_VDC.genclk.n19733 ;
    wire \ADC_VDC.genclk.n19734 ;
    wire \ADC_VDC.genclk.n19735 ;
    wire \ADC_VDC.genclk.n19736 ;
    wire \ADC_VDC.genclk.n19737 ;
    wire CONSTANT_ONE_NET;
    wire \ADC_VDC.genclk.n19738 ;
    wire \INVADC_VDC.genclk.t0on_i8C_net ;
    wire \ADC_VDC.genclk.n15051 ;
    wire \ADC_VDC.genclk.t0on_6 ;
    wire \ADC_VDC.genclk.t0on_1 ;
    wire \ADC_VDC.genclk.t0on_4 ;
    wire \ADC_VDC.genclk.t0on_0 ;
    wire \ADC_VDC.genclk.n21449_cascade_ ;
    wire \ADC_VDC.genclk.n21443 ;
    wire \ADC_VDC.genclk.t0on_12 ;
    wire \ADC_VDC.genclk.t0on_2 ;
    wire \ADC_VDC.genclk.t0on_7 ;
    wire \ADC_VDC.genclk.t0on_10 ;
    wire \ADC_VDC.genclk.n27_adj_1396 ;
    wire \ADC_VDC.genclk.t0on_3 ;
    wire \ADC_VDC.genclk.t0on_13 ;
    wire \ADC_VDC.genclk.t0on_5 ;
    wire \ADC_VDC.genclk.t0on_8 ;
    wire \ADC_VDC.genclk.n26_adj_1395 ;
    wire \ADC_VDC.genclk.div_state_1 ;
    wire \ADC_VDC.genclk.div_state_1__N_1274 ;
    wire \ADC_VDC.genclk.t0on_14 ;
    wire \ADC_VDC.genclk.t0on_9 ;
    wire \ADC_VDC.genclk.t0on_15 ;
    wire \ADC_VDC.genclk.t0on_11 ;
    wire \ADC_VDC.genclk.n28 ;
    wire _gnd_net_;

    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_main.zim_pll_inst .TEST_MODE=1'b0;
    defparam \pll_main.zim_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll_main.zim_pll_inst .FILTER_RANGE=3'b011;
    defparam \pll_main.zim_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_main.zim_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_main.zim_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll_main.zim_pll_inst .DIVR=4'b0000;
    defparam \pll_main.zim_pll_inst .DIVQ=3'b101;
    defparam \pll_main.zim_pll_inst .DIVF=7'b0011111;
    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll_main.zim_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(),
            .REFERENCECLK(N__19206),
            .RESETB(N__58564),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(clk_16MHz),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(clk_32MHz),
            .SCLK(GNDG0));
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged2_physical (
            .RDATA({dangling_wire_0,dangling_wire_1,buf_data_iac_19,dangling_wire_2,dangling_wire_3,dangling_wire_4,buf_data_vac_19,dangling_wire_5,dangling_wire_6,dangling_wire_7,buf_data_iac_18,dangling_wire_8,dangling_wire_9,dangling_wire_10,buf_data_vac_18,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__39015,N__38916,N__38829,N__38232,N__55983,N__47577,N__38352,N__45051,N__36435,N__36177}),
            .WADDR({dangling_wire_13,N__29544,N__29655,N__29754,N__28701,N__28809,N__28920,N__29025,N__29133,N__29241,N__29352}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__43230,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__25290,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__40716,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__27084,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__54379),
            .RE(N__58508),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .WE(N__27730));
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged7_physical (
            .RDATA({dangling_wire_42,dangling_wire_43,buf_data_iac_9,dangling_wire_44,dangling_wire_45,dangling_wire_46,buf_data_vac_9,dangling_wire_47,dangling_wire_48,dangling_wire_49,buf_data_iac_8,dangling_wire_50,dangling_wire_51,dangling_wire_52,buf_data_vac_8,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__38972,N__38873,N__38786,N__38192,N__55940,N__47531,N__38315,N__45008,N__36395,N__36137}),
            .WADDR({dangling_wire_55,N__29507,N__29618,N__29714,N__28658,N__28769,N__28883,N__28994,N__29099,N__29204,N__29318}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__37176,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__34941,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__43517,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__21576,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__54437),
            .RE(N__58607),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .WE(N__27707));
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged1_physical (
            .RDATA({dangling_wire_84,dangling_wire_85,buf_data_iac_21,dangling_wire_86,dangling_wire_87,dangling_wire_88,buf_data_vac_21,dangling_wire_89,dangling_wire_90,dangling_wire_91,buf_data_iac_20,dangling_wire_92,dangling_wire_93,dangling_wire_94,buf_data_vac_20,dangling_wire_95}),
            .RADDR({dangling_wire_96,N__39033,N__38934,N__38847,N__38250,N__56001,N__47595,N__38370,N__45069,N__36453,N__36195}),
            .WADDR({dangling_wire_97,N__29562,N__29673,N__29772,N__28719,N__28827,N__28938,N__29043,N__29151,N__29259,N__29370}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({dangling_wire_114,dangling_wire_115,N__25002,dangling_wire_116,dangling_wire_117,dangling_wire_118,N__22830,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__40386,dangling_wire_122,dangling_wire_123,dangling_wire_124,N__25098,dangling_wire_125}),
            .RCLKE(),
            .RCLK(N__54299),
            .RE(N__58359),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .WE(N__27758));
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged6_physical (
            .RDATA({dangling_wire_126,dangling_wire_127,buf_data_iac_11,dangling_wire_128,dangling_wire_129,dangling_wire_130,buf_data_vac_11,dangling_wire_131,dangling_wire_132,dangling_wire_133,buf_data_iac_10,dangling_wire_134,dangling_wire_135,dangling_wire_136,buf_data_vac_10,dangling_wire_137}),
            .RADDR({dangling_wire_138,N__38984,N__38885,N__38798,N__38204,N__55952,N__47543,N__38327,N__45020,N__36407,N__36149}),
            .WADDR({dangling_wire_139,N__29519,N__29630,N__29726,N__28670,N__28781,N__28895,N__29001,N__29109,N__29216,N__29328}),
            .MASK({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155}),
            .WDATA({dangling_wire_156,dangling_wire_157,N__52788,dangling_wire_158,dangling_wire_159,dangling_wire_160,N__50921,dangling_wire_161,dangling_wire_162,dangling_wire_163,N__46647,dangling_wire_164,dangling_wire_165,dangling_wire_166,N__35961,dangling_wire_167}),
            .RCLKE(),
            .RCLK(N__54435),
            .RE(N__58585),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .WE(N__27706));
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged0_physical (
            .RDATA({dangling_wire_168,dangling_wire_169,buf_data_iac_23,dangling_wire_170,dangling_wire_171,dangling_wire_172,buf_data_vac_23,dangling_wire_173,dangling_wire_174,dangling_wire_175,buf_data_iac_22,dangling_wire_176,dangling_wire_177,dangling_wire_178,buf_data_vac_22,dangling_wire_179}),
            .RADDR({dangling_wire_180,N__39039,N__38940,N__38853,N__38256,N__56007,N__47601,N__38376,N__45075,N__36459,N__36201}),
            .WADDR({dangling_wire_181,N__29568,N__29679,N__29778,N__28725,N__28833,N__28944,N__29049,N__29157,N__29265,N__29376}),
            .MASK({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .WDATA({dangling_wire_198,dangling_wire_199,N__25164,dangling_wire_200,dangling_wire_201,dangling_wire_202,N__24192,dangling_wire_203,dangling_wire_204,dangling_wire_205,N__31938,dangling_wire_206,dangling_wire_207,dangling_wire_208,N__40434,dangling_wire_209}),
            .RCLKE(),
            .RCLK(N__54284),
            .RE(N__58507),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .WE(N__27759));
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged5_physical (
            .RDATA({dangling_wire_210,dangling_wire_211,buf_data_iac_13,dangling_wire_212,dangling_wire_213,dangling_wire_214,buf_data_vac_13,dangling_wire_215,dangling_wire_216,dangling_wire_217,buf_data_iac_12,dangling_wire_218,dangling_wire_219,dangling_wire_220,buf_data_vac_12,dangling_wire_221}),
            .RADDR({dangling_wire_222,N__38996,N__38897,N__38810,N__38214,N__55964,N__47555,N__38334,N__45032,N__36417,N__36159}),
            .WADDR({dangling_wire_223,N__29526,N__29637,N__29736,N__28682,N__28791,N__28902,N__29007,N__29115,N__29223,N__29334}),
            .MASK({dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .WDATA({dangling_wire_240,dangling_wire_241,N__53832,dangling_wire_242,dangling_wire_243,dangling_wire_244,N__24927,dangling_wire_245,dangling_wire_246,dangling_wire_247,N__46268,dangling_wire_248,dangling_wire_249,dangling_wire_250,N__24861,dangling_wire_251}),
            .RCLKE(),
            .RCLK(N__54433),
            .RE(N__58566),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .WE(N__27708));
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged9_physical (
            .RDATA({dangling_wire_252,dangling_wire_253,buf_data_iac_5,dangling_wire_254,dangling_wire_255,dangling_wire_256,buf_data_vac_5,dangling_wire_257,dangling_wire_258,dangling_wire_259,buf_data_iac_4,dangling_wire_260,dangling_wire_261,dangling_wire_262,buf_data_vac_4,dangling_wire_263}),
            .RADDR({dangling_wire_264,N__38987,N__38888,N__38801,N__38201,N__55955,N__47552,N__38318,N__45023,N__36404,N__36146}),
            .WADDR({dangling_wire_265,N__29510,N__29621,N__29723,N__28673,N__28778,N__28886,N__28985,N__29096,N__29207,N__29315}),
            .MASK({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281}),
            .WDATA({dangling_wire_282,dangling_wire_283,N__20463,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__20484,dangling_wire_287,dangling_wire_288,dangling_wire_289,N__20406,dangling_wire_290,dangling_wire_291,dangling_wire_292,N__20430,dangling_wire_293}),
            .RCLKE(),
            .RCLK(N__54337),
            .RE(N__58584),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .WE(N__27756));
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged4_physical (
            .RDATA({dangling_wire_294,dangling_wire_295,buf_data_iac_15,dangling_wire_296,dangling_wire_297,dangling_wire_298,buf_data_vac_15,dangling_wire_299,dangling_wire_300,dangling_wire_301,buf_data_iac_14,dangling_wire_302,dangling_wire_303,dangling_wire_304,buf_data_vac_14,dangling_wire_305}),
            .RADDR({dangling_wire_306,N__39003,N__38904,N__38817,N__38220,N__55971,N__47565,N__38340,N__45039,N__36423,N__36165}),
            .WADDR({dangling_wire_307,N__29532,N__29643,N__29742,N__28689,N__28797,N__28908,N__29013,N__29121,N__29229,N__29340}),
            .MASK({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323}),
            .WDATA({dangling_wire_324,dangling_wire_325,N__52188,dangling_wire_326,dangling_wire_327,dangling_wire_328,N__50220,dangling_wire_329,dangling_wire_330,dangling_wire_331,N__47046,dangling_wire_332,dangling_wire_333,dangling_wire_334,N__46353,dangling_wire_335}),
            .RCLKE(),
            .RCLK(N__54425),
            .RE(N__58565),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .WE(N__27709));
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged8_physical (
            .RDATA({dangling_wire_336,dangling_wire_337,buf_data_iac_7,dangling_wire_338,dangling_wire_339,dangling_wire_340,buf_data_vac_7,dangling_wire_341,dangling_wire_342,dangling_wire_343,buf_data_iac_6,dangling_wire_344,dangling_wire_345,dangling_wire_346,buf_data_vac_6,dangling_wire_347}),
            .RADDR({dangling_wire_348,N__38999,N__38900,N__38813,N__38213,N__55967,N__47564,N__38330,N__45035,N__36416,N__36158}),
            .WADDR({dangling_wire_349,N__29522,N__29633,N__29735,N__28685,N__28790,N__28898,N__28997,N__29108,N__29219,N__29327}),
            .MASK({dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .WDATA({dangling_wire_366,dangling_wire_367,N__24834,dangling_wire_368,dangling_wire_369,dangling_wire_370,N__24297,dangling_wire_371,dangling_wire_372,dangling_wire_373,N__20649,dangling_wire_374,dangling_wire_375,dangling_wire_376,N__21546,dangling_wire_377}),
            .RCLKE(),
            .RCLK(N__54311),
            .RE(N__58560),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .WE(N__27757));
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged10_physical (
            .RDATA({dangling_wire_378,dangling_wire_379,buf_data_iac_3,dangling_wire_380,dangling_wire_381,dangling_wire_382,buf_data_vac_3,dangling_wire_383,dangling_wire_384,dangling_wire_385,buf_data_iac_2,dangling_wire_386,dangling_wire_387,dangling_wire_388,buf_data_vac_2,dangling_wire_389}),
            .RADDR({dangling_wire_390,N__39027,N__38928,N__38841,N__38244,N__55995,N__47589,N__38364,N__45063,N__36447,N__36189}),
            .WADDR({dangling_wire_391,N__29556,N__29667,N__29766,N__28713,N__28821,N__28932,N__29037,N__29145,N__29253,N__29364}),
            .MASK({dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407}),
            .WDATA({dangling_wire_408,dangling_wire_409,N__31050,dangling_wire_410,dangling_wire_411,dangling_wire_412,N__28371,dangling_wire_413,dangling_wire_414,dangling_wire_415,N__28179,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__27897,dangling_wire_419}),
            .RCLKE(),
            .RCLK(N__54325),
            .RE(N__58424),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .WE(N__27749));
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged3_physical (
            .RDATA({dangling_wire_420,dangling_wire_421,buf_data_iac_17,dangling_wire_422,dangling_wire_423,dangling_wire_424,buf_data_vac_17,dangling_wire_425,dangling_wire_426,dangling_wire_427,buf_data_iac_16,dangling_wire_428,dangling_wire_429,dangling_wire_430,buf_data_vac_16,dangling_wire_431}),
            .RADDR({dangling_wire_432,N__39009,N__38910,N__38823,N__38226,N__55977,N__47571,N__38346,N__45045,N__36429,N__36171}),
            .WADDR({dangling_wire_433,N__29538,N__29649,N__29748,N__28695,N__28803,N__28914,N__29019,N__29127,N__29235,N__29346}),
            .MASK({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449}),
            .WDATA({dangling_wire_450,dangling_wire_451,N__39768,dangling_wire_452,dangling_wire_453,dangling_wire_454,N__24393,dangling_wire_455,dangling_wire_456,dangling_wire_457,N__27348,dangling_wire_458,dangling_wire_459,dangling_wire_460,N__22683,dangling_wire_461}),
            .RCLKE(),
            .RCLK(N__54406),
            .RE(N__58509),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .WE(N__27729));
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged11_physical (
            .RDATA({dangling_wire_462,dangling_wire_463,buf_data_iac_1,dangling_wire_464,dangling_wire_465,dangling_wire_466,buf_data_vac_1,dangling_wire_467,dangling_wire_468,dangling_wire_469,buf_data_iac_0,dangling_wire_470,dangling_wire_471,dangling_wire_472,buf_data_vac_0,dangling_wire_473}),
            .RADDR({dangling_wire_474,N__39021,N__38922,N__38835,N__38238,N__55989,N__47583,N__38358,N__45057,N__36441,N__36183}),
            .WADDR({dangling_wire_475,N__29550,N__29661,N__29760,N__28707,N__28815,N__28926,N__29031,N__29139,N__29247,N__29358}),
            .MASK({dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .WDATA({dangling_wire_492,dangling_wire_493,N__32847,dangling_wire_494,dangling_wire_495,dangling_wire_496,N__33717,dangling_wire_497,dangling_wire_498,dangling_wire_499,N__26973,dangling_wire_500,dangling_wire_501,dangling_wire_502,N__26907,dangling_wire_503}),
            .RCLKE(),
            .RCLK(N__54351),
            .RE(N__58428),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .WE(N__27748));
    IO_PAD ipInertedIOPad_VAC_DRDY_iopad (
            .OE(N__59563),
            .DIN(N__59562),
            .DOUT(N__59561),
            .PACKAGEPIN(VAC_DRDY));
    defparam ipInertedIOPad_VAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_DRDY_preio (
            .PADOEN(N__59563),
            .PADOUT(N__59562),
            .PADIN(N__59561),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT1_iopad (
            .OE(N__59554),
            .DIN(N__59553),
            .DOUT(N__59552),
            .PACKAGEPIN(IAC_FLT1));
    defparam ipInertedIOPad_IAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT1_preio (
            .PADOEN(N__59554),
            .PADOUT(N__59553),
            .PADIN(N__59552),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44121),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK_iopad (
            .OE(N__59545),
            .DIN(N__59544),
            .DOUT(N__59543),
            .PACKAGEPIN(DDS_SCK));
    defparam ipInertedIOPad_DDS_SCK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK_preio (
            .PADOEN(N__59545),
            .PADOUT(N__59544),
            .PADIN(N__59543),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34197),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_166_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_166_iopad (
            .OE(N__59536),
            .DIN(N__59535),
            .DOUT(N__59534),
            .PACKAGEPIN(ICE_IOR_166));
    defparam ipInertedIOPad_ICE_IOR_166_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_166_preio (
            .PADOEN(N__59536),
            .PADOUT(N__59535),
            .PADIN(N__59534),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_119_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_119_iopad (
            .OE(N__59527),
            .DIN(N__59526),
            .DOUT(N__59525),
            .PACKAGEPIN(ICE_IOR_119));
    defparam ipInertedIOPad_ICE_IOR_119_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_119_preio (
            .PADOEN(N__59527),
            .PADOUT(N__59526),
            .PADIN(N__59525),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI_iopad (
            .OE(N__59518),
            .DIN(N__59517),
            .DOUT(N__59516),
            .PACKAGEPIN(DDS_MOSI));
    defparam ipInertedIOPad_DDS_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI_preio (
            .PADOEN(N__59518),
            .PADOUT(N__59517),
            .PADIN(N__59516),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36762),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MISO_iopad (
            .OE(N__59509),
            .DIN(N__59508),
            .DOUT(N__59507),
            .PACKAGEPIN(VAC_MISO));
    defparam ipInertedIOPad_VAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_MISO_preio (
            .PADOEN(N__59509),
            .PADOUT(N__59508),
            .PADIN(N__59507),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI1_iopad (
            .OE(N__59500),
            .DIN(N__59499),
            .DOUT(N__59498),
            .PACKAGEPIN(DDS_MOSI1));
    defparam ipInertedIOPad_DDS_MOSI1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI1_preio (
            .PADOEN(N__59500),
            .PADOUT(N__59499),
            .PADIN(N__59498),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24726),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_146_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_146_iopad (
            .OE(N__59491),
            .DIN(N__59490),
            .DOUT(N__59489),
            .PACKAGEPIN(ICE_IOR_146));
    defparam ipInertedIOPad_ICE_IOR_146_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_146_preio (
            .PADOEN(N__59491),
            .PADOUT(N__59490),
            .PADIN(N__59489),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_CLK_iopad (
            .OE(N__59482),
            .DIN(N__59481),
            .DOUT(N__59480),
            .PACKAGEPIN(VDC_CLK));
    defparam ipInertedIOPad_VDC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_CLK_preio (
            .PADOEN(N__59482),
            .PADOUT(N__59481),
            .PADIN(N__59480),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__53324),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_222_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_222_iopad (
            .OE(N__59473),
            .DIN(N__59472),
            .DOUT(N__59471),
            .PACKAGEPIN(ICE_IOT_222));
    defparam ipInertedIOPad_ICE_IOT_222_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_222_preio (
            .PADOEN(N__59473),
            .PADOUT(N__59472),
            .PADIN(N__59471),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CS_iopad (
            .OE(N__59464),
            .DIN(N__59463),
            .DOUT(N__59462),
            .PACKAGEPIN(IAC_CS));
    defparam ipInertedIOPad_IAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CS_preio (
            .PADOEN(N__59464),
            .PADOUT(N__59463),
            .PADIN(N__59462),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21213),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_18B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_18B_iopad (
            .OE(N__59455),
            .DIN(N__59454),
            .DOUT(N__59453),
            .PACKAGEPIN(ICE_IOL_18B));
    defparam ipInertedIOPad_ICE_IOL_18B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_18B_preio (
            .PADOEN(N__59455),
            .PADOUT(N__59454),
            .PADIN(N__59453),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13A_iopad (
            .OE(N__59446),
            .DIN(N__59445),
            .DOUT(N__59444),
            .PACKAGEPIN(ICE_IOL_13A));
    defparam ipInertedIOPad_ICE_IOL_13A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13A_preio (
            .PADOEN(N__59446),
            .PADOUT(N__59445),
            .PADIN(N__59444),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_81_iopad (
            .OE(N__59437),
            .DIN(N__59436),
            .DOUT(N__59435),
            .PACKAGEPIN(ICE_IOB_81));
    defparam ipInertedIOPad_ICE_IOB_81_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_81_preio (
            .PADOEN(N__59437),
            .PADOUT(N__59436),
            .PADIN(N__59435),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR1_iopad (
            .OE(N__59428),
            .DIN(N__59427),
            .DOUT(N__59426),
            .PACKAGEPIN(VAC_OSR1));
    defparam ipInertedIOPad_VAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR1_preio (
            .PADOEN(N__59428),
            .PADOUT(N__59427),
            .PADIN(N__59426),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23187),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MOSI_iopad (
            .OE(N__59419),
            .DIN(N__59418),
            .DOUT(N__59417),
            .PACKAGEPIN(IAC_MOSI));
    defparam ipInertedIOPad_IAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_MOSI_preio (
            .PADOEN(N__59419),
            .PADOUT(N__59418),
            .PADIN(N__59417),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS1_iopad (
            .OE(N__59410),
            .DIN(N__59409),
            .DOUT(N__59408),
            .PACKAGEPIN(DDS_CS1));
    defparam ipInertedIOPad_DDS_CS1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS1_preio (
            .PADOEN(N__59410),
            .PADOUT(N__59409),
            .PADIN(N__59408),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20304),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4B_iopad (
            .OE(N__59401),
            .DIN(N__59400),
            .DOUT(N__59399),
            .PACKAGEPIN(ICE_IOL_4B));
    defparam ipInertedIOPad_ICE_IOL_4B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4B_preio (
            .PADOEN(N__59401),
            .PADOUT(N__59400),
            .PADIN(N__59399),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_94_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_94_iopad (
            .OE(N__59392),
            .DIN(N__59391),
            .DOUT(N__59390),
            .PACKAGEPIN(ICE_IOB_94));
    defparam ipInertedIOPad_ICE_IOB_94_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_94_preio (
            .PADOEN(N__59392),
            .PADOUT(N__59391),
            .PADIN(N__59390),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CS_iopad (
            .OE(N__59383),
            .DIN(N__59382),
            .DOUT(N__59381),
            .PACKAGEPIN(VAC_CS));
    defparam ipInertedIOPad_VAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CS_preio (
            .PADOEN(N__59383),
            .PADOUT(N__59382),
            .PADIN(N__59381),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21126),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CLK_iopad (
            .OE(N__59374),
            .DIN(N__59373),
            .DOUT(N__59372),
            .PACKAGEPIN(VAC_CLK));
    defparam ipInertedIOPad_VAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CLK_preio (
            .PADOEN(N__59374),
            .PADOUT(N__59373),
            .PADIN(N__59372),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22998),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_CE0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_CE0_iopad (
            .OE(N__59365),
            .DIN(N__59364),
            .DOUT(N__59363),
            .PACKAGEPIN(ICE_SPI_CE0));
    defparam ipInertedIOPad_ICE_SPI_CE0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_CE0_preio (
            .PADOEN(N__59365),
            .PADOUT(N__59364),
            .PADIN(N__59363),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_CE0),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_167_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_167_iopad (
            .OE(N__59356),
            .DIN(N__59355),
            .DOUT(N__59354),
            .PACKAGEPIN(ICE_IOR_167));
    defparam ipInertedIOPad_ICE_IOR_167_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_167_preio (
            .PADOEN(N__59356),
            .PADOUT(N__59355),
            .PADIN(N__59354),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_118_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_118_iopad (
            .OE(N__59347),
            .DIN(N__59346),
            .DOUT(N__59345),
            .PACKAGEPIN(ICE_IOR_118));
    defparam ipInertedIOPad_ICE_IOR_118_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_118_preio (
            .PADOEN(N__59347),
            .PADOUT(N__59346),
            .PADIN(N__59345),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_SDO_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_SDO_iopad (
            .OE(N__59338),
            .DIN(N__59337),
            .DOUT(N__59336),
            .PACKAGEPIN(RTD_SDO));
    defparam ipInertedIOPad_RTD_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_SDO_preio (
            .PADOEN(N__59338),
            .PADOUT(N__59337),
            .PADIN(N__59336),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_SDO),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR0_iopad (
            .OE(N__59329),
            .DIN(N__59328),
            .DOUT(N__59327),
            .PACKAGEPIN(IAC_OSR0));
    defparam ipInertedIOPad_IAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR0_preio (
            .PADOEN(N__59329),
            .PADOUT(N__59328),
            .PADIN(N__59327),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27636),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SCLK_iopad (
            .OE(N__59320),
            .DIN(N__59319),
            .DOUT(N__59318),
            .PACKAGEPIN(VDC_SCLK));
    defparam ipInertedIOPad_VDC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_SCLK_preio (
            .PADOEN(N__59320),
            .PADOUT(N__59319),
            .PADIN(N__59318),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25851),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT1_iopad (
            .OE(N__59311),
            .DIN(N__59310),
            .DOUT(N__59309),
            .PACKAGEPIN(VAC_FLT1));
    defparam ipInertedIOPad_VAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT1_preio (
            .PADOEN(N__59311),
            .PADOUT(N__59310),
            .PADIN(N__59309),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25365),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_MOSI_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_MOSI_iopad (
            .OE(N__59302),
            .DIN(N__59301),
            .DOUT(N__59300),
            .PACKAGEPIN(ICE_SPI_MOSI));
    defparam ipInertedIOPad_ICE_SPI_MOSI_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_MOSI_preio (
            .PADOEN(N__59302),
            .PADOUT(N__59301),
            .PADIN(N__59300),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_MOSI),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_165_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_165_iopad (
            .OE(N__59293),
            .DIN(N__59292),
            .DOUT(N__59291),
            .PACKAGEPIN(ICE_IOR_165));
    defparam ipInertedIOPad_ICE_IOR_165_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_165_preio (
            .PADOEN(N__59293),
            .PADOUT(N__59292),
            .PADIN(N__59291),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_147_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_147_iopad (
            .OE(N__59284),
            .DIN(N__59283),
            .DOUT(N__59282),
            .PACKAGEPIN(ICE_IOR_147));
    defparam ipInertedIOPad_ICE_IOR_147_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_147_preio (
            .PADOEN(N__59284),
            .PADOUT(N__59283),
            .PADIN(N__59282),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_14A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_14A_iopad (
            .OE(N__59275),
            .DIN(N__59274),
            .DOUT(N__59273),
            .PACKAGEPIN(ICE_IOL_14A));
    defparam ipInertedIOPad_ICE_IOL_14A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_14A_preio (
            .PADOEN(N__59275),
            .PADOUT(N__59274),
            .PADIN(N__59273),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13B_iopad (
            .OE(N__59266),
            .DIN(N__59265),
            .DOUT(N__59264),
            .PACKAGEPIN(ICE_IOL_13B));
    defparam ipInertedIOPad_ICE_IOL_13B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13B_preio (
            .PADOEN(N__59266),
            .PADOUT(N__59265),
            .PADIN(N__59264),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_91_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_91_iopad (
            .OE(N__59257),
            .DIN(N__59256),
            .DOUT(N__59255),
            .PACKAGEPIN(ICE_IOB_91));
    defparam ipInertedIOPad_ICE_IOB_91_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_91_preio (
            .PADOEN(N__59257),
            .PADOUT(N__59256),
            .PADIN(N__59255),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_0_iopad (
            .OE(N__59248),
            .DIN(N__59247),
            .DOUT(N__59246),
            .PACKAGEPIN(ICE_GPMO_0));
    defparam ipInertedIOPad_ICE_GPMO_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_0_preio (
            .PADOEN(N__59248),
            .PADOUT(N__59247),
            .PADIN(N__59246),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_RNG_0_iopad (
            .OE(N__59239),
            .DIN(N__59238),
            .DOUT(N__59237),
            .PACKAGEPIN(DDS_RNG_0));
    defparam ipInertedIOPad_DDS_RNG_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_RNG_0_preio (
            .PADOEN(N__59239),
            .PADOUT(N__59238),
            .PADIN(N__59237),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36365),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_RNG0_iopad (
            .OE(N__59230),
            .DIN(N__59229),
            .DOUT(N__59228),
            .PACKAGEPIN(VDC_RNG0));
    defparam ipInertedIOPad_VDC_RNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_RNG0_preio (
            .PADOEN(N__59230),
            .PADOUT(N__59229),
            .PADIN(N__59228),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31866),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_SCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_SCLK_iopad (
            .OE(N__59221),
            .DIN(N__59220),
            .DOUT(N__59219),
            .PACKAGEPIN(ICE_SPI_SCLK));
    defparam ipInertedIOPad_ICE_SPI_SCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_SCLK_preio (
            .PADOEN(N__59221),
            .PADOUT(N__59220),
            .PADIN(N__59219),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_SCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_152_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_152_iopad (
            .OE(N__59212),
            .DIN(N__59211),
            .DOUT(N__59210),
            .PACKAGEPIN(ICE_IOR_152));
    defparam ipInertedIOPad_ICE_IOR_152_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_152_preio (
            .PADOEN(N__59212),
            .PADOUT(N__59211),
            .PADIN(N__59210),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12A_iopad (
            .OE(N__59203),
            .DIN(N__59202),
            .DOUT(N__59201),
            .PACKAGEPIN(ICE_IOL_12A));
    defparam ipInertedIOPad_ICE_IOL_12A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12A_preio (
            .PADOEN(N__59203),
            .PADOUT(N__59202),
            .PADIN(N__59201),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_DRDY_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_DRDY_iopad (
            .OE(N__59194),
            .DIN(N__59193),
            .DOUT(N__59192),
            .PACKAGEPIN(RTD_DRDY));
    defparam ipInertedIOPad_RTD_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_DRDY_preio (
            .PADOEN(N__59194),
            .PADOUT(N__59193),
            .PADIN(N__59192),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_SPI_MISO_iopad (
            .OE(N__59185),
            .DIN(N__59184),
            .DOUT(N__59183),
            .PACKAGEPIN(ICE_SPI_MISO));
    defparam ipInertedIOPad_ICE_SPI_MISO_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_SPI_MISO_preio (
            .PADOEN(N__59185),
            .PADOUT(N__59184),
            .PADIN(N__59183),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34143),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_177_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_177_iopad (
            .OE(N__59176),
            .DIN(N__59175),
            .DOUT(N__59174),
            .PACKAGEPIN(ICE_IOT_177));
    defparam ipInertedIOPad_ICE_IOT_177_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_177_preio (
            .PADOEN(N__59176),
            .PADOUT(N__59175),
            .PADIN(N__59174),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_141_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_141_iopad (
            .OE(N__59167),
            .DIN(N__59166),
            .DOUT(N__59165),
            .PACKAGEPIN(ICE_IOR_141));
    defparam ipInertedIOPad_ICE_IOR_141_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_141_preio (
            .PADOEN(N__59167),
            .PADOUT(N__59166),
            .PADIN(N__59165),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_80_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_80_iopad (
            .OE(N__59158),
            .DIN(N__59157),
            .DOUT(N__59156),
            .PACKAGEPIN(ICE_IOB_80));
    defparam ipInertedIOPad_ICE_IOB_80_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_80_preio (
            .PADOEN(N__59158),
            .PADOUT(N__59157),
            .PADIN(N__59156),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_102_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_102_iopad (
            .OE(N__59149),
            .DIN(N__59148),
            .DOUT(N__59147),
            .PACKAGEPIN(ICE_IOB_102));
    defparam ipInertedIOPad_ICE_IOB_102_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_102_preio (
            .PADOEN(N__59149),
            .PADOUT(N__59148),
            .PADIN(N__59147),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_2_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_2_iopad (
            .OE(N__59140),
            .DIN(N__59139),
            .DOUT(N__59138),
            .PACKAGEPIN(ICE_GPMO_2));
    defparam ipInertedIOPad_ICE_GPMO_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_2_preio (
            .PADOEN(N__59140),
            .PADOUT(N__59139),
            .PADIN(N__59138),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_2),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_GPMI_0_iopad (
            .OE(N__59131),
            .DIN(N__59130),
            .DOUT(N__59129),
            .PACKAGEPIN(ICE_GPMI_0));
    defparam ipInertedIOPad_ICE_GPMI_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_GPMI_0_preio (
            .PADOEN(N__59131),
            .PADOUT(N__59130),
            .PADIN(N__59129),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__35928),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MISO_iopad (
            .OE(N__59122),
            .DIN(N__59121),
            .DOUT(N__59120),
            .PACKAGEPIN(IAC_MISO));
    defparam ipInertedIOPad_IAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_MISO_preio (
            .PADOEN(N__59122),
            .PADOUT(N__59121),
            .PADIN(N__59120),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR0_iopad (
            .OE(N__59113),
            .DIN(N__59112),
            .DOUT(N__59111),
            .PACKAGEPIN(VAC_OSR0));
    defparam ipInertedIOPad_VAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR0_preio (
            .PADOEN(N__59113),
            .PADOUT(N__59112),
            .PADIN(N__59111),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__41400),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MOSI_iopad (
            .OE(N__59104),
            .DIN(N__59103),
            .DOUT(N__59102),
            .PACKAGEPIN(VAC_MOSI));
    defparam ipInertedIOPad_VAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_MOSI_preio (
            .PADOEN(N__59104),
            .PADOUT(N__59103),
            .PADIN(N__59102),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TEST_LED_iopad (
            .OE(N__59095),
            .DIN(N__59094),
            .DOUT(N__59093),
            .PACKAGEPIN(TEST_LED));
    defparam ipInertedIOPad_TEST_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_TEST_LED_preio (
            .PADOEN(N__59095),
            .PADOUT(N__59094),
            .PADIN(N__59093),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__39207),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_148_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_148_iopad (
            .OE(N__59086),
            .DIN(N__59085),
            .DOUT(N__59084),
            .PACKAGEPIN(ICE_IOR_148));
    defparam ipInertedIOPad_ICE_IOR_148_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_148_preio (
            .PADOEN(N__59086),
            .PADOUT(N__59085),
            .PADIN(N__59084),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_STAT_COMM_iopad (
            .OE(N__59077),
            .DIN(N__59076),
            .DOUT(N__59075),
            .PACKAGEPIN(STAT_COMM));
    defparam ipInertedIOPad_STAT_COMM_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_STAT_COMM_preio (
            .PADOEN(N__59077),
            .PADOUT(N__59076),
            .PADIN(N__59075),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19191),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SYSCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SYSCLK_iopad (
            .OE(N__59068),
            .DIN(N__59067),
            .DOUT(N__59066),
            .PACKAGEPIN(ICE_SYSCLK));
    defparam ipInertedIOPad_ICE_SYSCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SYSCLK_preio (
            .PADOEN(N__59068),
            .PADOUT(N__59067),
            .PADIN(N__59066),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SYSCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_161_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_161_iopad (
            .OE(N__59059),
            .DIN(N__59058),
            .DOUT(N__59057),
            .PACKAGEPIN(ICE_IOR_161));
    defparam ipInertedIOPad_ICE_IOR_161_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_161_preio (
            .PADOEN(N__59059),
            .PADOUT(N__59058),
            .PADIN(N__59057),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_95_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_95_iopad (
            .OE(N__59050),
            .DIN(N__59049),
            .DOUT(N__59048),
            .PACKAGEPIN(ICE_IOB_95));
    defparam ipInertedIOPad_ICE_IOB_95_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_95_preio (
            .PADOEN(N__59050),
            .PADOUT(N__59049),
            .PADIN(N__59048),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_82_iopad (
            .OE(N__59041),
            .DIN(N__59040),
            .DOUT(N__59039),
            .PACKAGEPIN(ICE_IOB_82));
    defparam ipInertedIOPad_ICE_IOB_82_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_82_preio (
            .PADOEN(N__59041),
            .PADOUT(N__59040),
            .PADIN(N__59039),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_104_iopad (
            .OE(N__59032),
            .DIN(N__59031),
            .DOUT(N__59030),
            .PACKAGEPIN(ICE_IOB_104));
    defparam ipInertedIOPad_ICE_IOB_104_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_104_preio (
            .PADOEN(N__59032),
            .PADOUT(N__59031),
            .PADIN(N__59030),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CLK_iopad (
            .OE(N__59023),
            .DIN(N__59022),
            .DOUT(N__59021),
            .PACKAGEPIN(IAC_CLK));
    defparam ipInertedIOPad_IAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CLK_preio (
            .PADOEN(N__59023),
            .PADOUT(N__59022),
            .PADIN(N__59021),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22994),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS_iopad (
            .OE(N__59014),
            .DIN(N__59013),
            .DOUT(N__59012),
            .PACKAGEPIN(DDS_CS));
    defparam ipInertedIOPad_DDS_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS_preio (
            .PADOEN(N__59014),
            .PADOUT(N__59013),
            .PADIN(N__59012),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36741),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG0_iopad (
            .OE(N__59005),
            .DIN(N__59004),
            .DOUT(N__59003),
            .PACKAGEPIN(SELIRNG0));
    defparam ipInertedIOPad_SELIRNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG0_preio (
            .PADOEN(N__59005),
            .PADOUT(N__59004),
            .PADIN(N__59003),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31782),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SDI_iopad (
            .OE(N__58996),
            .DIN(N__58995),
            .DOUT(N__58994),
            .PACKAGEPIN(RTD_SDI));
    defparam ipInertedIOPad_RTD_SDI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SDI_preio (
            .PADOEN(N__58996),
            .PADOUT(N__58995),
            .PADIN(N__58994),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19254),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_221_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_221_iopad (
            .OE(N__58987),
            .DIN(N__58986),
            .DOUT(N__58985),
            .PACKAGEPIN(ICE_IOT_221));
    defparam ipInertedIOPad_ICE_IOT_221_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_221_preio (
            .PADOEN(N__58987),
            .PADOUT(N__58986),
            .PADIN(N__58985),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_197_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_197_iopad (
            .OE(N__58978),
            .DIN(N__58977),
            .DOUT(N__58976),
            .PACKAGEPIN(ICE_IOT_197));
    defparam ipInertedIOPad_ICE_IOT_197_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_197_preio (
            .PADOEN(N__58978),
            .PADOUT(N__58977),
            .PADIN(N__58976),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK_iopad (
            .OE(N__58969),
            .DIN(N__58968),
            .DOUT(N__58967),
            .PACKAGEPIN(DDS_MCLK));
    defparam ipInertedIOPad_DDS_MCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK_preio (
            .PADOEN(N__58969),
            .PADOUT(N__58968),
            .PADIN(N__58967),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__38649),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SCLK_iopad (
            .OE(N__58960),
            .DIN(N__58959),
            .DOUT(N__58958),
            .PACKAGEPIN(RTD_SCLK));
    defparam ipInertedIOPad_RTD_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SCLK_preio (
            .PADOEN(N__58960),
            .PADOUT(N__58959),
            .PADIN(N__58958),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19224),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_CS_iopad (
            .OE(N__58951),
            .DIN(N__58950),
            .DOUT(N__58949),
            .PACKAGEPIN(RTD_CS));
    defparam ipInertedIOPad_RTD_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_CS_preio (
            .PADOEN(N__58951),
            .PADOUT(N__58950),
            .PADIN(N__58949),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19581),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_137_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_137_iopad (
            .OE(N__58942),
            .DIN(N__58941),
            .DOUT(N__58940),
            .PACKAGEPIN(ICE_IOR_137));
    defparam ipInertedIOPad_ICE_IOR_137_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_137_preio (
            .PADOEN(N__58942),
            .PADOUT(N__58941),
            .PADIN(N__58940),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR1_iopad (
            .OE(N__58933),
            .DIN(N__58932),
            .DOUT(N__58931),
            .PACKAGEPIN(IAC_OSR1));
    defparam ipInertedIOPad_IAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR1_preio (
            .PADOEN(N__58933),
            .PADOUT(N__58932),
            .PADIN(N__58931),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__39807),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT0_iopad (
            .OE(N__58924),
            .DIN(N__58923),
            .DOUT(N__58922),
            .PACKAGEPIN(VAC_FLT0));
    defparam ipInertedIOPad_VAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT0_preio (
            .PADOEN(N__58924),
            .PADOUT(N__58923),
            .PADIN(N__58922),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31902),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_144_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_144_iopad (
            .OE(N__58915),
            .DIN(N__58914),
            .DOUT(N__58913),
            .PACKAGEPIN(ICE_IOR_144));
    defparam ipInertedIOPad_ICE_IOR_144_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_144_preio (
            .PADOEN(N__58915),
            .PADOUT(N__58914),
            .PADIN(N__58913),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_128_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_128_iopad (
            .OE(N__58906),
            .DIN(N__58905),
            .DOUT(N__58904),
            .PACKAGEPIN(ICE_IOR_128));
    defparam ipInertedIOPad_ICE_IOR_128_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_128_preio (
            .PADOEN(N__58906),
            .PADOUT(N__58905),
            .PADIN(N__58904),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_1_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_1_iopad (
            .OE(N__58897),
            .DIN(N__58896),
            .DOUT(N__58895),
            .PACKAGEPIN(ICE_GPMO_1));
    defparam ipInertedIOPad_ICE_GPMO_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_1_preio (
            .PADOEN(N__58897),
            .PADOUT(N__58896),
            .PADIN(N__58895),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_SCLK_iopad (
            .OE(N__58888),
            .DIN(N__58887),
            .DOUT(N__58886),
            .PACKAGEPIN(IAC_SCLK));
    defparam ipInertedIOPad_IAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_SCLK_preio (
            .PADOEN(N__58888),
            .PADOUT(N__58887),
            .PADIN(N__58886),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23322),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_EIS_SYNCCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_EIS_SYNCCLK_iopad (
            .OE(N__58879),
            .DIN(N__58878),
            .DOUT(N__58877),
            .PACKAGEPIN(EIS_SYNCCLK));
    defparam ipInertedIOPad_EIS_SYNCCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_EIS_SYNCCLK_preio (
            .PADOEN(N__58879),
            .PADOUT(N__58878),
            .PADIN(N__58877),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(EIS_SYNCCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_139_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_139_iopad (
            .OE(N__58870),
            .DIN(N__58869),
            .DOUT(N__58868),
            .PACKAGEPIN(ICE_IOR_139));
    defparam ipInertedIOPad_ICE_IOR_139_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_139_preio (
            .PADOEN(N__58870),
            .PADOUT(N__58869),
            .PADIN(N__58868),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4A_iopad (
            .OE(N__58861),
            .DIN(N__58860),
            .DOUT(N__58859),
            .PACKAGEPIN(ICE_IOL_4A));
    defparam ipInertedIOPad_ICE_IOL_4A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4A_preio (
            .PADOEN(N__58861),
            .PADOUT(N__58860),
            .PADIN(N__58859),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_SCLK_iopad (
            .OE(N__58852),
            .DIN(N__58851),
            .DOUT(N__58850),
            .PACKAGEPIN(VAC_SCLK));
    defparam ipInertedIOPad_VAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_SCLK_preio (
            .PADOEN(N__58852),
            .PADOUT(N__58851),
            .PADIN(N__58850),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21957),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_THERMOSTAT_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_THERMOSTAT_iopad (
            .OE(N__58843),
            .DIN(N__58842),
            .DOUT(N__58841),
            .PACKAGEPIN(THERMOSTAT));
    defparam ipInertedIOPad_THERMOSTAT_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_THERMOSTAT_preio (
            .PADOEN(N__58843),
            .PADOUT(N__58842),
            .PADIN(N__58841),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(THERMOSTAT),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_164_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_164_iopad (
            .OE(N__58834),
            .DIN(N__58833),
            .DOUT(N__58832),
            .PACKAGEPIN(ICE_IOR_164));
    defparam ipInertedIOPad_ICE_IOR_164_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_164_preio (
            .PADOEN(N__58834),
            .PADOUT(N__58833),
            .PADIN(N__58832),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_103_iopad (
            .OE(N__58825),
            .DIN(N__58824),
            .DOUT(N__58823),
            .PACKAGEPIN(ICE_IOB_103));
    defparam ipInertedIOPad_ICE_IOB_103_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_103_preio (
            .PADOEN(N__58825),
            .PADOUT(N__58824),
            .PADIN(N__58823),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AMPV_POW_iopad (
            .OE(N__58816),
            .DIN(N__58815),
            .DOUT(N__58814),
            .PACKAGEPIN(AMPV_POW));
    defparam ipInertedIOPad_AMPV_POW_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AMPV_POW_preio (
            .PADOEN(N__58816),
            .PADOUT(N__58815),
            .PADIN(N__58814),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23058),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SDO_iopad (
            .OE(N__58807),
            .DIN(N__58806),
            .DOUT(N__58805),
            .PACKAGEPIN(VDC_SDO));
    defparam ipInertedIOPad_VDC_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDC_SDO_preio (
            .PADOEN(N__58807),
            .PADOUT(N__58806),
            .PADIN(N__58805),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VDC_SDO),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_174_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_174_iopad (
            .OE(N__58798),
            .DIN(N__58797),
            .DOUT(N__58796),
            .PACKAGEPIN(ICE_IOT_174));
    defparam ipInertedIOPad_ICE_IOT_174_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_174_preio (
            .PADOEN(N__58798),
            .PADOUT(N__58797),
            .PADIN(N__58796),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_140_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_140_iopad (
            .OE(N__58789),
            .DIN(N__58788),
            .DOUT(N__58787),
            .PACKAGEPIN(ICE_IOR_140));
    defparam ipInertedIOPad_ICE_IOR_140_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_140_preio (
            .PADOEN(N__58789),
            .PADOUT(N__58788),
            .PADIN(N__58787),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_96_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_96_iopad (
            .OE(N__58780),
            .DIN(N__58779),
            .DOUT(N__58778),
            .PACKAGEPIN(ICE_IOB_96));
    defparam ipInertedIOPad_ICE_IOB_96_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_96_preio (
            .PADOEN(N__58780),
            .PADOUT(N__58779),
            .PADIN(N__58778),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_CONT_SD_iopad (
            .OE(N__58771),
            .DIN(N__58770),
            .DOUT(N__58769),
            .PACKAGEPIN(CONT_SD));
    defparam ipInertedIOPad_CONT_SD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_CONT_SD_preio (
            .PADOEN(N__58771),
            .PADOUT(N__58770),
            .PADIN(N__58769),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44592),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AC_ADC_SYNC_iopad (
            .OE(N__58762),
            .DIN(N__58761),
            .DOUT(N__58760),
            .PACKAGEPIN(AC_ADC_SYNC));
    defparam ipInertedIOPad_AC_ADC_SYNC_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AC_ADC_SYNC_preio (
            .PADOEN(N__58762),
            .PADOUT(N__58761),
            .PADIN(N__58760),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21282),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG1_iopad (
            .OE(N__58753),
            .DIN(N__58752),
            .DOUT(N__58751),
            .PACKAGEPIN(SELIRNG1));
    defparam ipInertedIOPad_SELIRNG1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG1_preio (
            .PADOEN(N__58753),
            .PADOUT(N__58752),
            .PADIN(N__58751),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__41964),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12B_iopad (
            .OE(N__58744),
            .DIN(N__58743),
            .DOUT(N__58742),
            .PACKAGEPIN(ICE_IOL_12B));
    defparam ipInertedIOPad_ICE_IOL_12B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12B_preio (
            .PADOEN(N__58744),
            .PADOUT(N__58743),
            .PADIN(N__58742),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_160_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_160_iopad (
            .OE(N__58735),
            .DIN(N__58734),
            .DOUT(N__58733),
            .PACKAGEPIN(ICE_IOR_160));
    defparam ipInertedIOPad_ICE_IOR_160_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_160_preio (
            .PADOEN(N__58735),
            .PADOUT(N__58734),
            .PADIN(N__58733),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_136_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_136_iopad (
            .OE(N__58726),
            .DIN(N__58725),
            .DOUT(N__58724),
            .PACKAGEPIN(ICE_IOR_136));
    defparam ipInertedIOPad_ICE_IOR_136_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_136_preio (
            .PADOEN(N__58726),
            .PADOUT(N__58725),
            .PADIN(N__58724),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK1_iopad (
            .OE(N__58717),
            .DIN(N__58716),
            .DOUT(N__58715),
            .PACKAGEPIN(DDS_MCLK1));
    defparam ipInertedIOPad_DDS_MCLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK1_preio (
            .PADOEN(N__58717),
            .PADOUT(N__58716),
            .PADIN(N__58715),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19596),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_198_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_198_iopad (
            .OE(N__58708),
            .DIN(N__58707),
            .DOUT(N__58706),
            .PACKAGEPIN(ICE_IOT_198));
    defparam ipInertedIOPad_ICE_IOT_198_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_198_preio (
            .PADOEN(N__58708),
            .PADOUT(N__58707),
            .PADIN(N__58706),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_173_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_173_iopad (
            .OE(N__58699),
            .DIN(N__58698),
            .DOUT(N__58697),
            .PACKAGEPIN(ICE_IOT_173));
    defparam ipInertedIOPad_ICE_IOT_173_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_173_preio (
            .PADOEN(N__58699),
            .PADOUT(N__58698),
            .PADIN(N__58697),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_DRDY_iopad (
            .OE(N__58690),
            .DIN(N__58689),
            .DOUT(N__58688),
            .PACKAGEPIN(IAC_DRDY));
    defparam ipInertedIOPad_IAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_DRDY_preio (
            .PADOEN(N__58690),
            .PADOUT(N__58689),
            .PADIN(N__58688),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_DRDY),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_178_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_178_iopad (
            .OE(N__58681),
            .DIN(N__58680),
            .DOUT(N__58679),
            .PACKAGEPIN(ICE_IOT_178));
    defparam ipInertedIOPad_ICE_IOT_178_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_178_preio (
            .PADOEN(N__58681),
            .PADOUT(N__58680),
            .PADIN(N__58679),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_138_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_138_iopad (
            .OE(N__58672),
            .DIN(N__58671),
            .DOUT(N__58670),
            .PACKAGEPIN(ICE_IOR_138));
    defparam ipInertedIOPad_ICE_IOR_138_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_138_preio (
            .PADOEN(N__58672),
            .PADOUT(N__58671),
            .PADIN(N__58670),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_120_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_120_iopad (
            .OE(N__58663),
            .DIN(N__58662),
            .DOUT(N__58661),
            .PACKAGEPIN(ICE_IOR_120));
    defparam ipInertedIOPad_ICE_IOR_120_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_120_preio (
            .PADOEN(N__58663),
            .PADOUT(N__58662),
            .PADIN(N__58661),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT0_iopad (
            .OE(N__58654),
            .DIN(N__58653),
            .DOUT(N__58652),
            .PACKAGEPIN(IAC_FLT0));
    defparam ipInertedIOPad_IAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT0_preio (
            .PADOEN(N__58654),
            .PADOUT(N__58653),
            .PADIN(N__58652),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44685),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK1_iopad (
            .OE(N__58645),
            .DIN(N__58644),
            .DOUT(N__58643),
            .PACKAGEPIN(DDS_SCK1));
    defparam ipInertedIOPad_DDS_SCK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK1_preio (
            .PADOEN(N__58645),
            .PADOUT(N__58644),
            .PADIN(N__58643),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27132),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__14719 (
            .O(N__58626),
            .I(\ADC_VDC.genclk.n19737 ));
    CascadeMux I__14718 (
            .O(N__58623),
            .I(N__58617));
    CascadeMux I__14717 (
            .O(N__58622),
            .I(N__58613));
    CascadeMux I__14716 (
            .O(N__58621),
            .I(N__58609));
    InMux I__14715 (
            .O(N__58620),
            .I(N__58592));
    InMux I__14714 (
            .O(N__58617),
            .I(N__58592));
    InMux I__14713 (
            .O(N__58616),
            .I(N__58592));
    InMux I__14712 (
            .O(N__58613),
            .I(N__58592));
    InMux I__14711 (
            .O(N__58612),
            .I(N__58592));
    InMux I__14710 (
            .O(N__58609),
            .I(N__58592));
    InMux I__14709 (
            .O(N__58608),
            .I(N__58592));
    SRMux I__14708 (
            .O(N__58607),
            .I(N__58589));
    LocalMux I__14707 (
            .O(N__58592),
            .I(N__58586));
    LocalMux I__14706 (
            .O(N__58589),
            .I(N__58581));
    Span4Mux_v I__14705 (
            .O(N__58586),
            .I(N__58570));
    SRMux I__14704 (
            .O(N__58585),
            .I(N__58567));
    SRMux I__14703 (
            .O(N__58584),
            .I(N__58561));
    Span4Mux_h I__14702 (
            .O(N__58581),
            .I(N__58557));
    CascadeMux I__14701 (
            .O(N__58580),
            .I(N__58554));
    CascadeMux I__14700 (
            .O(N__58579),
            .I(N__58550));
    CascadeMux I__14699 (
            .O(N__58578),
            .I(N__58546));
    CascadeMux I__14698 (
            .O(N__58577),
            .I(N__58542));
    CascadeMux I__14697 (
            .O(N__58576),
            .I(N__58538));
    CascadeMux I__14696 (
            .O(N__58575),
            .I(N__58534));
    CascadeMux I__14695 (
            .O(N__58574),
            .I(N__58530));
    CascadeMux I__14694 (
            .O(N__58573),
            .I(N__58526));
    Span4Mux_h I__14693 (
            .O(N__58570),
            .I(N__58519));
    LocalMux I__14692 (
            .O(N__58567),
            .I(N__58516));
    SRMux I__14691 (
            .O(N__58566),
            .I(N__58513));
    SRMux I__14690 (
            .O(N__58565),
            .I(N__58510));
    IoInMux I__14689 (
            .O(N__58564),
            .I(N__58504));
    LocalMux I__14688 (
            .O(N__58561),
            .I(N__58497));
    SRMux I__14687 (
            .O(N__58560),
            .I(N__58494));
    Span4Mux_v I__14686 (
            .O(N__58557),
            .I(N__58491));
    InMux I__14685 (
            .O(N__58554),
            .I(N__58476));
    InMux I__14684 (
            .O(N__58553),
            .I(N__58476));
    InMux I__14683 (
            .O(N__58550),
            .I(N__58476));
    InMux I__14682 (
            .O(N__58549),
            .I(N__58476));
    InMux I__14681 (
            .O(N__58546),
            .I(N__58476));
    InMux I__14680 (
            .O(N__58545),
            .I(N__58476));
    InMux I__14679 (
            .O(N__58542),
            .I(N__58476));
    InMux I__14678 (
            .O(N__58541),
            .I(N__58459));
    InMux I__14677 (
            .O(N__58538),
            .I(N__58459));
    InMux I__14676 (
            .O(N__58537),
            .I(N__58459));
    InMux I__14675 (
            .O(N__58534),
            .I(N__58459));
    InMux I__14674 (
            .O(N__58533),
            .I(N__58459));
    InMux I__14673 (
            .O(N__58530),
            .I(N__58459));
    InMux I__14672 (
            .O(N__58529),
            .I(N__58459));
    InMux I__14671 (
            .O(N__58526),
            .I(N__58459));
    CascadeMux I__14670 (
            .O(N__58525),
            .I(N__58456));
    CascadeMux I__14669 (
            .O(N__58524),
            .I(N__58452));
    CascadeMux I__14668 (
            .O(N__58523),
            .I(N__58448));
    CascadeMux I__14667 (
            .O(N__58522),
            .I(N__58444));
    Span4Mux_h I__14666 (
            .O(N__58519),
            .I(N__58435));
    Span4Mux_v I__14665 (
            .O(N__58516),
            .I(N__58435));
    LocalMux I__14664 (
            .O(N__58513),
            .I(N__58435));
    LocalMux I__14663 (
            .O(N__58510),
            .I(N__58435));
    SRMux I__14662 (
            .O(N__58509),
            .I(N__58432));
    SRMux I__14661 (
            .O(N__58508),
            .I(N__58429));
    SRMux I__14660 (
            .O(N__58507),
            .I(N__58425));
    LocalMux I__14659 (
            .O(N__58504),
            .I(N__58421));
    CascadeMux I__14658 (
            .O(N__58503),
            .I(N__58417));
    CascadeMux I__14657 (
            .O(N__58502),
            .I(N__58413));
    CascadeMux I__14656 (
            .O(N__58501),
            .I(N__58409));
    CascadeMux I__14655 (
            .O(N__58500),
            .I(N__58405));
    Span4Mux_h I__14654 (
            .O(N__58497),
            .I(N__58400));
    LocalMux I__14653 (
            .O(N__58494),
            .I(N__58400));
    Span4Mux_v I__14652 (
            .O(N__58491),
            .I(N__58397));
    LocalMux I__14651 (
            .O(N__58476),
            .I(N__58394));
    LocalMux I__14650 (
            .O(N__58459),
            .I(N__58391));
    InMux I__14649 (
            .O(N__58456),
            .I(N__58376));
    InMux I__14648 (
            .O(N__58455),
            .I(N__58376));
    InMux I__14647 (
            .O(N__58452),
            .I(N__58376));
    InMux I__14646 (
            .O(N__58451),
            .I(N__58376));
    InMux I__14645 (
            .O(N__58448),
            .I(N__58376));
    InMux I__14644 (
            .O(N__58447),
            .I(N__58376));
    InMux I__14643 (
            .O(N__58444),
            .I(N__58376));
    Span4Mux_v I__14642 (
            .O(N__58435),
            .I(N__58369));
    LocalMux I__14641 (
            .O(N__58432),
            .I(N__58369));
    LocalMux I__14640 (
            .O(N__58429),
            .I(N__58369));
    SRMux I__14639 (
            .O(N__58428),
            .I(N__58366));
    LocalMux I__14638 (
            .O(N__58425),
            .I(N__58363));
    SRMux I__14637 (
            .O(N__58424),
            .I(N__58360));
    IoSpan4Mux I__14636 (
            .O(N__58421),
            .I(N__58356));
    InMux I__14635 (
            .O(N__58420),
            .I(N__58339));
    InMux I__14634 (
            .O(N__58417),
            .I(N__58339));
    InMux I__14633 (
            .O(N__58416),
            .I(N__58339));
    InMux I__14632 (
            .O(N__58413),
            .I(N__58339));
    InMux I__14631 (
            .O(N__58412),
            .I(N__58339));
    InMux I__14630 (
            .O(N__58409),
            .I(N__58339));
    InMux I__14629 (
            .O(N__58408),
            .I(N__58339));
    InMux I__14628 (
            .O(N__58405),
            .I(N__58339));
    Span4Mux_v I__14627 (
            .O(N__58400),
            .I(N__58336));
    Span4Mux_v I__14626 (
            .O(N__58397),
            .I(N__58326));
    Span4Mux_h I__14625 (
            .O(N__58394),
            .I(N__58326));
    Span4Mux_v I__14624 (
            .O(N__58391),
            .I(N__58326));
    LocalMux I__14623 (
            .O(N__58376),
            .I(N__58326));
    Span4Mux_v I__14622 (
            .O(N__58369),
            .I(N__58317));
    LocalMux I__14621 (
            .O(N__58366),
            .I(N__58317));
    Span4Mux_v I__14620 (
            .O(N__58363),
            .I(N__58317));
    LocalMux I__14619 (
            .O(N__58360),
            .I(N__58317));
    SRMux I__14618 (
            .O(N__58359),
            .I(N__58314));
    Span4Mux_s0_v I__14617 (
            .O(N__58356),
            .I(N__58311));
    LocalMux I__14616 (
            .O(N__58339),
            .I(N__58308));
    Sp12to4 I__14615 (
            .O(N__58336),
            .I(N__58305));
    InMux I__14614 (
            .O(N__58335),
            .I(N__58302));
    Span4Mux_v I__14613 (
            .O(N__58326),
            .I(N__58299));
    Span4Mux_v I__14612 (
            .O(N__58317),
            .I(N__58294));
    LocalMux I__14611 (
            .O(N__58314),
            .I(N__58294));
    Sp12to4 I__14610 (
            .O(N__58311),
            .I(N__58288));
    Span12Mux_s10_h I__14609 (
            .O(N__58308),
            .I(N__58288));
    Span12Mux_h I__14608 (
            .O(N__58305),
            .I(N__58283));
    LocalMux I__14607 (
            .O(N__58302),
            .I(N__58283));
    Sp12to4 I__14606 (
            .O(N__58299),
            .I(N__58278));
    Sp12to4 I__14605 (
            .O(N__58294),
            .I(N__58278));
    InMux I__14604 (
            .O(N__58293),
            .I(N__58275));
    Odrv12 I__14603 (
            .O(N__58288),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__14602 (
            .O(N__58283),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__14601 (
            .O(N__58278),
            .I(CONSTANT_ONE_NET));
    LocalMux I__14600 (
            .O(N__58275),
            .I(CONSTANT_ONE_NET));
    InMux I__14599 (
            .O(N__58266),
            .I(\ADC_VDC.genclk.n19738 ));
    SRMux I__14598 (
            .O(N__58263),
            .I(N__58260));
    LocalMux I__14597 (
            .O(N__58260),
            .I(N__58255));
    SRMux I__14596 (
            .O(N__58259),
            .I(N__58252));
    SRMux I__14595 (
            .O(N__58258),
            .I(N__58249));
    Span4Mux_v I__14594 (
            .O(N__58255),
            .I(N__58244));
    LocalMux I__14593 (
            .O(N__58252),
            .I(N__58244));
    LocalMux I__14592 (
            .O(N__58249),
            .I(N__58240));
    Span4Mux_h I__14591 (
            .O(N__58244),
            .I(N__58237));
    SRMux I__14590 (
            .O(N__58243),
            .I(N__58234));
    Span4Mux_v I__14589 (
            .O(N__58240),
            .I(N__58231));
    Sp12to4 I__14588 (
            .O(N__58237),
            .I(N__58226));
    LocalMux I__14587 (
            .O(N__58234),
            .I(N__58226));
    Odrv4 I__14586 (
            .O(N__58231),
            .I(\ADC_VDC.genclk.n15051 ));
    Odrv12 I__14585 (
            .O(N__58226),
            .I(\ADC_VDC.genclk.n15051 ));
    CascadeMux I__14584 (
            .O(N__58221),
            .I(N__58218));
    InMux I__14583 (
            .O(N__58218),
            .I(N__58214));
    InMux I__14582 (
            .O(N__58217),
            .I(N__58211));
    LocalMux I__14581 (
            .O(N__58214),
            .I(\ADC_VDC.genclk.t0on_6 ));
    LocalMux I__14580 (
            .O(N__58211),
            .I(\ADC_VDC.genclk.t0on_6 ));
    InMux I__14579 (
            .O(N__58206),
            .I(N__58202));
    InMux I__14578 (
            .O(N__58205),
            .I(N__58199));
    LocalMux I__14577 (
            .O(N__58202),
            .I(\ADC_VDC.genclk.t0on_1 ));
    LocalMux I__14576 (
            .O(N__58199),
            .I(\ADC_VDC.genclk.t0on_1 ));
    CascadeMux I__14575 (
            .O(N__58194),
            .I(N__58190));
    CascadeMux I__14574 (
            .O(N__58193),
            .I(N__58187));
    InMux I__14573 (
            .O(N__58190),
            .I(N__58184));
    InMux I__14572 (
            .O(N__58187),
            .I(N__58181));
    LocalMux I__14571 (
            .O(N__58184),
            .I(\ADC_VDC.genclk.t0on_4 ));
    LocalMux I__14570 (
            .O(N__58181),
            .I(\ADC_VDC.genclk.t0on_4 ));
    InMux I__14569 (
            .O(N__58176),
            .I(N__58172));
    InMux I__14568 (
            .O(N__58175),
            .I(N__58169));
    LocalMux I__14567 (
            .O(N__58172),
            .I(\ADC_VDC.genclk.t0on_0 ));
    LocalMux I__14566 (
            .O(N__58169),
            .I(\ADC_VDC.genclk.t0on_0 ));
    CascadeMux I__14565 (
            .O(N__58164),
            .I(\ADC_VDC.genclk.n21449_cascade_ ));
    CascadeMux I__14564 (
            .O(N__58161),
            .I(N__58157));
    CascadeMux I__14563 (
            .O(N__58160),
            .I(N__58154));
    InMux I__14562 (
            .O(N__58157),
            .I(N__58151));
    InMux I__14561 (
            .O(N__58154),
            .I(N__58148));
    LocalMux I__14560 (
            .O(N__58151),
            .I(N__58145));
    LocalMux I__14559 (
            .O(N__58148),
            .I(N__58142));
    Span4Mux_h I__14558 (
            .O(N__58145),
            .I(N__58139));
    Span4Mux_h I__14557 (
            .O(N__58142),
            .I(N__58136));
    Odrv4 I__14556 (
            .O(N__58139),
            .I(\ADC_VDC.genclk.n21443 ));
    Odrv4 I__14555 (
            .O(N__58136),
            .I(\ADC_VDC.genclk.n21443 ));
    InMux I__14554 (
            .O(N__58131),
            .I(N__58127));
    InMux I__14553 (
            .O(N__58130),
            .I(N__58124));
    LocalMux I__14552 (
            .O(N__58127),
            .I(\ADC_VDC.genclk.t0on_12 ));
    LocalMux I__14551 (
            .O(N__58124),
            .I(\ADC_VDC.genclk.t0on_12 ));
    CascadeMux I__14550 (
            .O(N__58119),
            .I(N__58116));
    InMux I__14549 (
            .O(N__58116),
            .I(N__58112));
    InMux I__14548 (
            .O(N__58115),
            .I(N__58109));
    LocalMux I__14547 (
            .O(N__58112),
            .I(\ADC_VDC.genclk.t0on_2 ));
    LocalMux I__14546 (
            .O(N__58109),
            .I(\ADC_VDC.genclk.t0on_2 ));
    CascadeMux I__14545 (
            .O(N__58104),
            .I(N__58100));
    InMux I__14544 (
            .O(N__58103),
            .I(N__58097));
    InMux I__14543 (
            .O(N__58100),
            .I(N__58094));
    LocalMux I__14542 (
            .O(N__58097),
            .I(\ADC_VDC.genclk.t0on_7 ));
    LocalMux I__14541 (
            .O(N__58094),
            .I(\ADC_VDC.genclk.t0on_7 ));
    InMux I__14540 (
            .O(N__58089),
            .I(N__58085));
    InMux I__14539 (
            .O(N__58088),
            .I(N__58082));
    LocalMux I__14538 (
            .O(N__58085),
            .I(\ADC_VDC.genclk.t0on_10 ));
    LocalMux I__14537 (
            .O(N__58082),
            .I(\ADC_VDC.genclk.t0on_10 ));
    InMux I__14536 (
            .O(N__58077),
            .I(N__58074));
    LocalMux I__14535 (
            .O(N__58074),
            .I(\ADC_VDC.genclk.n27_adj_1396 ));
    InMux I__14534 (
            .O(N__58071),
            .I(N__58067));
    InMux I__14533 (
            .O(N__58070),
            .I(N__58064));
    LocalMux I__14532 (
            .O(N__58067),
            .I(\ADC_VDC.genclk.t0on_3 ));
    LocalMux I__14531 (
            .O(N__58064),
            .I(\ADC_VDC.genclk.t0on_3 ));
    CascadeMux I__14530 (
            .O(N__58059),
            .I(N__58056));
    InMux I__14529 (
            .O(N__58056),
            .I(N__58052));
    InMux I__14528 (
            .O(N__58055),
            .I(N__58049));
    LocalMux I__14527 (
            .O(N__58052),
            .I(\ADC_VDC.genclk.t0on_13 ));
    LocalMux I__14526 (
            .O(N__58049),
            .I(\ADC_VDC.genclk.t0on_13 ));
    CascadeMux I__14525 (
            .O(N__58044),
            .I(N__58040));
    InMux I__14524 (
            .O(N__58043),
            .I(N__58037));
    InMux I__14523 (
            .O(N__58040),
            .I(N__58034));
    LocalMux I__14522 (
            .O(N__58037),
            .I(\ADC_VDC.genclk.t0on_5 ));
    LocalMux I__14521 (
            .O(N__58034),
            .I(\ADC_VDC.genclk.t0on_5 ));
    InMux I__14520 (
            .O(N__58029),
            .I(N__58025));
    InMux I__14519 (
            .O(N__58028),
            .I(N__58022));
    LocalMux I__14518 (
            .O(N__58025),
            .I(\ADC_VDC.genclk.t0on_8 ));
    LocalMux I__14517 (
            .O(N__58022),
            .I(\ADC_VDC.genclk.t0on_8 ));
    InMux I__14516 (
            .O(N__58017),
            .I(N__58014));
    LocalMux I__14515 (
            .O(N__58014),
            .I(\ADC_VDC.genclk.n26_adj_1395 ));
    InMux I__14514 (
            .O(N__58011),
            .I(N__58007));
    InMux I__14513 (
            .O(N__58010),
            .I(N__57999));
    LocalMux I__14512 (
            .O(N__58007),
            .I(N__57996));
    InMux I__14511 (
            .O(N__58006),
            .I(N__57993));
    InMux I__14510 (
            .O(N__58005),
            .I(N__57986));
    InMux I__14509 (
            .O(N__58004),
            .I(N__57986));
    InMux I__14508 (
            .O(N__58003),
            .I(N__57986));
    InMux I__14507 (
            .O(N__58002),
            .I(N__57983));
    LocalMux I__14506 (
            .O(N__57999),
            .I(N__57978));
    Span4Mux_h I__14505 (
            .O(N__57996),
            .I(N__57978));
    LocalMux I__14504 (
            .O(N__57993),
            .I(N__57975));
    LocalMux I__14503 (
            .O(N__57986),
            .I(N__57972));
    LocalMux I__14502 (
            .O(N__57983),
            .I(\ADC_VDC.genclk.div_state_1 ));
    Odrv4 I__14501 (
            .O(N__57978),
            .I(\ADC_VDC.genclk.div_state_1 ));
    Odrv4 I__14500 (
            .O(N__57975),
            .I(\ADC_VDC.genclk.div_state_1 ));
    Odrv4 I__14499 (
            .O(N__57972),
            .I(\ADC_VDC.genclk.div_state_1 ));
    CEMux I__14498 (
            .O(N__57963),
            .I(N__57960));
    LocalMux I__14497 (
            .O(N__57960),
            .I(N__57956));
    CEMux I__14496 (
            .O(N__57959),
            .I(N__57953));
    Span4Mux_v I__14495 (
            .O(N__57956),
            .I(N__57950));
    LocalMux I__14494 (
            .O(N__57953),
            .I(N__57947));
    Span4Mux_h I__14493 (
            .O(N__57950),
            .I(N__57944));
    Span4Mux_h I__14492 (
            .O(N__57947),
            .I(N__57941));
    Odrv4 I__14491 (
            .O(N__57944),
            .I(\ADC_VDC.genclk.div_state_1__N_1274 ));
    Odrv4 I__14490 (
            .O(N__57941),
            .I(\ADC_VDC.genclk.div_state_1__N_1274 ));
    InMux I__14489 (
            .O(N__57936),
            .I(N__57932));
    InMux I__14488 (
            .O(N__57935),
            .I(N__57929));
    LocalMux I__14487 (
            .O(N__57932),
            .I(\ADC_VDC.genclk.t0on_14 ));
    LocalMux I__14486 (
            .O(N__57929),
            .I(\ADC_VDC.genclk.t0on_14 ));
    CascadeMux I__14485 (
            .O(N__57924),
            .I(N__57921));
    InMux I__14484 (
            .O(N__57921),
            .I(N__57917));
    InMux I__14483 (
            .O(N__57920),
            .I(N__57914));
    LocalMux I__14482 (
            .O(N__57917),
            .I(\ADC_VDC.genclk.t0on_9 ));
    LocalMux I__14481 (
            .O(N__57914),
            .I(\ADC_VDC.genclk.t0on_9 ));
    CascadeMux I__14480 (
            .O(N__57909),
            .I(N__57905));
    InMux I__14479 (
            .O(N__57908),
            .I(N__57902));
    InMux I__14478 (
            .O(N__57905),
            .I(N__57899));
    LocalMux I__14477 (
            .O(N__57902),
            .I(\ADC_VDC.genclk.t0on_15 ));
    LocalMux I__14476 (
            .O(N__57899),
            .I(\ADC_VDC.genclk.t0on_15 ));
    CascadeMux I__14475 (
            .O(N__57894),
            .I(N__57891));
    InMux I__14474 (
            .O(N__57891),
            .I(N__57887));
    InMux I__14473 (
            .O(N__57890),
            .I(N__57884));
    LocalMux I__14472 (
            .O(N__57887),
            .I(\ADC_VDC.genclk.t0on_11 ));
    LocalMux I__14471 (
            .O(N__57884),
            .I(\ADC_VDC.genclk.t0on_11 ));
    InMux I__14470 (
            .O(N__57879),
            .I(N__57876));
    LocalMux I__14469 (
            .O(N__57876),
            .I(N__57873));
    Odrv4 I__14468 (
            .O(N__57873),
            .I(\ADC_VDC.genclk.n28 ));
    InMux I__14467 (
            .O(N__57870),
            .I(\ADC_VDC.genclk.n19728 ));
    InMux I__14466 (
            .O(N__57867),
            .I(\ADC_VDC.genclk.n19729 ));
    InMux I__14465 (
            .O(N__57864),
            .I(\ADC_VDC.genclk.n19730 ));
    InMux I__14464 (
            .O(N__57861),
            .I(bfn_22_8_0_));
    InMux I__14463 (
            .O(N__57858),
            .I(\ADC_VDC.genclk.n19732 ));
    InMux I__14462 (
            .O(N__57855),
            .I(\ADC_VDC.genclk.n19733 ));
    InMux I__14461 (
            .O(N__57852),
            .I(\ADC_VDC.genclk.n19734 ));
    InMux I__14460 (
            .O(N__57849),
            .I(\ADC_VDC.genclk.n19735 ));
    InMux I__14459 (
            .O(N__57846),
            .I(\ADC_VDC.genclk.n19736 ));
    InMux I__14458 (
            .O(N__57843),
            .I(N__57840));
    LocalMux I__14457 (
            .O(N__57840),
            .I(buf_data_iac_13));
    InMux I__14456 (
            .O(N__57837),
            .I(N__57834));
    LocalMux I__14455 (
            .O(N__57834),
            .I(n21350));
    InMux I__14454 (
            .O(N__57831),
            .I(N__57828));
    LocalMux I__14453 (
            .O(N__57828),
            .I(buf_data_iac_9));
    CascadeMux I__14452 (
            .O(N__57825),
            .I(N__57809));
    InMux I__14451 (
            .O(N__57824),
            .I(N__57797));
    InMux I__14450 (
            .O(N__57823),
            .I(N__57789));
    InMux I__14449 (
            .O(N__57822),
            .I(N__57773));
    InMux I__14448 (
            .O(N__57821),
            .I(N__57770));
    InMux I__14447 (
            .O(N__57820),
            .I(N__57767));
    CascadeMux I__14446 (
            .O(N__57819),
            .I(N__57764));
    InMux I__14445 (
            .O(N__57818),
            .I(N__57760));
    InMux I__14444 (
            .O(N__57817),
            .I(N__57751));
    InMux I__14443 (
            .O(N__57816),
            .I(N__57744));
    InMux I__14442 (
            .O(N__57815),
            .I(N__57741));
    InMux I__14441 (
            .O(N__57814),
            .I(N__57729));
    InMux I__14440 (
            .O(N__57813),
            .I(N__57729));
    InMux I__14439 (
            .O(N__57812),
            .I(N__57729));
    InMux I__14438 (
            .O(N__57809),
            .I(N__57724));
    InMux I__14437 (
            .O(N__57808),
            .I(N__57724));
    InMux I__14436 (
            .O(N__57807),
            .I(N__57717));
    InMux I__14435 (
            .O(N__57806),
            .I(N__57717));
    InMux I__14434 (
            .O(N__57805),
            .I(N__57717));
    InMux I__14433 (
            .O(N__57804),
            .I(N__57714));
    InMux I__14432 (
            .O(N__57803),
            .I(N__57705));
    InMux I__14431 (
            .O(N__57802),
            .I(N__57705));
    InMux I__14430 (
            .O(N__57801),
            .I(N__57705));
    InMux I__14429 (
            .O(N__57800),
            .I(N__57705));
    LocalMux I__14428 (
            .O(N__57797),
            .I(N__57702));
    InMux I__14427 (
            .O(N__57796),
            .I(N__57695));
    InMux I__14426 (
            .O(N__57795),
            .I(N__57690));
    InMux I__14425 (
            .O(N__57794),
            .I(N__57690));
    InMux I__14424 (
            .O(N__57793),
            .I(N__57685));
    InMux I__14423 (
            .O(N__57792),
            .I(N__57685));
    LocalMux I__14422 (
            .O(N__57789),
            .I(N__57682));
    InMux I__14421 (
            .O(N__57788),
            .I(N__57675));
    InMux I__14420 (
            .O(N__57787),
            .I(N__57675));
    InMux I__14419 (
            .O(N__57786),
            .I(N__57675));
    InMux I__14418 (
            .O(N__57785),
            .I(N__57672));
    InMux I__14417 (
            .O(N__57784),
            .I(N__57669));
    InMux I__14416 (
            .O(N__57783),
            .I(N__57662));
    InMux I__14415 (
            .O(N__57782),
            .I(N__57658));
    InMux I__14414 (
            .O(N__57781),
            .I(N__57655));
    InMux I__14413 (
            .O(N__57780),
            .I(N__57648));
    InMux I__14412 (
            .O(N__57779),
            .I(N__57643));
    InMux I__14411 (
            .O(N__57778),
            .I(N__57643));
    InMux I__14410 (
            .O(N__57777),
            .I(N__57638));
    InMux I__14409 (
            .O(N__57776),
            .I(N__57635));
    LocalMux I__14408 (
            .O(N__57773),
            .I(N__57632));
    LocalMux I__14407 (
            .O(N__57770),
            .I(N__57627));
    LocalMux I__14406 (
            .O(N__57767),
            .I(N__57627));
    InMux I__14405 (
            .O(N__57764),
            .I(N__57619));
    InMux I__14404 (
            .O(N__57763),
            .I(N__57619));
    LocalMux I__14403 (
            .O(N__57760),
            .I(N__57611));
    InMux I__14402 (
            .O(N__57759),
            .I(N__57608));
    InMux I__14401 (
            .O(N__57758),
            .I(N__57605));
    InMux I__14400 (
            .O(N__57757),
            .I(N__57600));
    InMux I__14399 (
            .O(N__57756),
            .I(N__57597));
    InMux I__14398 (
            .O(N__57755),
            .I(N__57594));
    InMux I__14397 (
            .O(N__57754),
            .I(N__57585));
    LocalMux I__14396 (
            .O(N__57751),
            .I(N__57582));
    InMux I__14395 (
            .O(N__57750),
            .I(N__57579));
    InMux I__14394 (
            .O(N__57749),
            .I(N__57576));
    InMux I__14393 (
            .O(N__57748),
            .I(N__57573));
    InMux I__14392 (
            .O(N__57747),
            .I(N__57569));
    LocalMux I__14391 (
            .O(N__57744),
            .I(N__57564));
    LocalMux I__14390 (
            .O(N__57741),
            .I(N__57564));
    InMux I__14389 (
            .O(N__57740),
            .I(N__57561));
    InMux I__14388 (
            .O(N__57739),
            .I(N__57558));
    InMux I__14387 (
            .O(N__57738),
            .I(N__57555));
    InMux I__14386 (
            .O(N__57737),
            .I(N__57550));
    InMux I__14385 (
            .O(N__57736),
            .I(N__57547));
    LocalMux I__14384 (
            .O(N__57729),
            .I(N__57544));
    LocalMux I__14383 (
            .O(N__57724),
            .I(N__57539));
    LocalMux I__14382 (
            .O(N__57717),
            .I(N__57539));
    LocalMux I__14381 (
            .O(N__57714),
            .I(N__57532));
    LocalMux I__14380 (
            .O(N__57705),
            .I(N__57532));
    Span4Mux_h I__14379 (
            .O(N__57702),
            .I(N__57532));
    InMux I__14378 (
            .O(N__57701),
            .I(N__57527));
    InMux I__14377 (
            .O(N__57700),
            .I(N__57527));
    InMux I__14376 (
            .O(N__57699),
            .I(N__57524));
    InMux I__14375 (
            .O(N__57698),
            .I(N__57521));
    LocalMux I__14374 (
            .O(N__57695),
            .I(N__57508));
    LocalMux I__14373 (
            .O(N__57690),
            .I(N__57508));
    LocalMux I__14372 (
            .O(N__57685),
            .I(N__57508));
    Span4Mux_h I__14371 (
            .O(N__57682),
            .I(N__57508));
    LocalMux I__14370 (
            .O(N__57675),
            .I(N__57508));
    LocalMux I__14369 (
            .O(N__57672),
            .I(N__57508));
    LocalMux I__14368 (
            .O(N__57669),
            .I(N__57505));
    InMux I__14367 (
            .O(N__57668),
            .I(N__57500));
    InMux I__14366 (
            .O(N__57667),
            .I(N__57500));
    InMux I__14365 (
            .O(N__57666),
            .I(N__57493));
    InMux I__14364 (
            .O(N__57665),
            .I(N__57493));
    LocalMux I__14363 (
            .O(N__57662),
            .I(N__57490));
    InMux I__14362 (
            .O(N__57661),
            .I(N__57487));
    LocalMux I__14361 (
            .O(N__57658),
            .I(N__57484));
    LocalMux I__14360 (
            .O(N__57655),
            .I(N__57481));
    InMux I__14359 (
            .O(N__57654),
            .I(N__57478));
    InMux I__14358 (
            .O(N__57653),
            .I(N__57467));
    InMux I__14357 (
            .O(N__57652),
            .I(N__57467));
    InMux I__14356 (
            .O(N__57651),
            .I(N__57467));
    LocalMux I__14355 (
            .O(N__57648),
            .I(N__57462));
    LocalMux I__14354 (
            .O(N__57643),
            .I(N__57462));
    InMux I__14353 (
            .O(N__57642),
            .I(N__57459));
    InMux I__14352 (
            .O(N__57641),
            .I(N__57456));
    LocalMux I__14351 (
            .O(N__57638),
            .I(N__57451));
    LocalMux I__14350 (
            .O(N__57635),
            .I(N__57451));
    Span4Mux_v I__14349 (
            .O(N__57632),
            .I(N__57446));
    Span4Mux_h I__14348 (
            .O(N__57627),
            .I(N__57446));
    InMux I__14347 (
            .O(N__57626),
            .I(N__57443));
    InMux I__14346 (
            .O(N__57625),
            .I(N__57440));
    InMux I__14345 (
            .O(N__57624),
            .I(N__57437));
    LocalMux I__14344 (
            .O(N__57619),
            .I(N__57434));
    InMux I__14343 (
            .O(N__57618),
            .I(N__57423));
    InMux I__14342 (
            .O(N__57617),
            .I(N__57423));
    InMux I__14341 (
            .O(N__57616),
            .I(N__57423));
    InMux I__14340 (
            .O(N__57615),
            .I(N__57423));
    InMux I__14339 (
            .O(N__57614),
            .I(N__57423));
    Span4Mux_h I__14338 (
            .O(N__57611),
            .I(N__57416));
    LocalMux I__14337 (
            .O(N__57608),
            .I(N__57416));
    LocalMux I__14336 (
            .O(N__57605),
            .I(N__57416));
    InMux I__14335 (
            .O(N__57604),
            .I(N__57411));
    InMux I__14334 (
            .O(N__57603),
            .I(N__57411));
    LocalMux I__14333 (
            .O(N__57600),
            .I(N__57404));
    LocalMux I__14332 (
            .O(N__57597),
            .I(N__57404));
    LocalMux I__14331 (
            .O(N__57594),
            .I(N__57404));
    InMux I__14330 (
            .O(N__57593),
            .I(N__57399));
    InMux I__14329 (
            .O(N__57592),
            .I(N__57399));
    InMux I__14328 (
            .O(N__57591),
            .I(N__57394));
    InMux I__14327 (
            .O(N__57590),
            .I(N__57394));
    InMux I__14326 (
            .O(N__57589),
            .I(N__57389));
    InMux I__14325 (
            .O(N__57588),
            .I(N__57389));
    LocalMux I__14324 (
            .O(N__57585),
            .I(N__57370));
    Sp12to4 I__14323 (
            .O(N__57582),
            .I(N__57370));
    LocalMux I__14322 (
            .O(N__57579),
            .I(N__57370));
    LocalMux I__14321 (
            .O(N__57576),
            .I(N__57370));
    LocalMux I__14320 (
            .O(N__57573),
            .I(N__57370));
    InMux I__14319 (
            .O(N__57572),
            .I(N__57367));
    LocalMux I__14318 (
            .O(N__57569),
            .I(N__57362));
    Sp12to4 I__14317 (
            .O(N__57564),
            .I(N__57362));
    LocalMux I__14316 (
            .O(N__57561),
            .I(N__57355));
    LocalMux I__14315 (
            .O(N__57558),
            .I(N__57355));
    LocalMux I__14314 (
            .O(N__57555),
            .I(N__57355));
    InMux I__14313 (
            .O(N__57554),
            .I(N__57352));
    InMux I__14312 (
            .O(N__57553),
            .I(N__57349));
    LocalMux I__14311 (
            .O(N__57550),
            .I(N__57346));
    LocalMux I__14310 (
            .O(N__57547),
            .I(N__57335));
    Span4Mux_h I__14309 (
            .O(N__57544),
            .I(N__57335));
    Span4Mux_h I__14308 (
            .O(N__57539),
            .I(N__57335));
    Span4Mux_v I__14307 (
            .O(N__57532),
            .I(N__57335));
    LocalMux I__14306 (
            .O(N__57527),
            .I(N__57335));
    LocalMux I__14305 (
            .O(N__57524),
            .I(N__57330));
    LocalMux I__14304 (
            .O(N__57521),
            .I(N__57330));
    Span4Mux_v I__14303 (
            .O(N__57508),
            .I(N__57323));
    Span4Mux_h I__14302 (
            .O(N__57505),
            .I(N__57323));
    LocalMux I__14301 (
            .O(N__57500),
            .I(N__57323));
    InMux I__14300 (
            .O(N__57499),
            .I(N__57320));
    InMux I__14299 (
            .O(N__57498),
            .I(N__57317));
    LocalMux I__14298 (
            .O(N__57493),
            .I(N__57312));
    Span4Mux_v I__14297 (
            .O(N__57490),
            .I(N__57312));
    LocalMux I__14296 (
            .O(N__57487),
            .I(N__57303));
    Span4Mux_h I__14295 (
            .O(N__57484),
            .I(N__57303));
    Span4Mux_h I__14294 (
            .O(N__57481),
            .I(N__57303));
    LocalMux I__14293 (
            .O(N__57478),
            .I(N__57303));
    InMux I__14292 (
            .O(N__57477),
            .I(N__57300));
    InMux I__14291 (
            .O(N__57476),
            .I(N__57293));
    InMux I__14290 (
            .O(N__57475),
            .I(N__57293));
    InMux I__14289 (
            .O(N__57474),
            .I(N__57293));
    LocalMux I__14288 (
            .O(N__57467),
            .I(N__57288));
    Span4Mux_v I__14287 (
            .O(N__57462),
            .I(N__57288));
    LocalMux I__14286 (
            .O(N__57459),
            .I(N__57281));
    LocalMux I__14285 (
            .O(N__57456),
            .I(N__57281));
    Span4Mux_v I__14284 (
            .O(N__57451),
            .I(N__57281));
    Span4Mux_v I__14283 (
            .O(N__57446),
            .I(N__57278));
    LocalMux I__14282 (
            .O(N__57443),
            .I(N__57263));
    LocalMux I__14281 (
            .O(N__57440),
            .I(N__57263));
    LocalMux I__14280 (
            .O(N__57437),
            .I(N__57263));
    Span4Mux_h I__14279 (
            .O(N__57434),
            .I(N__57263));
    LocalMux I__14278 (
            .O(N__57423),
            .I(N__57263));
    Span4Mux_v I__14277 (
            .O(N__57416),
            .I(N__57263));
    LocalMux I__14276 (
            .O(N__57411),
            .I(N__57263));
    Span4Mux_h I__14275 (
            .O(N__57404),
            .I(N__57258));
    LocalMux I__14274 (
            .O(N__57399),
            .I(N__57251));
    LocalMux I__14273 (
            .O(N__57394),
            .I(N__57251));
    LocalMux I__14272 (
            .O(N__57389),
            .I(N__57251));
    InMux I__14271 (
            .O(N__57388),
            .I(N__57246));
    InMux I__14270 (
            .O(N__57387),
            .I(N__57246));
    InMux I__14269 (
            .O(N__57386),
            .I(N__57241));
    InMux I__14268 (
            .O(N__57385),
            .I(N__57241));
    InMux I__14267 (
            .O(N__57384),
            .I(N__57232));
    InMux I__14266 (
            .O(N__57383),
            .I(N__57232));
    InMux I__14265 (
            .O(N__57382),
            .I(N__57232));
    InMux I__14264 (
            .O(N__57381),
            .I(N__57232));
    Span12Mux_v I__14263 (
            .O(N__57370),
            .I(N__57225));
    LocalMux I__14262 (
            .O(N__57367),
            .I(N__57225));
    Span12Mux_v I__14261 (
            .O(N__57362),
            .I(N__57225));
    Span12Mux_h I__14260 (
            .O(N__57355),
            .I(N__57222));
    LocalMux I__14259 (
            .O(N__57352),
            .I(N__57215));
    LocalMux I__14258 (
            .O(N__57349),
            .I(N__57215));
    Span12Mux_h I__14257 (
            .O(N__57346),
            .I(N__57215));
    Span4Mux_h I__14256 (
            .O(N__57335),
            .I(N__57208));
    Span4Mux_h I__14255 (
            .O(N__57330),
            .I(N__57208));
    Span4Mux_h I__14254 (
            .O(N__57323),
            .I(N__57208));
    LocalMux I__14253 (
            .O(N__57320),
            .I(N__57199));
    LocalMux I__14252 (
            .O(N__57317),
            .I(N__57199));
    Span4Mux_h I__14251 (
            .O(N__57312),
            .I(N__57199));
    Span4Mux_v I__14250 (
            .O(N__57303),
            .I(N__57199));
    LocalMux I__14249 (
            .O(N__57300),
            .I(N__57186));
    LocalMux I__14248 (
            .O(N__57293),
            .I(N__57186));
    Span4Mux_h I__14247 (
            .O(N__57288),
            .I(N__57186));
    Span4Mux_h I__14246 (
            .O(N__57281),
            .I(N__57186));
    Span4Mux_v I__14245 (
            .O(N__57278),
            .I(N__57186));
    Span4Mux_v I__14244 (
            .O(N__57263),
            .I(N__57186));
    InMux I__14243 (
            .O(N__57262),
            .I(N__57181));
    InMux I__14242 (
            .O(N__57261),
            .I(N__57181));
    Odrv4 I__14241 (
            .O(N__57258),
            .I(comm_cmd_0));
    Odrv4 I__14240 (
            .O(N__57251),
            .I(comm_cmd_0));
    LocalMux I__14239 (
            .O(N__57246),
            .I(comm_cmd_0));
    LocalMux I__14238 (
            .O(N__57241),
            .I(comm_cmd_0));
    LocalMux I__14237 (
            .O(N__57232),
            .I(comm_cmd_0));
    Odrv12 I__14236 (
            .O(N__57225),
            .I(comm_cmd_0));
    Odrv12 I__14235 (
            .O(N__57222),
            .I(comm_cmd_0));
    Odrv12 I__14234 (
            .O(N__57215),
            .I(comm_cmd_0));
    Odrv4 I__14233 (
            .O(N__57208),
            .I(comm_cmd_0));
    Odrv4 I__14232 (
            .O(N__57199),
            .I(comm_cmd_0));
    Odrv4 I__14231 (
            .O(N__57186),
            .I(comm_cmd_0));
    LocalMux I__14230 (
            .O(N__57181),
            .I(comm_cmd_0));
    InMux I__14229 (
            .O(N__57156),
            .I(N__57153));
    LocalMux I__14228 (
            .O(N__57153),
            .I(N__57150));
    Span12Mux_v I__14227 (
            .O(N__57150),
            .I(N__57147));
    Odrv12 I__14226 (
            .O(N__57147),
            .I(n21529));
    CascadeMux I__14225 (
            .O(N__57144),
            .I(N__57140));
    CascadeMux I__14224 (
            .O(N__57143),
            .I(N__57135));
    InMux I__14223 (
            .O(N__57140),
            .I(N__57127));
    InMux I__14222 (
            .O(N__57139),
            .I(N__57127));
    InMux I__14221 (
            .O(N__57138),
            .I(N__57119));
    InMux I__14220 (
            .O(N__57135),
            .I(N__57115));
    InMux I__14219 (
            .O(N__57134),
            .I(N__57110));
    InMux I__14218 (
            .O(N__57133),
            .I(N__57110));
    CascadeMux I__14217 (
            .O(N__57132),
            .I(N__57105));
    LocalMux I__14216 (
            .O(N__57127),
            .I(N__57102));
    InMux I__14215 (
            .O(N__57126),
            .I(N__57099));
    InMux I__14214 (
            .O(N__57125),
            .I(N__57082));
    InMux I__14213 (
            .O(N__57124),
            .I(N__57082));
    InMux I__14212 (
            .O(N__57123),
            .I(N__57079));
    InMux I__14211 (
            .O(N__57122),
            .I(N__57076));
    LocalMux I__14210 (
            .O(N__57119),
            .I(N__57073));
    SRMux I__14209 (
            .O(N__57118),
            .I(N__57070));
    LocalMux I__14208 (
            .O(N__57115),
            .I(N__57056));
    LocalMux I__14207 (
            .O(N__57110),
            .I(N__57053));
    CascadeMux I__14206 (
            .O(N__57109),
            .I(N__57050));
    CascadeMux I__14205 (
            .O(N__57108),
            .I(N__57046));
    InMux I__14204 (
            .O(N__57105),
            .I(N__57043));
    Span4Mux_v I__14203 (
            .O(N__57102),
            .I(N__57038));
    LocalMux I__14202 (
            .O(N__57099),
            .I(N__57038));
    InMux I__14201 (
            .O(N__57098),
            .I(N__57035));
    InMux I__14200 (
            .O(N__57097),
            .I(N__57032));
    InMux I__14199 (
            .O(N__57096),
            .I(N__57029));
    CascadeMux I__14198 (
            .O(N__57095),
            .I(N__57025));
    InMux I__14197 (
            .O(N__57094),
            .I(N__57016));
    InMux I__14196 (
            .O(N__57093),
            .I(N__57016));
    InMux I__14195 (
            .O(N__57092),
            .I(N__57008));
    InMux I__14194 (
            .O(N__57091),
            .I(N__57008));
    InMux I__14193 (
            .O(N__57090),
            .I(N__57005));
    InMux I__14192 (
            .O(N__57089),
            .I(N__57001));
    CascadeMux I__14191 (
            .O(N__57088),
            .I(N__56996));
    CascadeMux I__14190 (
            .O(N__57087),
            .I(N__56993));
    LocalMux I__14189 (
            .O(N__57082),
            .I(N__56983));
    LocalMux I__14188 (
            .O(N__57079),
            .I(N__56983));
    LocalMux I__14187 (
            .O(N__57076),
            .I(N__56983));
    Span4Mux_h I__14186 (
            .O(N__57073),
            .I(N__56983));
    LocalMux I__14185 (
            .O(N__57070),
            .I(N__56980));
    InMux I__14184 (
            .O(N__57069),
            .I(N__56973));
    InMux I__14183 (
            .O(N__57068),
            .I(N__56973));
    InMux I__14182 (
            .O(N__57067),
            .I(N__56973));
    InMux I__14181 (
            .O(N__57066),
            .I(N__56968));
    InMux I__14180 (
            .O(N__57065),
            .I(N__56968));
    InMux I__14179 (
            .O(N__57064),
            .I(N__56959));
    InMux I__14178 (
            .O(N__57063),
            .I(N__56959));
    InMux I__14177 (
            .O(N__57062),
            .I(N__56959));
    InMux I__14176 (
            .O(N__57061),
            .I(N__56959));
    InMux I__14175 (
            .O(N__57060),
            .I(N__56948));
    InMux I__14174 (
            .O(N__57059),
            .I(N__56948));
    Span4Mux_h I__14173 (
            .O(N__57056),
            .I(N__56940));
    Span4Mux_h I__14172 (
            .O(N__57053),
            .I(N__56940));
    InMux I__14171 (
            .O(N__57050),
            .I(N__56937));
    InMux I__14170 (
            .O(N__57049),
            .I(N__56920));
    InMux I__14169 (
            .O(N__57046),
            .I(N__56917));
    LocalMux I__14168 (
            .O(N__57043),
            .I(N__56914));
    Span4Mux_h I__14167 (
            .O(N__57038),
            .I(N__56905));
    LocalMux I__14166 (
            .O(N__57035),
            .I(N__56905));
    LocalMux I__14165 (
            .O(N__57032),
            .I(N__56905));
    LocalMux I__14164 (
            .O(N__57029),
            .I(N__56905));
    CascadeMux I__14163 (
            .O(N__57028),
            .I(N__56902));
    InMux I__14162 (
            .O(N__57025),
            .I(N__56888));
    InMux I__14161 (
            .O(N__57024),
            .I(N__56888));
    InMux I__14160 (
            .O(N__57023),
            .I(N__56888));
    InMux I__14159 (
            .O(N__57022),
            .I(N__56888));
    InMux I__14158 (
            .O(N__57021),
            .I(N__56888));
    LocalMux I__14157 (
            .O(N__57016),
            .I(N__56885));
    InMux I__14156 (
            .O(N__57015),
            .I(N__56878));
    InMux I__14155 (
            .O(N__57014),
            .I(N__56878));
    InMux I__14154 (
            .O(N__57013),
            .I(N__56878));
    LocalMux I__14153 (
            .O(N__57008),
            .I(N__56875));
    LocalMux I__14152 (
            .O(N__57005),
            .I(N__56872));
    CascadeMux I__14151 (
            .O(N__57004),
            .I(N__56869));
    LocalMux I__14150 (
            .O(N__57001),
            .I(N__56860));
    InMux I__14149 (
            .O(N__57000),
            .I(N__56857));
    InMux I__14148 (
            .O(N__56999),
            .I(N__56854));
    InMux I__14147 (
            .O(N__56996),
            .I(N__56845));
    InMux I__14146 (
            .O(N__56993),
            .I(N__56845));
    InMux I__14145 (
            .O(N__56992),
            .I(N__56845));
    Span4Mux_v I__14144 (
            .O(N__56983),
            .I(N__56842));
    Span4Mux_v I__14143 (
            .O(N__56980),
            .I(N__56835));
    LocalMux I__14142 (
            .O(N__56973),
            .I(N__56835));
    LocalMux I__14141 (
            .O(N__56968),
            .I(N__56835));
    LocalMux I__14140 (
            .O(N__56959),
            .I(N__56832));
    InMux I__14139 (
            .O(N__56958),
            .I(N__56827));
    InMux I__14138 (
            .O(N__56957),
            .I(N__56811));
    InMux I__14137 (
            .O(N__56956),
            .I(N__56811));
    InMux I__14136 (
            .O(N__56955),
            .I(N__56811));
    InMux I__14135 (
            .O(N__56954),
            .I(N__56811));
    InMux I__14134 (
            .O(N__56953),
            .I(N__56811));
    LocalMux I__14133 (
            .O(N__56948),
            .I(N__56808));
    InMux I__14132 (
            .O(N__56947),
            .I(N__56801));
    InMux I__14131 (
            .O(N__56946),
            .I(N__56801));
    InMux I__14130 (
            .O(N__56945),
            .I(N__56801));
    Span4Mux_v I__14129 (
            .O(N__56940),
            .I(N__56796));
    LocalMux I__14128 (
            .O(N__56937),
            .I(N__56796));
    InMux I__14127 (
            .O(N__56936),
            .I(N__56787));
    InMux I__14126 (
            .O(N__56935),
            .I(N__56787));
    InMux I__14125 (
            .O(N__56934),
            .I(N__56787));
    InMux I__14124 (
            .O(N__56933),
            .I(N__56787));
    InMux I__14123 (
            .O(N__56932),
            .I(N__56778));
    InMux I__14122 (
            .O(N__56931),
            .I(N__56778));
    InMux I__14121 (
            .O(N__56930),
            .I(N__56778));
    InMux I__14120 (
            .O(N__56929),
            .I(N__56778));
    InMux I__14119 (
            .O(N__56928),
            .I(N__56773));
    InMux I__14118 (
            .O(N__56927),
            .I(N__56773));
    InMux I__14117 (
            .O(N__56926),
            .I(N__56768));
    InMux I__14116 (
            .O(N__56925),
            .I(N__56768));
    InMux I__14115 (
            .O(N__56924),
            .I(N__56763));
    InMux I__14114 (
            .O(N__56923),
            .I(N__56763));
    LocalMux I__14113 (
            .O(N__56920),
            .I(N__56760));
    LocalMux I__14112 (
            .O(N__56917),
            .I(N__56757));
    Span4Mux_h I__14111 (
            .O(N__56914),
            .I(N__56752));
    Span4Mux_v I__14110 (
            .O(N__56905),
            .I(N__56752));
    InMux I__14109 (
            .O(N__56902),
            .I(N__56743));
    InMux I__14108 (
            .O(N__56901),
            .I(N__56743));
    InMux I__14107 (
            .O(N__56900),
            .I(N__56743));
    InMux I__14106 (
            .O(N__56899),
            .I(N__56743));
    LocalMux I__14105 (
            .O(N__56888),
            .I(N__56732));
    Span4Mux_h I__14104 (
            .O(N__56885),
            .I(N__56732));
    LocalMux I__14103 (
            .O(N__56878),
            .I(N__56732));
    Span4Mux_h I__14102 (
            .O(N__56875),
            .I(N__56732));
    Span4Mux_v I__14101 (
            .O(N__56872),
            .I(N__56732));
    InMux I__14100 (
            .O(N__56869),
            .I(N__56727));
    InMux I__14099 (
            .O(N__56868),
            .I(N__56727));
    InMux I__14098 (
            .O(N__56867),
            .I(N__56724));
    InMux I__14097 (
            .O(N__56866),
            .I(N__56715));
    InMux I__14096 (
            .O(N__56865),
            .I(N__56715));
    InMux I__14095 (
            .O(N__56864),
            .I(N__56715));
    InMux I__14094 (
            .O(N__56863),
            .I(N__56715));
    Sp12to4 I__14093 (
            .O(N__56860),
            .I(N__56708));
    LocalMux I__14092 (
            .O(N__56857),
            .I(N__56708));
    LocalMux I__14091 (
            .O(N__56854),
            .I(N__56708));
    InMux I__14090 (
            .O(N__56853),
            .I(N__56703));
    InMux I__14089 (
            .O(N__56852),
            .I(N__56703));
    LocalMux I__14088 (
            .O(N__56845),
            .I(N__56694));
    Span4Mux_v I__14087 (
            .O(N__56842),
            .I(N__56694));
    Span4Mux_h I__14086 (
            .O(N__56835),
            .I(N__56694));
    Span4Mux_h I__14085 (
            .O(N__56832),
            .I(N__56694));
    InMux I__14084 (
            .O(N__56831),
            .I(N__56689));
    InMux I__14083 (
            .O(N__56830),
            .I(N__56686));
    LocalMux I__14082 (
            .O(N__56827),
            .I(N__56683));
    InMux I__14081 (
            .O(N__56826),
            .I(N__56676));
    InMux I__14080 (
            .O(N__56825),
            .I(N__56676));
    InMux I__14079 (
            .O(N__56824),
            .I(N__56676));
    InMux I__14078 (
            .O(N__56823),
            .I(N__56671));
    InMux I__14077 (
            .O(N__56822),
            .I(N__56671));
    LocalMux I__14076 (
            .O(N__56811),
            .I(N__56668));
    Sp12to4 I__14075 (
            .O(N__56808),
            .I(N__56651));
    LocalMux I__14074 (
            .O(N__56801),
            .I(N__56651));
    Sp12to4 I__14073 (
            .O(N__56796),
            .I(N__56651));
    LocalMux I__14072 (
            .O(N__56787),
            .I(N__56651));
    LocalMux I__14071 (
            .O(N__56778),
            .I(N__56651));
    LocalMux I__14070 (
            .O(N__56773),
            .I(N__56651));
    LocalMux I__14069 (
            .O(N__56768),
            .I(N__56651));
    LocalMux I__14068 (
            .O(N__56763),
            .I(N__56651));
    Span4Mux_h I__14067 (
            .O(N__56760),
            .I(N__56640));
    Span4Mux_v I__14066 (
            .O(N__56757),
            .I(N__56640));
    Span4Mux_h I__14065 (
            .O(N__56752),
            .I(N__56640));
    LocalMux I__14064 (
            .O(N__56743),
            .I(N__56640));
    Span4Mux_v I__14063 (
            .O(N__56732),
            .I(N__56640));
    LocalMux I__14062 (
            .O(N__56727),
            .I(N__56629));
    LocalMux I__14061 (
            .O(N__56724),
            .I(N__56629));
    LocalMux I__14060 (
            .O(N__56715),
            .I(N__56629));
    Span12Mux_v I__14059 (
            .O(N__56708),
            .I(N__56629));
    LocalMux I__14058 (
            .O(N__56703),
            .I(N__56629));
    Span4Mux_h I__14057 (
            .O(N__56694),
            .I(N__56626));
    InMux I__14056 (
            .O(N__56693),
            .I(N__56621));
    InMux I__14055 (
            .O(N__56692),
            .I(N__56621));
    LocalMux I__14054 (
            .O(N__56689),
            .I(comm_state_3));
    LocalMux I__14053 (
            .O(N__56686),
            .I(comm_state_3));
    Odrv4 I__14052 (
            .O(N__56683),
            .I(comm_state_3));
    LocalMux I__14051 (
            .O(N__56676),
            .I(comm_state_3));
    LocalMux I__14050 (
            .O(N__56671),
            .I(comm_state_3));
    Odrv4 I__14049 (
            .O(N__56668),
            .I(comm_state_3));
    Odrv12 I__14048 (
            .O(N__56651),
            .I(comm_state_3));
    Odrv4 I__14047 (
            .O(N__56640),
            .I(comm_state_3));
    Odrv12 I__14046 (
            .O(N__56629),
            .I(comm_state_3));
    Odrv4 I__14045 (
            .O(N__56626),
            .I(comm_state_3));
    LocalMux I__14044 (
            .O(N__56621),
            .I(comm_state_3));
    CascadeMux I__14043 (
            .O(N__56598),
            .I(N__56595));
    InMux I__14042 (
            .O(N__56595),
            .I(N__56591));
    InMux I__14041 (
            .O(N__56594),
            .I(N__56588));
    LocalMux I__14040 (
            .O(N__56591),
            .I(N__56585));
    LocalMux I__14039 (
            .O(N__56588),
            .I(N__56582));
    Span4Mux_v I__14038 (
            .O(N__56585),
            .I(N__56579));
    Span4Mux_v I__14037 (
            .O(N__56582),
            .I(N__56576));
    Span4Mux_h I__14036 (
            .O(N__56579),
            .I(N__56571));
    Span4Mux_h I__14035 (
            .O(N__56576),
            .I(N__56571));
    Odrv4 I__14034 (
            .O(N__56571),
            .I(n17489));
    CascadeMux I__14033 (
            .O(N__56568),
            .I(N__56564));
    CascadeMux I__14032 (
            .O(N__56567),
            .I(N__56541));
    InMux I__14031 (
            .O(N__56564),
            .I(N__56532));
    InMux I__14030 (
            .O(N__56563),
            .I(N__56532));
    InMux I__14029 (
            .O(N__56562),
            .I(N__56532));
    InMux I__14028 (
            .O(N__56561),
            .I(N__56527));
    InMux I__14027 (
            .O(N__56560),
            .I(N__56527));
    InMux I__14026 (
            .O(N__56559),
            .I(N__56520));
    InMux I__14025 (
            .O(N__56558),
            .I(N__56520));
    InMux I__14024 (
            .O(N__56557),
            .I(N__56520));
    CascadeMux I__14023 (
            .O(N__56556),
            .I(N__56513));
    InMux I__14022 (
            .O(N__56555),
            .I(N__56509));
    InMux I__14021 (
            .O(N__56554),
            .I(N__56506));
    CascadeMux I__14020 (
            .O(N__56553),
            .I(N__56501));
    InMux I__14019 (
            .O(N__56552),
            .I(N__56494));
    InMux I__14018 (
            .O(N__56551),
            .I(N__56489));
    InMux I__14017 (
            .O(N__56550),
            .I(N__56489));
    CascadeMux I__14016 (
            .O(N__56549),
            .I(N__56485));
    CascadeMux I__14015 (
            .O(N__56548),
            .I(N__56468));
    InMux I__14014 (
            .O(N__56547),
            .I(N__56459));
    InMux I__14013 (
            .O(N__56546),
            .I(N__56459));
    InMux I__14012 (
            .O(N__56545),
            .I(N__56459));
    InMux I__14011 (
            .O(N__56544),
            .I(N__56456));
    InMux I__14010 (
            .O(N__56541),
            .I(N__56453));
    CascadeMux I__14009 (
            .O(N__56540),
            .I(N__56447));
    CascadeMux I__14008 (
            .O(N__56539),
            .I(N__56442));
    LocalMux I__14007 (
            .O(N__56532),
            .I(N__56433));
    LocalMux I__14006 (
            .O(N__56527),
            .I(N__56433));
    LocalMux I__14005 (
            .O(N__56520),
            .I(N__56433));
    InMux I__14004 (
            .O(N__56519),
            .I(N__56430));
    CascadeMux I__14003 (
            .O(N__56518),
            .I(N__56427));
    CascadeMux I__14002 (
            .O(N__56517),
            .I(N__56424));
    CascadeMux I__14001 (
            .O(N__56516),
            .I(N__56421));
    InMux I__14000 (
            .O(N__56513),
            .I(N__56414));
    InMux I__13999 (
            .O(N__56512),
            .I(N__56414));
    LocalMux I__13998 (
            .O(N__56509),
            .I(N__56409));
    LocalMux I__13997 (
            .O(N__56506),
            .I(N__56409));
    InMux I__13996 (
            .O(N__56505),
            .I(N__56406));
    InMux I__13995 (
            .O(N__56504),
            .I(N__56401));
    InMux I__13994 (
            .O(N__56501),
            .I(N__56401));
    InMux I__13993 (
            .O(N__56500),
            .I(N__56395));
    InMux I__13992 (
            .O(N__56499),
            .I(N__56395));
    InMux I__13991 (
            .O(N__56498),
            .I(N__56390));
    InMux I__13990 (
            .O(N__56497),
            .I(N__56390));
    LocalMux I__13989 (
            .O(N__56494),
            .I(N__56387));
    LocalMux I__13988 (
            .O(N__56489),
            .I(N__56384));
    InMux I__13987 (
            .O(N__56488),
            .I(N__56379));
    InMux I__13986 (
            .O(N__56485),
            .I(N__56379));
    InMux I__13985 (
            .O(N__56484),
            .I(N__56364));
    InMux I__13984 (
            .O(N__56483),
            .I(N__56364));
    InMux I__13983 (
            .O(N__56482),
            .I(N__56364));
    InMux I__13982 (
            .O(N__56481),
            .I(N__56364));
    InMux I__13981 (
            .O(N__56480),
            .I(N__56364));
    InMux I__13980 (
            .O(N__56479),
            .I(N__56364));
    InMux I__13979 (
            .O(N__56478),
            .I(N__56364));
    CascadeMux I__13978 (
            .O(N__56477),
            .I(N__56361));
    CascadeMux I__13977 (
            .O(N__56476),
            .I(N__56358));
    InMux I__13976 (
            .O(N__56475),
            .I(N__56351));
    InMux I__13975 (
            .O(N__56474),
            .I(N__56351));
    CascadeMux I__13974 (
            .O(N__56473),
            .I(N__56348));
    CascadeMux I__13973 (
            .O(N__56472),
            .I(N__56345));
    InMux I__13972 (
            .O(N__56471),
            .I(N__56334));
    InMux I__13971 (
            .O(N__56468),
            .I(N__56334));
    InMux I__13970 (
            .O(N__56467),
            .I(N__56334));
    InMux I__13969 (
            .O(N__56466),
            .I(N__56334));
    LocalMux I__13968 (
            .O(N__56459),
            .I(N__56331));
    LocalMux I__13967 (
            .O(N__56456),
            .I(N__56328));
    LocalMux I__13966 (
            .O(N__56453),
            .I(N__56325));
    InMux I__13965 (
            .O(N__56452),
            .I(N__56322));
    InMux I__13964 (
            .O(N__56451),
            .I(N__56317));
    InMux I__13963 (
            .O(N__56450),
            .I(N__56312));
    InMux I__13962 (
            .O(N__56447),
            .I(N__56305));
    InMux I__13961 (
            .O(N__56446),
            .I(N__56305));
    InMux I__13960 (
            .O(N__56445),
            .I(N__56305));
    InMux I__13959 (
            .O(N__56442),
            .I(N__56298));
    InMux I__13958 (
            .O(N__56441),
            .I(N__56298));
    InMux I__13957 (
            .O(N__56440),
            .I(N__56298));
    Span4Mux_v I__13956 (
            .O(N__56433),
            .I(N__56293));
    LocalMux I__13955 (
            .O(N__56430),
            .I(N__56293));
    InMux I__13954 (
            .O(N__56427),
            .I(N__56288));
    InMux I__13953 (
            .O(N__56424),
            .I(N__56281));
    InMux I__13952 (
            .O(N__56421),
            .I(N__56281));
    InMux I__13951 (
            .O(N__56420),
            .I(N__56281));
    InMux I__13950 (
            .O(N__56419),
            .I(N__56278));
    LocalMux I__13949 (
            .O(N__56414),
            .I(N__56275));
    Span4Mux_v I__13948 (
            .O(N__56409),
            .I(N__56272));
    LocalMux I__13947 (
            .O(N__56406),
            .I(N__56267));
    LocalMux I__13946 (
            .O(N__56401),
            .I(N__56267));
    InMux I__13945 (
            .O(N__56400),
            .I(N__56264));
    LocalMux I__13944 (
            .O(N__56395),
            .I(N__56253));
    LocalMux I__13943 (
            .O(N__56390),
            .I(N__56253));
    Span4Mux_h I__13942 (
            .O(N__56387),
            .I(N__56253));
    Span4Mux_h I__13941 (
            .O(N__56384),
            .I(N__56253));
    LocalMux I__13940 (
            .O(N__56379),
            .I(N__56253));
    LocalMux I__13939 (
            .O(N__56364),
            .I(N__56250));
    InMux I__13938 (
            .O(N__56361),
            .I(N__56247));
    InMux I__13937 (
            .O(N__56358),
            .I(N__56240));
    InMux I__13936 (
            .O(N__56357),
            .I(N__56240));
    InMux I__13935 (
            .O(N__56356),
            .I(N__56240));
    LocalMux I__13934 (
            .O(N__56351),
            .I(N__56237));
    InMux I__13933 (
            .O(N__56348),
            .I(N__56232));
    InMux I__13932 (
            .O(N__56345),
            .I(N__56232));
    CascadeMux I__13931 (
            .O(N__56344),
            .I(N__56229));
    CascadeMux I__13930 (
            .O(N__56343),
            .I(N__56224));
    LocalMux I__13929 (
            .O(N__56334),
            .I(N__56215));
    Span4Mux_v I__13928 (
            .O(N__56331),
            .I(N__56215));
    Span4Mux_h I__13927 (
            .O(N__56328),
            .I(N__56212));
    Span4Mux_h I__13926 (
            .O(N__56325),
            .I(N__56207));
    LocalMux I__13925 (
            .O(N__56322),
            .I(N__56207));
    CascadeMux I__13924 (
            .O(N__56321),
            .I(N__56204));
    CascadeMux I__13923 (
            .O(N__56320),
            .I(N__56199));
    LocalMux I__13922 (
            .O(N__56317),
            .I(N__56196));
    InMux I__13921 (
            .O(N__56316),
            .I(N__56191));
    InMux I__13920 (
            .O(N__56315),
            .I(N__56191));
    LocalMux I__13919 (
            .O(N__56312),
            .I(N__56188));
    LocalMux I__13918 (
            .O(N__56305),
            .I(N__56181));
    LocalMux I__13917 (
            .O(N__56298),
            .I(N__56181));
    Span4Mux_h I__13916 (
            .O(N__56293),
            .I(N__56181));
    CascadeMux I__13915 (
            .O(N__56292),
            .I(N__56176));
    CascadeMux I__13914 (
            .O(N__56291),
            .I(N__56171));
    LocalMux I__13913 (
            .O(N__56288),
            .I(N__56165));
    LocalMux I__13912 (
            .O(N__56281),
            .I(N__56160));
    LocalMux I__13911 (
            .O(N__56278),
            .I(N__56160));
    Span4Mux_v I__13910 (
            .O(N__56275),
            .I(N__56157));
    Span4Mux_h I__13909 (
            .O(N__56272),
            .I(N__56146));
    Span4Mux_v I__13908 (
            .O(N__56267),
            .I(N__56146));
    LocalMux I__13907 (
            .O(N__56264),
            .I(N__56146));
    Span4Mux_v I__13906 (
            .O(N__56253),
            .I(N__56146));
    Span4Mux_v I__13905 (
            .O(N__56250),
            .I(N__56146));
    LocalMux I__13904 (
            .O(N__56247),
            .I(N__56143));
    LocalMux I__13903 (
            .O(N__56240),
            .I(N__56136));
    Span4Mux_v I__13902 (
            .O(N__56237),
            .I(N__56136));
    LocalMux I__13901 (
            .O(N__56232),
            .I(N__56136));
    InMux I__13900 (
            .O(N__56229),
            .I(N__56129));
    InMux I__13899 (
            .O(N__56228),
            .I(N__56129));
    InMux I__13898 (
            .O(N__56227),
            .I(N__56129));
    InMux I__13897 (
            .O(N__56224),
            .I(N__56124));
    InMux I__13896 (
            .O(N__56223),
            .I(N__56124));
    InMux I__13895 (
            .O(N__56222),
            .I(N__56121));
    InMux I__13894 (
            .O(N__56221),
            .I(N__56116));
    InMux I__13893 (
            .O(N__56220),
            .I(N__56116));
    Span4Mux_h I__13892 (
            .O(N__56215),
            .I(N__56109));
    Span4Mux_v I__13891 (
            .O(N__56212),
            .I(N__56109));
    Span4Mux_v I__13890 (
            .O(N__56207),
            .I(N__56109));
    InMux I__13889 (
            .O(N__56204),
            .I(N__56100));
    InMux I__13888 (
            .O(N__56203),
            .I(N__56100));
    InMux I__13887 (
            .O(N__56202),
            .I(N__56100));
    InMux I__13886 (
            .O(N__56199),
            .I(N__56100));
    Span4Mux_h I__13885 (
            .O(N__56196),
            .I(N__56091));
    LocalMux I__13884 (
            .O(N__56191),
            .I(N__56091));
    Span4Mux_v I__13883 (
            .O(N__56188),
            .I(N__56091));
    Span4Mux_h I__13882 (
            .O(N__56181),
            .I(N__56091));
    InMux I__13881 (
            .O(N__56180),
            .I(N__56084));
    InMux I__13880 (
            .O(N__56179),
            .I(N__56084));
    InMux I__13879 (
            .O(N__56176),
            .I(N__56084));
    InMux I__13878 (
            .O(N__56175),
            .I(N__56075));
    InMux I__13877 (
            .O(N__56174),
            .I(N__56075));
    InMux I__13876 (
            .O(N__56171),
            .I(N__56075));
    InMux I__13875 (
            .O(N__56170),
            .I(N__56075));
    InMux I__13874 (
            .O(N__56169),
            .I(N__56070));
    InMux I__13873 (
            .O(N__56168),
            .I(N__56070));
    Span4Mux_h I__13872 (
            .O(N__56165),
            .I(N__56065));
    Span4Mux_h I__13871 (
            .O(N__56160),
            .I(N__56065));
    Span4Mux_v I__13870 (
            .O(N__56157),
            .I(N__56054));
    Span4Mux_h I__13869 (
            .O(N__56146),
            .I(N__56054));
    Span4Mux_v I__13868 (
            .O(N__56143),
            .I(N__56054));
    Span4Mux_v I__13867 (
            .O(N__56136),
            .I(N__56054));
    LocalMux I__13866 (
            .O(N__56129),
            .I(N__56054));
    LocalMux I__13865 (
            .O(N__56124),
            .I(n9306));
    LocalMux I__13864 (
            .O(N__56121),
            .I(n9306));
    LocalMux I__13863 (
            .O(N__56116),
            .I(n9306));
    Odrv4 I__13862 (
            .O(N__56109),
            .I(n9306));
    LocalMux I__13861 (
            .O(N__56100),
            .I(n9306));
    Odrv4 I__13860 (
            .O(N__56091),
            .I(n9306));
    LocalMux I__13859 (
            .O(N__56084),
            .I(n9306));
    LocalMux I__13858 (
            .O(N__56075),
            .I(n9306));
    LocalMux I__13857 (
            .O(N__56070),
            .I(n9306));
    Odrv4 I__13856 (
            .O(N__56065),
            .I(n9306));
    Odrv4 I__13855 (
            .O(N__56054),
            .I(n9306));
    InMux I__13854 (
            .O(N__56031),
            .I(N__56027));
    InMux I__13853 (
            .O(N__56030),
            .I(N__56024));
    LocalMux I__13852 (
            .O(N__56027),
            .I(N__56021));
    LocalMux I__13851 (
            .O(N__56024),
            .I(N__56018));
    Span4Mux_v I__13850 (
            .O(N__56021),
            .I(N__56015));
    Span4Mux_v I__13849 (
            .O(N__56018),
            .I(N__56010));
    Span4Mux_h I__13848 (
            .O(N__56015),
            .I(N__56010));
    Odrv4 I__13847 (
            .O(N__56010),
            .I(n17487));
    CascadeMux I__13846 (
            .O(N__56007),
            .I(N__56004));
    CascadeBuf I__13845 (
            .O(N__56004),
            .I(N__56001));
    CascadeMux I__13844 (
            .O(N__56001),
            .I(N__55998));
    CascadeBuf I__13843 (
            .O(N__55998),
            .I(N__55995));
    CascadeMux I__13842 (
            .O(N__55995),
            .I(N__55992));
    CascadeBuf I__13841 (
            .O(N__55992),
            .I(N__55989));
    CascadeMux I__13840 (
            .O(N__55989),
            .I(N__55986));
    CascadeBuf I__13839 (
            .O(N__55986),
            .I(N__55983));
    CascadeMux I__13838 (
            .O(N__55983),
            .I(N__55980));
    CascadeBuf I__13837 (
            .O(N__55980),
            .I(N__55977));
    CascadeMux I__13836 (
            .O(N__55977),
            .I(N__55974));
    CascadeBuf I__13835 (
            .O(N__55974),
            .I(N__55971));
    CascadeMux I__13834 (
            .O(N__55971),
            .I(N__55968));
    CascadeBuf I__13833 (
            .O(N__55968),
            .I(N__55964));
    CascadeMux I__13832 (
            .O(N__55967),
            .I(N__55961));
    CascadeMux I__13831 (
            .O(N__55964),
            .I(N__55958));
    CascadeBuf I__13830 (
            .O(N__55961),
            .I(N__55955));
    CascadeBuf I__13829 (
            .O(N__55958),
            .I(N__55952));
    CascadeMux I__13828 (
            .O(N__55955),
            .I(N__55949));
    CascadeMux I__13827 (
            .O(N__55952),
            .I(N__55946));
    InMux I__13826 (
            .O(N__55949),
            .I(N__55943));
    CascadeBuf I__13825 (
            .O(N__55946),
            .I(N__55940));
    LocalMux I__13824 (
            .O(N__55943),
            .I(N__55937));
    CascadeMux I__13823 (
            .O(N__55940),
            .I(N__55934));
    Span12Mux_h I__13822 (
            .O(N__55937),
            .I(N__55931));
    InMux I__13821 (
            .O(N__55934),
            .I(N__55928));
    Span12Mux_v I__13820 (
            .O(N__55931),
            .I(N__55925));
    LocalMux I__13819 (
            .O(N__55928),
            .I(N__55922));
    Odrv12 I__13818 (
            .O(N__55925),
            .I(data_index_9_N_216_5));
    Odrv4 I__13817 (
            .O(N__55922),
            .I(data_index_9_N_216_5));
    InMux I__13816 (
            .O(N__55917),
            .I(bfn_22_7_0_));
    InMux I__13815 (
            .O(N__55914),
            .I(\ADC_VDC.genclk.n19724 ));
    InMux I__13814 (
            .O(N__55911),
            .I(\ADC_VDC.genclk.n19725 ));
    InMux I__13813 (
            .O(N__55908),
            .I(\ADC_VDC.genclk.n19726 ));
    InMux I__13812 (
            .O(N__55905),
            .I(\ADC_VDC.genclk.n19727 ));
    InMux I__13811 (
            .O(N__55902),
            .I(N__55897));
    InMux I__13810 (
            .O(N__55901),
            .I(N__55894));
    InMux I__13809 (
            .O(N__55900),
            .I(N__55891));
    LocalMux I__13808 (
            .O(N__55897),
            .I(N__55888));
    LocalMux I__13807 (
            .O(N__55894),
            .I(N__55885));
    LocalMux I__13806 (
            .O(N__55891),
            .I(N__55882));
    Odrv4 I__13805 (
            .O(N__55888),
            .I(\comm_spi.n14600 ));
    Odrv4 I__13804 (
            .O(N__55885),
            .I(\comm_spi.n14600 ));
    Odrv4 I__13803 (
            .O(N__55882),
            .I(\comm_spi.n14600 ));
    InMux I__13802 (
            .O(N__55875),
            .I(N__55862));
    InMux I__13801 (
            .O(N__55874),
            .I(N__55859));
    CascadeMux I__13800 (
            .O(N__55873),
            .I(N__55854));
    CascadeMux I__13799 (
            .O(N__55872),
            .I(N__55851));
    CascadeMux I__13798 (
            .O(N__55871),
            .I(N__55844));
    SRMux I__13797 (
            .O(N__55870),
            .I(N__55840));
    SRMux I__13796 (
            .O(N__55869),
            .I(N__55837));
    InMux I__13795 (
            .O(N__55868),
            .I(N__55834));
    InMux I__13794 (
            .O(N__55867),
            .I(N__55828));
    InMux I__13793 (
            .O(N__55866),
            .I(N__55824));
    InMux I__13792 (
            .O(N__55865),
            .I(N__55821));
    LocalMux I__13791 (
            .O(N__55862),
            .I(N__55811));
    LocalMux I__13790 (
            .O(N__55859),
            .I(N__55811));
    InMux I__13789 (
            .O(N__55858),
            .I(N__55795));
    InMux I__13788 (
            .O(N__55857),
            .I(N__55795));
    InMux I__13787 (
            .O(N__55854),
            .I(N__55795));
    InMux I__13786 (
            .O(N__55851),
            .I(N__55795));
    InMux I__13785 (
            .O(N__55850),
            .I(N__55795));
    InMux I__13784 (
            .O(N__55849),
            .I(N__55795));
    InMux I__13783 (
            .O(N__55848),
            .I(N__55795));
    InMux I__13782 (
            .O(N__55847),
            .I(N__55792));
    InMux I__13781 (
            .O(N__55844),
            .I(N__55787));
    InMux I__13780 (
            .O(N__55843),
            .I(N__55787));
    LocalMux I__13779 (
            .O(N__55840),
            .I(N__55782));
    LocalMux I__13778 (
            .O(N__55837),
            .I(N__55782));
    LocalMux I__13777 (
            .O(N__55834),
            .I(N__55779));
    InMux I__13776 (
            .O(N__55833),
            .I(N__55772));
    InMux I__13775 (
            .O(N__55832),
            .I(N__55772));
    InMux I__13774 (
            .O(N__55831),
            .I(N__55769));
    LocalMux I__13773 (
            .O(N__55828),
            .I(N__55766));
    InMux I__13772 (
            .O(N__55827),
            .I(N__55760));
    LocalMux I__13771 (
            .O(N__55824),
            .I(N__55752));
    LocalMux I__13770 (
            .O(N__55821),
            .I(N__55752));
    SRMux I__13769 (
            .O(N__55820),
            .I(N__55749));
    InMux I__13768 (
            .O(N__55819),
            .I(N__55742));
    InMux I__13767 (
            .O(N__55818),
            .I(N__55742));
    InMux I__13766 (
            .O(N__55817),
            .I(N__55742));
    InMux I__13765 (
            .O(N__55816),
            .I(N__55739));
    Span4Mux_h I__13764 (
            .O(N__55811),
            .I(N__55736));
    InMux I__13763 (
            .O(N__55810),
            .I(N__55733));
    LocalMux I__13762 (
            .O(N__55795),
            .I(N__55730));
    LocalMux I__13761 (
            .O(N__55792),
            .I(N__55725));
    LocalMux I__13760 (
            .O(N__55787),
            .I(N__55725));
    Span4Mux_h I__13759 (
            .O(N__55782),
            .I(N__55720));
    Span4Mux_h I__13758 (
            .O(N__55779),
            .I(N__55720));
    InMux I__13757 (
            .O(N__55778),
            .I(N__55717));
    InMux I__13756 (
            .O(N__55777),
            .I(N__55714));
    LocalMux I__13755 (
            .O(N__55772),
            .I(N__55709));
    LocalMux I__13754 (
            .O(N__55769),
            .I(N__55709));
    Span4Mux_v I__13753 (
            .O(N__55766),
            .I(N__55706));
    InMux I__13752 (
            .O(N__55765),
            .I(N__55699));
    InMux I__13751 (
            .O(N__55764),
            .I(N__55699));
    InMux I__13750 (
            .O(N__55763),
            .I(N__55699));
    LocalMux I__13749 (
            .O(N__55760),
            .I(N__55696));
    InMux I__13748 (
            .O(N__55759),
            .I(N__55689));
    InMux I__13747 (
            .O(N__55758),
            .I(N__55689));
    InMux I__13746 (
            .O(N__55757),
            .I(N__55689));
    Span4Mux_h I__13745 (
            .O(N__55752),
            .I(N__55680));
    LocalMux I__13744 (
            .O(N__55749),
            .I(N__55680));
    LocalMux I__13743 (
            .O(N__55742),
            .I(N__55680));
    LocalMux I__13742 (
            .O(N__55739),
            .I(N__55680));
    Span4Mux_v I__13741 (
            .O(N__55736),
            .I(N__55677));
    LocalMux I__13740 (
            .O(N__55733),
            .I(N__55674));
    Span4Mux_h I__13739 (
            .O(N__55730),
            .I(N__55667));
    Span4Mux_h I__13738 (
            .O(N__55725),
            .I(N__55667));
    Span4Mux_h I__13737 (
            .O(N__55720),
            .I(N__55667));
    LocalMux I__13736 (
            .O(N__55717),
            .I(N__55656));
    LocalMux I__13735 (
            .O(N__55714),
            .I(N__55656));
    Span12Mux_v I__13734 (
            .O(N__55709),
            .I(N__55656));
    Sp12to4 I__13733 (
            .O(N__55706),
            .I(N__55656));
    LocalMux I__13732 (
            .O(N__55699),
            .I(N__55656));
    Span4Mux_v I__13731 (
            .O(N__55696),
            .I(N__55649));
    LocalMux I__13730 (
            .O(N__55689),
            .I(N__55649));
    Span4Mux_v I__13729 (
            .O(N__55680),
            .I(N__55649));
    Odrv4 I__13728 (
            .O(N__55677),
            .I(comm_clear));
    Odrv4 I__13727 (
            .O(N__55674),
            .I(comm_clear));
    Odrv4 I__13726 (
            .O(N__55667),
            .I(comm_clear));
    Odrv12 I__13725 (
            .O(N__55656),
            .I(comm_clear));
    Odrv4 I__13724 (
            .O(N__55649),
            .I(comm_clear));
    InMux I__13723 (
            .O(N__55638),
            .I(N__55633));
    InMux I__13722 (
            .O(N__55637),
            .I(N__55630));
    InMux I__13721 (
            .O(N__55636),
            .I(N__55627));
    LocalMux I__13720 (
            .O(N__55633),
            .I(N__55624));
    LocalMux I__13719 (
            .O(N__55630),
            .I(N__55621));
    LocalMux I__13718 (
            .O(N__55627),
            .I(N__55618));
    Span4Mux_v I__13717 (
            .O(N__55624),
            .I(N__55615));
    Span4Mux_h I__13716 (
            .O(N__55621),
            .I(N__55611));
    Span4Mux_h I__13715 (
            .O(N__55618),
            .I(N__55608));
    Span4Mux_h I__13714 (
            .O(N__55615),
            .I(N__55605));
    InMux I__13713 (
            .O(N__55614),
            .I(N__55602));
    Span4Mux_h I__13712 (
            .O(N__55611),
            .I(N__55598));
    Span4Mux_v I__13711 (
            .O(N__55608),
            .I(N__55595));
    Sp12to4 I__13710 (
            .O(N__55605),
            .I(N__55590));
    LocalMux I__13709 (
            .O(N__55602),
            .I(N__55590));
    InMux I__13708 (
            .O(N__55601),
            .I(N__55587));
    Sp12to4 I__13707 (
            .O(N__55598),
            .I(N__55578));
    Sp12to4 I__13706 (
            .O(N__55595),
            .I(N__55578));
    Span12Mux_s10_h I__13705 (
            .O(N__55590),
            .I(N__55578));
    LocalMux I__13704 (
            .O(N__55587),
            .I(N__55578));
    Span12Mux_v I__13703 (
            .O(N__55578),
            .I(N__55575));
    Odrv12 I__13702 (
            .O(N__55575),
            .I(ICE_SPI_MOSI));
    SRMux I__13701 (
            .O(N__55572),
            .I(N__55569));
    LocalMux I__13700 (
            .O(N__55569),
            .I(N__55566));
    Span4Mux_h I__13699 (
            .O(N__55566),
            .I(N__55563));
    Odrv4 I__13698 (
            .O(N__55563),
            .I(\comm_spi.imosi_N_752 ));
    InMux I__13697 (
            .O(N__55560),
            .I(N__55557));
    LocalMux I__13696 (
            .O(N__55557),
            .I(N__55553));
    CascadeMux I__13695 (
            .O(N__55556),
            .I(N__55538));
    Span4Mux_h I__13694 (
            .O(N__55553),
            .I(N__55535));
    InMux I__13693 (
            .O(N__55552),
            .I(N__55526));
    InMux I__13692 (
            .O(N__55551),
            .I(N__55526));
    InMux I__13691 (
            .O(N__55550),
            .I(N__55526));
    InMux I__13690 (
            .O(N__55549),
            .I(N__55526));
    InMux I__13689 (
            .O(N__55548),
            .I(N__55519));
    InMux I__13688 (
            .O(N__55547),
            .I(N__55507));
    InMux I__13687 (
            .O(N__55546),
            .I(N__55504));
    InMux I__13686 (
            .O(N__55545),
            .I(N__55501));
    InMux I__13685 (
            .O(N__55544),
            .I(N__55492));
    InMux I__13684 (
            .O(N__55543),
            .I(N__55492));
    InMux I__13683 (
            .O(N__55542),
            .I(N__55492));
    InMux I__13682 (
            .O(N__55541),
            .I(N__55489));
    InMux I__13681 (
            .O(N__55538),
            .I(N__55486));
    Span4Mux_h I__13680 (
            .O(N__55535),
            .I(N__55481));
    LocalMux I__13679 (
            .O(N__55526),
            .I(N__55481));
    InMux I__13678 (
            .O(N__55525),
            .I(N__55473));
    InMux I__13677 (
            .O(N__55524),
            .I(N__55473));
    InMux I__13676 (
            .O(N__55523),
            .I(N__55473));
    InMux I__13675 (
            .O(N__55522),
            .I(N__55470));
    LocalMux I__13674 (
            .O(N__55519),
            .I(N__55467));
    InMux I__13673 (
            .O(N__55518),
            .I(N__55464));
    InMux I__13672 (
            .O(N__55517),
            .I(N__55459));
    InMux I__13671 (
            .O(N__55516),
            .I(N__55459));
    InMux I__13670 (
            .O(N__55515),
            .I(N__55452));
    InMux I__13669 (
            .O(N__55514),
            .I(N__55452));
    InMux I__13668 (
            .O(N__55513),
            .I(N__55452));
    CascadeMux I__13667 (
            .O(N__55512),
            .I(N__55448));
    CascadeMux I__13666 (
            .O(N__55511),
            .I(N__55444));
    CascadeMux I__13665 (
            .O(N__55510),
            .I(N__55441));
    LocalMux I__13664 (
            .O(N__55507),
            .I(N__55434));
    LocalMux I__13663 (
            .O(N__55504),
            .I(N__55434));
    LocalMux I__13662 (
            .O(N__55501),
            .I(N__55434));
    InMux I__13661 (
            .O(N__55500),
            .I(N__55431));
    InMux I__13660 (
            .O(N__55499),
            .I(N__55426));
    LocalMux I__13659 (
            .O(N__55492),
            .I(N__55423));
    LocalMux I__13658 (
            .O(N__55489),
            .I(N__55418));
    LocalMux I__13657 (
            .O(N__55486),
            .I(N__55415));
    Span4Mux_v I__13656 (
            .O(N__55481),
            .I(N__55412));
    InMux I__13655 (
            .O(N__55480),
            .I(N__55409));
    LocalMux I__13654 (
            .O(N__55473),
            .I(N__55397));
    LocalMux I__13653 (
            .O(N__55470),
            .I(N__55397));
    Span4Mux_v I__13652 (
            .O(N__55467),
            .I(N__55397));
    LocalMux I__13651 (
            .O(N__55464),
            .I(N__55394));
    LocalMux I__13650 (
            .O(N__55459),
            .I(N__55391));
    LocalMux I__13649 (
            .O(N__55452),
            .I(N__55388));
    InMux I__13648 (
            .O(N__55451),
            .I(N__55385));
    InMux I__13647 (
            .O(N__55448),
            .I(N__55380));
    InMux I__13646 (
            .O(N__55447),
            .I(N__55380));
    InMux I__13645 (
            .O(N__55444),
            .I(N__55375));
    InMux I__13644 (
            .O(N__55441),
            .I(N__55375));
    Span4Mux_v I__13643 (
            .O(N__55434),
            .I(N__55370));
    LocalMux I__13642 (
            .O(N__55431),
            .I(N__55370));
    InMux I__13641 (
            .O(N__55430),
            .I(N__55365));
    InMux I__13640 (
            .O(N__55429),
            .I(N__55365));
    LocalMux I__13639 (
            .O(N__55426),
            .I(N__55360));
    Span4Mux_h I__13638 (
            .O(N__55423),
            .I(N__55360));
    InMux I__13637 (
            .O(N__55422),
            .I(N__55357));
    InMux I__13636 (
            .O(N__55421),
            .I(N__55354));
    Span4Mux_v I__13635 (
            .O(N__55418),
            .I(N__55339));
    Span4Mux_h I__13634 (
            .O(N__55415),
            .I(N__55339));
    Span4Mux_h I__13633 (
            .O(N__55412),
            .I(N__55339));
    LocalMux I__13632 (
            .O(N__55409),
            .I(N__55339));
    InMux I__13631 (
            .O(N__55408),
            .I(N__55336));
    InMux I__13630 (
            .O(N__55407),
            .I(N__55331));
    InMux I__13629 (
            .O(N__55406),
            .I(N__55331));
    InMux I__13628 (
            .O(N__55405),
            .I(N__55326));
    InMux I__13627 (
            .O(N__55404),
            .I(N__55326));
    Span4Mux_v I__13626 (
            .O(N__55397),
            .I(N__55317));
    Span4Mux_v I__13625 (
            .O(N__55394),
            .I(N__55317));
    Span4Mux_h I__13624 (
            .O(N__55391),
            .I(N__55317));
    Span4Mux_v I__13623 (
            .O(N__55388),
            .I(N__55317));
    LocalMux I__13622 (
            .O(N__55385),
            .I(N__55314));
    LocalMux I__13621 (
            .O(N__55380),
            .I(N__55309));
    LocalMux I__13620 (
            .O(N__55375),
            .I(N__55309));
    Span4Mux_h I__13619 (
            .O(N__55370),
            .I(N__55302));
    LocalMux I__13618 (
            .O(N__55365),
            .I(N__55302));
    Span4Mux_v I__13617 (
            .O(N__55360),
            .I(N__55302));
    LocalMux I__13616 (
            .O(N__55357),
            .I(N__55299));
    LocalMux I__13615 (
            .O(N__55354),
            .I(N__55296));
    InMux I__13614 (
            .O(N__55353),
            .I(N__55287));
    InMux I__13613 (
            .O(N__55352),
            .I(N__55287));
    InMux I__13612 (
            .O(N__55351),
            .I(N__55287));
    InMux I__13611 (
            .O(N__55350),
            .I(N__55287));
    InMux I__13610 (
            .O(N__55349),
            .I(N__55282));
    InMux I__13609 (
            .O(N__55348),
            .I(N__55282));
    Span4Mux_v I__13608 (
            .O(N__55339),
            .I(N__55277));
    LocalMux I__13607 (
            .O(N__55336),
            .I(N__55277));
    LocalMux I__13606 (
            .O(N__55331),
            .I(N__55270));
    LocalMux I__13605 (
            .O(N__55326),
            .I(N__55270));
    Sp12to4 I__13604 (
            .O(N__55317),
            .I(N__55270));
    Span4Mux_h I__13603 (
            .O(N__55314),
            .I(N__55263));
    Span4Mux_v I__13602 (
            .O(N__55309),
            .I(N__55263));
    Span4Mux_v I__13601 (
            .O(N__55302),
            .I(N__55263));
    Odrv4 I__13600 (
            .O(N__55299),
            .I(comm_state_2));
    Odrv12 I__13599 (
            .O(N__55296),
            .I(comm_state_2));
    LocalMux I__13598 (
            .O(N__55287),
            .I(comm_state_2));
    LocalMux I__13597 (
            .O(N__55282),
            .I(comm_state_2));
    Odrv4 I__13596 (
            .O(N__55277),
            .I(comm_state_2));
    Odrv12 I__13595 (
            .O(N__55270),
            .I(comm_state_2));
    Odrv4 I__13594 (
            .O(N__55263),
            .I(comm_state_2));
    CascadeMux I__13593 (
            .O(N__55248),
            .I(N__55245));
    InMux I__13592 (
            .O(N__55245),
            .I(N__55242));
    LocalMux I__13591 (
            .O(N__55242),
            .I(comm_length_0));
    CascadeMux I__13590 (
            .O(N__55239),
            .I(N__55236));
    InMux I__13589 (
            .O(N__55236),
            .I(N__55225));
    InMux I__13588 (
            .O(N__55235),
            .I(N__55225));
    InMux I__13587 (
            .O(N__55234),
            .I(N__55220));
    InMux I__13586 (
            .O(N__55233),
            .I(N__55220));
    InMux I__13585 (
            .O(N__55232),
            .I(N__55205));
    InMux I__13584 (
            .O(N__55231),
            .I(N__55200));
    InMux I__13583 (
            .O(N__55230),
            .I(N__55200));
    LocalMux I__13582 (
            .O(N__55225),
            .I(N__55195));
    LocalMux I__13581 (
            .O(N__55220),
            .I(N__55195));
    InMux I__13580 (
            .O(N__55219),
            .I(N__55190));
    InMux I__13579 (
            .O(N__55218),
            .I(N__55190));
    InMux I__13578 (
            .O(N__55217),
            .I(N__55184));
    InMux I__13577 (
            .O(N__55216),
            .I(N__55177));
    InMux I__13576 (
            .O(N__55215),
            .I(N__55177));
    InMux I__13575 (
            .O(N__55214),
            .I(N__55177));
    CascadeMux I__13574 (
            .O(N__55213),
            .I(N__55166));
    CascadeMux I__13573 (
            .O(N__55212),
            .I(N__55142));
    CascadeMux I__13572 (
            .O(N__55211),
            .I(N__55137));
    CascadeMux I__13571 (
            .O(N__55210),
            .I(N__55133));
    CascadeMux I__13570 (
            .O(N__55209),
            .I(N__55129));
    InMux I__13569 (
            .O(N__55208),
            .I(N__55126));
    LocalMux I__13568 (
            .O(N__55205),
            .I(N__55116));
    LocalMux I__13567 (
            .O(N__55200),
            .I(N__55116));
    Span4Mux_v I__13566 (
            .O(N__55195),
            .I(N__55116));
    LocalMux I__13565 (
            .O(N__55190),
            .I(N__55116));
    InMux I__13564 (
            .O(N__55189),
            .I(N__55109));
    InMux I__13563 (
            .O(N__55188),
            .I(N__55109));
    InMux I__13562 (
            .O(N__55187),
            .I(N__55109));
    LocalMux I__13561 (
            .O(N__55184),
            .I(N__55104));
    LocalMux I__13560 (
            .O(N__55177),
            .I(N__55104));
    InMux I__13559 (
            .O(N__55176),
            .I(N__55101));
    InMux I__13558 (
            .O(N__55175),
            .I(N__55098));
    InMux I__13557 (
            .O(N__55174),
            .I(N__55095));
    InMux I__13556 (
            .O(N__55173),
            .I(N__55092));
    InMux I__13555 (
            .O(N__55172),
            .I(N__55085));
    InMux I__13554 (
            .O(N__55171),
            .I(N__55085));
    InMux I__13553 (
            .O(N__55170),
            .I(N__55085));
    InMux I__13552 (
            .O(N__55169),
            .I(N__55082));
    InMux I__13551 (
            .O(N__55166),
            .I(N__55071));
    InMux I__13550 (
            .O(N__55165),
            .I(N__55071));
    InMux I__13549 (
            .O(N__55164),
            .I(N__55071));
    InMux I__13548 (
            .O(N__55163),
            .I(N__55071));
    InMux I__13547 (
            .O(N__55162),
            .I(N__55071));
    InMux I__13546 (
            .O(N__55161),
            .I(N__55066));
    InMux I__13545 (
            .O(N__55160),
            .I(N__55066));
    InMux I__13544 (
            .O(N__55159),
            .I(N__55063));
    InMux I__13543 (
            .O(N__55158),
            .I(N__55060));
    InMux I__13542 (
            .O(N__55157),
            .I(N__55053));
    InMux I__13541 (
            .O(N__55156),
            .I(N__55050));
    InMux I__13540 (
            .O(N__55155),
            .I(N__55047));
    InMux I__13539 (
            .O(N__55154),
            .I(N__55042));
    InMux I__13538 (
            .O(N__55153),
            .I(N__55042));
    InMux I__13537 (
            .O(N__55152),
            .I(N__55037));
    InMux I__13536 (
            .O(N__55151),
            .I(N__55037));
    InMux I__13535 (
            .O(N__55150),
            .I(N__55029));
    InMux I__13534 (
            .O(N__55149),
            .I(N__55029));
    InMux I__13533 (
            .O(N__55148),
            .I(N__55026));
    CascadeMux I__13532 (
            .O(N__55147),
            .I(N__55023));
    CascadeMux I__13531 (
            .O(N__55146),
            .I(N__55019));
    InMux I__13530 (
            .O(N__55145),
            .I(N__55012));
    InMux I__13529 (
            .O(N__55142),
            .I(N__55012));
    InMux I__13528 (
            .O(N__55141),
            .I(N__55012));
    InMux I__13527 (
            .O(N__55140),
            .I(N__55009));
    InMux I__13526 (
            .O(N__55137),
            .I(N__55006));
    InMux I__13525 (
            .O(N__55136),
            .I(N__55003));
    InMux I__13524 (
            .O(N__55133),
            .I(N__54996));
    InMux I__13523 (
            .O(N__55132),
            .I(N__54996));
    InMux I__13522 (
            .O(N__55129),
            .I(N__54996));
    LocalMux I__13521 (
            .O(N__55126),
            .I(N__54993));
    InMux I__13520 (
            .O(N__55125),
            .I(N__54990));
    Span4Mux_v I__13519 (
            .O(N__55116),
            .I(N__54985));
    LocalMux I__13518 (
            .O(N__55109),
            .I(N__54985));
    Span4Mux_v I__13517 (
            .O(N__55104),
            .I(N__54980));
    LocalMux I__13516 (
            .O(N__55101),
            .I(N__54980));
    LocalMux I__13515 (
            .O(N__55098),
            .I(N__54975));
    LocalMux I__13514 (
            .O(N__55095),
            .I(N__54968));
    LocalMux I__13513 (
            .O(N__55092),
            .I(N__54968));
    LocalMux I__13512 (
            .O(N__55085),
            .I(N__54968));
    LocalMux I__13511 (
            .O(N__55082),
            .I(N__54965));
    LocalMux I__13510 (
            .O(N__55071),
            .I(N__54962));
    LocalMux I__13509 (
            .O(N__55066),
            .I(N__54959));
    LocalMux I__13508 (
            .O(N__55063),
            .I(N__54956));
    LocalMux I__13507 (
            .O(N__55060),
            .I(N__54953));
    InMux I__13506 (
            .O(N__55059),
            .I(N__54950));
    InMux I__13505 (
            .O(N__55058),
            .I(N__54947));
    InMux I__13504 (
            .O(N__55057),
            .I(N__54944));
    InMux I__13503 (
            .O(N__55056),
            .I(N__54941));
    LocalMux I__13502 (
            .O(N__55053),
            .I(N__54930));
    LocalMux I__13501 (
            .O(N__55050),
            .I(N__54930));
    LocalMux I__13500 (
            .O(N__55047),
            .I(N__54930));
    LocalMux I__13499 (
            .O(N__55042),
            .I(N__54930));
    LocalMux I__13498 (
            .O(N__55037),
            .I(N__54930));
    InMux I__13497 (
            .O(N__55036),
            .I(N__54925));
    InMux I__13496 (
            .O(N__55035),
            .I(N__54925));
    InMux I__13495 (
            .O(N__55034),
            .I(N__54922));
    LocalMux I__13494 (
            .O(N__55029),
            .I(N__54917));
    LocalMux I__13493 (
            .O(N__55026),
            .I(N__54917));
    InMux I__13492 (
            .O(N__55023),
            .I(N__54914));
    InMux I__13491 (
            .O(N__55022),
            .I(N__54910));
    InMux I__13490 (
            .O(N__55019),
            .I(N__54907));
    LocalMux I__13489 (
            .O(N__55012),
            .I(N__54904));
    LocalMux I__13488 (
            .O(N__55009),
            .I(N__54895));
    LocalMux I__13487 (
            .O(N__55006),
            .I(N__54895));
    LocalMux I__13486 (
            .O(N__55003),
            .I(N__54895));
    LocalMux I__13485 (
            .O(N__54996),
            .I(N__54895));
    Span4Mux_v I__13484 (
            .O(N__54993),
            .I(N__54892));
    LocalMux I__13483 (
            .O(N__54990),
            .I(N__54885));
    Span4Mux_h I__13482 (
            .O(N__54985),
            .I(N__54885));
    Span4Mux_v I__13481 (
            .O(N__54980),
            .I(N__54885));
    InMux I__13480 (
            .O(N__54979),
            .I(N__54879));
    InMux I__13479 (
            .O(N__54978),
            .I(N__54879));
    Span4Mux_v I__13478 (
            .O(N__54975),
            .I(N__54874));
    Span4Mux_v I__13477 (
            .O(N__54968),
            .I(N__54874));
    Span4Mux_v I__13476 (
            .O(N__54965),
            .I(N__54869));
    Span4Mux_v I__13475 (
            .O(N__54962),
            .I(N__54869));
    Span4Mux_v I__13474 (
            .O(N__54959),
            .I(N__54865));
    Span4Mux_v I__13473 (
            .O(N__54956),
            .I(N__54860));
    Span4Mux_v I__13472 (
            .O(N__54953),
            .I(N__54860));
    LocalMux I__13471 (
            .O(N__54950),
            .I(N__54857));
    LocalMux I__13470 (
            .O(N__54947),
            .I(N__54852));
    LocalMux I__13469 (
            .O(N__54944),
            .I(N__54852));
    LocalMux I__13468 (
            .O(N__54941),
            .I(N__54849));
    Span4Mux_v I__13467 (
            .O(N__54930),
            .I(N__54838));
    LocalMux I__13466 (
            .O(N__54925),
            .I(N__54838));
    LocalMux I__13465 (
            .O(N__54922),
            .I(N__54838));
    Span4Mux_h I__13464 (
            .O(N__54917),
            .I(N__54838));
    LocalMux I__13463 (
            .O(N__54914),
            .I(N__54838));
    InMux I__13462 (
            .O(N__54913),
            .I(N__54832));
    LocalMux I__13461 (
            .O(N__54910),
            .I(N__54827));
    LocalMux I__13460 (
            .O(N__54907),
            .I(N__54827));
    Span4Mux_h I__13459 (
            .O(N__54904),
            .I(N__54818));
    Span4Mux_v I__13458 (
            .O(N__54895),
            .I(N__54818));
    Span4Mux_v I__13457 (
            .O(N__54892),
            .I(N__54818));
    Span4Mux_v I__13456 (
            .O(N__54885),
            .I(N__54818));
    InMux I__13455 (
            .O(N__54884),
            .I(N__54815));
    LocalMux I__13454 (
            .O(N__54879),
            .I(N__54808));
    Span4Mux_h I__13453 (
            .O(N__54874),
            .I(N__54808));
    Span4Mux_h I__13452 (
            .O(N__54869),
            .I(N__54808));
    InMux I__13451 (
            .O(N__54868),
            .I(N__54805));
    Span4Mux_h I__13450 (
            .O(N__54865),
            .I(N__54800));
    Span4Mux_h I__13449 (
            .O(N__54860),
            .I(N__54800));
    Span4Mux_h I__13448 (
            .O(N__54857),
            .I(N__54791));
    Span4Mux_h I__13447 (
            .O(N__54852),
            .I(N__54791));
    Span4Mux_v I__13446 (
            .O(N__54849),
            .I(N__54791));
    Span4Mux_h I__13445 (
            .O(N__54838),
            .I(N__54791));
    InMux I__13444 (
            .O(N__54837),
            .I(N__54784));
    InMux I__13443 (
            .O(N__54836),
            .I(N__54784));
    InMux I__13442 (
            .O(N__54835),
            .I(N__54784));
    LocalMux I__13441 (
            .O(N__54832),
            .I(comm_cmd_1));
    Odrv12 I__13440 (
            .O(N__54827),
            .I(comm_cmd_1));
    Odrv4 I__13439 (
            .O(N__54818),
            .I(comm_cmd_1));
    LocalMux I__13438 (
            .O(N__54815),
            .I(comm_cmd_1));
    Odrv4 I__13437 (
            .O(N__54808),
            .I(comm_cmd_1));
    LocalMux I__13436 (
            .O(N__54805),
            .I(comm_cmd_1));
    Odrv4 I__13435 (
            .O(N__54800),
            .I(comm_cmd_1));
    Odrv4 I__13434 (
            .O(N__54791),
            .I(comm_cmd_1));
    LocalMux I__13433 (
            .O(N__54784),
            .I(comm_cmd_1));
    InMux I__13432 (
            .O(N__54765),
            .I(N__54750));
    InMux I__13431 (
            .O(N__54764),
            .I(N__54741));
    InMux I__13430 (
            .O(N__54763),
            .I(N__54738));
    InMux I__13429 (
            .O(N__54762),
            .I(N__54733));
    InMux I__13428 (
            .O(N__54761),
            .I(N__54733));
    InMux I__13427 (
            .O(N__54760),
            .I(N__54728));
    InMux I__13426 (
            .O(N__54759),
            .I(N__54728));
    InMux I__13425 (
            .O(N__54758),
            .I(N__54723));
    InMux I__13424 (
            .O(N__54757),
            .I(N__54723));
    InMux I__13423 (
            .O(N__54756),
            .I(N__54720));
    InMux I__13422 (
            .O(N__54755),
            .I(N__54716));
    InMux I__13421 (
            .O(N__54754),
            .I(N__54713));
    InMux I__13420 (
            .O(N__54753),
            .I(N__54708));
    LocalMux I__13419 (
            .O(N__54750),
            .I(N__54703));
    InMux I__13418 (
            .O(N__54749),
            .I(N__54698));
    InMux I__13417 (
            .O(N__54748),
            .I(N__54698));
    InMux I__13416 (
            .O(N__54747),
            .I(N__54688));
    InMux I__13415 (
            .O(N__54746),
            .I(N__54683));
    InMux I__13414 (
            .O(N__54745),
            .I(N__54680));
    InMux I__13413 (
            .O(N__54744),
            .I(N__54677));
    LocalMux I__13412 (
            .O(N__54741),
            .I(N__54672));
    LocalMux I__13411 (
            .O(N__54738),
            .I(N__54672));
    LocalMux I__13410 (
            .O(N__54733),
            .I(N__54665));
    LocalMux I__13409 (
            .O(N__54728),
            .I(N__54665));
    LocalMux I__13408 (
            .O(N__54723),
            .I(N__54665));
    LocalMux I__13407 (
            .O(N__54720),
            .I(N__54662));
    InMux I__13406 (
            .O(N__54719),
            .I(N__54659));
    LocalMux I__13405 (
            .O(N__54716),
            .I(N__54654));
    LocalMux I__13404 (
            .O(N__54713),
            .I(N__54654));
    InMux I__13403 (
            .O(N__54712),
            .I(N__54648));
    InMux I__13402 (
            .O(N__54711),
            .I(N__54648));
    LocalMux I__13401 (
            .O(N__54708),
            .I(N__54645));
    InMux I__13400 (
            .O(N__54707),
            .I(N__54641));
    InMux I__13399 (
            .O(N__54706),
            .I(N__54638));
    Span4Mux_h I__13398 (
            .O(N__54703),
            .I(N__54635));
    LocalMux I__13397 (
            .O(N__54698),
            .I(N__54632));
    InMux I__13396 (
            .O(N__54697),
            .I(N__54628));
    InMux I__13395 (
            .O(N__54696),
            .I(N__54625));
    InMux I__13394 (
            .O(N__54695),
            .I(N__54622));
    InMux I__13393 (
            .O(N__54694),
            .I(N__54619));
    InMux I__13392 (
            .O(N__54693),
            .I(N__54614));
    InMux I__13391 (
            .O(N__54692),
            .I(N__54614));
    InMux I__13390 (
            .O(N__54691),
            .I(N__54611));
    LocalMux I__13389 (
            .O(N__54688),
            .I(N__54608));
    InMux I__13388 (
            .O(N__54687),
            .I(N__54603));
    InMux I__13387 (
            .O(N__54686),
            .I(N__54603));
    LocalMux I__13386 (
            .O(N__54683),
            .I(N__54598));
    LocalMux I__13385 (
            .O(N__54680),
            .I(N__54595));
    LocalMux I__13384 (
            .O(N__54677),
            .I(N__54588));
    Span4Mux_v I__13383 (
            .O(N__54672),
            .I(N__54588));
    Span4Mux_v I__13382 (
            .O(N__54665),
            .I(N__54588));
    Span4Mux_v I__13381 (
            .O(N__54662),
            .I(N__54585));
    LocalMux I__13380 (
            .O(N__54659),
            .I(N__54582));
    Span4Mux_h I__13379 (
            .O(N__54654),
            .I(N__54579));
    InMux I__13378 (
            .O(N__54653),
            .I(N__54576));
    LocalMux I__13377 (
            .O(N__54648),
            .I(N__54573));
    Sp12to4 I__13376 (
            .O(N__54645),
            .I(N__54570));
    InMux I__13375 (
            .O(N__54644),
            .I(N__54566));
    LocalMux I__13374 (
            .O(N__54641),
            .I(N__54563));
    LocalMux I__13373 (
            .O(N__54638),
            .I(N__54558));
    Span4Mux_v I__13372 (
            .O(N__54635),
            .I(N__54558));
    Span4Mux_h I__13371 (
            .O(N__54632),
            .I(N__54555));
    InMux I__13370 (
            .O(N__54631),
            .I(N__54551));
    LocalMux I__13369 (
            .O(N__54628),
            .I(N__54546));
    LocalMux I__13368 (
            .O(N__54625),
            .I(N__54546));
    LocalMux I__13367 (
            .O(N__54622),
            .I(N__54539));
    LocalMux I__13366 (
            .O(N__54619),
            .I(N__54539));
    LocalMux I__13365 (
            .O(N__54614),
            .I(N__54539));
    LocalMux I__13364 (
            .O(N__54611),
            .I(N__54532));
    Span4Mux_h I__13363 (
            .O(N__54608),
            .I(N__54532));
    LocalMux I__13362 (
            .O(N__54603),
            .I(N__54532));
    InMux I__13361 (
            .O(N__54602),
            .I(N__54529));
    InMux I__13360 (
            .O(N__54601),
            .I(N__54526));
    Span4Mux_h I__13359 (
            .O(N__54598),
            .I(N__54517));
    Span4Mux_v I__13358 (
            .O(N__54595),
            .I(N__54517));
    Span4Mux_h I__13357 (
            .O(N__54588),
            .I(N__54517));
    Span4Mux_v I__13356 (
            .O(N__54585),
            .I(N__54517));
    Span4Mux_h I__13355 (
            .O(N__54582),
            .I(N__54512));
    Span4Mux_v I__13354 (
            .O(N__54579),
            .I(N__54512));
    LocalMux I__13353 (
            .O(N__54576),
            .I(N__54505));
    Span12Mux_v I__13352 (
            .O(N__54573),
            .I(N__54505));
    Span12Mux_v I__13351 (
            .O(N__54570),
            .I(N__54505));
    InMux I__13350 (
            .O(N__54569),
            .I(N__54502));
    LocalMux I__13349 (
            .O(N__54566),
            .I(N__54493));
    Span4Mux_v I__13348 (
            .O(N__54563),
            .I(N__54493));
    Span4Mux_h I__13347 (
            .O(N__54558),
            .I(N__54493));
    Span4Mux_h I__13346 (
            .O(N__54555),
            .I(N__54493));
    InMux I__13345 (
            .O(N__54554),
            .I(N__54490));
    LocalMux I__13344 (
            .O(N__54551),
            .I(N__54481));
    Span4Mux_v I__13343 (
            .O(N__54546),
            .I(N__54481));
    Span4Mux_v I__13342 (
            .O(N__54539),
            .I(N__54481));
    Span4Mux_v I__13341 (
            .O(N__54532),
            .I(N__54481));
    LocalMux I__13340 (
            .O(N__54529),
            .I(N__54478));
    LocalMux I__13339 (
            .O(N__54526),
            .I(comm_cmd_3));
    Odrv4 I__13338 (
            .O(N__54517),
            .I(comm_cmd_3));
    Odrv4 I__13337 (
            .O(N__54512),
            .I(comm_cmd_3));
    Odrv12 I__13336 (
            .O(N__54505),
            .I(comm_cmd_3));
    LocalMux I__13335 (
            .O(N__54502),
            .I(comm_cmd_3));
    Odrv4 I__13334 (
            .O(N__54493),
            .I(comm_cmd_3));
    LocalMux I__13333 (
            .O(N__54490),
            .I(comm_cmd_3));
    Odrv4 I__13332 (
            .O(N__54481),
            .I(comm_cmd_3));
    Odrv12 I__13331 (
            .O(N__54478),
            .I(comm_cmd_3));
    CascadeMux I__13330 (
            .O(N__54459),
            .I(N__54456));
    InMux I__13329 (
            .O(N__54456),
            .I(N__54453));
    LocalMux I__13328 (
            .O(N__54453),
            .I(N__54450));
    Span4Mux_h I__13327 (
            .O(N__54450),
            .I(N__54446));
    InMux I__13326 (
            .O(N__54449),
            .I(N__54443));
    Odrv4 I__13325 (
            .O(N__54446),
            .I(comm_length_1));
    LocalMux I__13324 (
            .O(N__54443),
            .I(comm_length_1));
    ClkMux I__13323 (
            .O(N__54438),
            .I(N__53928));
    ClkMux I__13322 (
            .O(N__54437),
            .I(N__53928));
    ClkMux I__13321 (
            .O(N__54436),
            .I(N__53928));
    ClkMux I__13320 (
            .O(N__54435),
            .I(N__53928));
    ClkMux I__13319 (
            .O(N__54434),
            .I(N__53928));
    ClkMux I__13318 (
            .O(N__54433),
            .I(N__53928));
    ClkMux I__13317 (
            .O(N__54432),
            .I(N__53928));
    ClkMux I__13316 (
            .O(N__54431),
            .I(N__53928));
    ClkMux I__13315 (
            .O(N__54430),
            .I(N__53928));
    ClkMux I__13314 (
            .O(N__54429),
            .I(N__53928));
    ClkMux I__13313 (
            .O(N__54428),
            .I(N__53928));
    ClkMux I__13312 (
            .O(N__54427),
            .I(N__53928));
    ClkMux I__13311 (
            .O(N__54426),
            .I(N__53928));
    ClkMux I__13310 (
            .O(N__54425),
            .I(N__53928));
    ClkMux I__13309 (
            .O(N__54424),
            .I(N__53928));
    ClkMux I__13308 (
            .O(N__54423),
            .I(N__53928));
    ClkMux I__13307 (
            .O(N__54422),
            .I(N__53928));
    ClkMux I__13306 (
            .O(N__54421),
            .I(N__53928));
    ClkMux I__13305 (
            .O(N__54420),
            .I(N__53928));
    ClkMux I__13304 (
            .O(N__54419),
            .I(N__53928));
    ClkMux I__13303 (
            .O(N__54418),
            .I(N__53928));
    ClkMux I__13302 (
            .O(N__54417),
            .I(N__53928));
    ClkMux I__13301 (
            .O(N__54416),
            .I(N__53928));
    ClkMux I__13300 (
            .O(N__54415),
            .I(N__53928));
    ClkMux I__13299 (
            .O(N__54414),
            .I(N__53928));
    ClkMux I__13298 (
            .O(N__54413),
            .I(N__53928));
    ClkMux I__13297 (
            .O(N__54412),
            .I(N__53928));
    ClkMux I__13296 (
            .O(N__54411),
            .I(N__53928));
    ClkMux I__13295 (
            .O(N__54410),
            .I(N__53928));
    ClkMux I__13294 (
            .O(N__54409),
            .I(N__53928));
    ClkMux I__13293 (
            .O(N__54408),
            .I(N__53928));
    ClkMux I__13292 (
            .O(N__54407),
            .I(N__53928));
    ClkMux I__13291 (
            .O(N__54406),
            .I(N__53928));
    ClkMux I__13290 (
            .O(N__54405),
            .I(N__53928));
    ClkMux I__13289 (
            .O(N__54404),
            .I(N__53928));
    ClkMux I__13288 (
            .O(N__54403),
            .I(N__53928));
    ClkMux I__13287 (
            .O(N__54402),
            .I(N__53928));
    ClkMux I__13286 (
            .O(N__54401),
            .I(N__53928));
    ClkMux I__13285 (
            .O(N__54400),
            .I(N__53928));
    ClkMux I__13284 (
            .O(N__54399),
            .I(N__53928));
    ClkMux I__13283 (
            .O(N__54398),
            .I(N__53928));
    ClkMux I__13282 (
            .O(N__54397),
            .I(N__53928));
    ClkMux I__13281 (
            .O(N__54396),
            .I(N__53928));
    ClkMux I__13280 (
            .O(N__54395),
            .I(N__53928));
    ClkMux I__13279 (
            .O(N__54394),
            .I(N__53928));
    ClkMux I__13278 (
            .O(N__54393),
            .I(N__53928));
    ClkMux I__13277 (
            .O(N__54392),
            .I(N__53928));
    ClkMux I__13276 (
            .O(N__54391),
            .I(N__53928));
    ClkMux I__13275 (
            .O(N__54390),
            .I(N__53928));
    ClkMux I__13274 (
            .O(N__54389),
            .I(N__53928));
    ClkMux I__13273 (
            .O(N__54388),
            .I(N__53928));
    ClkMux I__13272 (
            .O(N__54387),
            .I(N__53928));
    ClkMux I__13271 (
            .O(N__54386),
            .I(N__53928));
    ClkMux I__13270 (
            .O(N__54385),
            .I(N__53928));
    ClkMux I__13269 (
            .O(N__54384),
            .I(N__53928));
    ClkMux I__13268 (
            .O(N__54383),
            .I(N__53928));
    ClkMux I__13267 (
            .O(N__54382),
            .I(N__53928));
    ClkMux I__13266 (
            .O(N__54381),
            .I(N__53928));
    ClkMux I__13265 (
            .O(N__54380),
            .I(N__53928));
    ClkMux I__13264 (
            .O(N__54379),
            .I(N__53928));
    ClkMux I__13263 (
            .O(N__54378),
            .I(N__53928));
    ClkMux I__13262 (
            .O(N__54377),
            .I(N__53928));
    ClkMux I__13261 (
            .O(N__54376),
            .I(N__53928));
    ClkMux I__13260 (
            .O(N__54375),
            .I(N__53928));
    ClkMux I__13259 (
            .O(N__54374),
            .I(N__53928));
    ClkMux I__13258 (
            .O(N__54373),
            .I(N__53928));
    ClkMux I__13257 (
            .O(N__54372),
            .I(N__53928));
    ClkMux I__13256 (
            .O(N__54371),
            .I(N__53928));
    ClkMux I__13255 (
            .O(N__54370),
            .I(N__53928));
    ClkMux I__13254 (
            .O(N__54369),
            .I(N__53928));
    ClkMux I__13253 (
            .O(N__54368),
            .I(N__53928));
    ClkMux I__13252 (
            .O(N__54367),
            .I(N__53928));
    ClkMux I__13251 (
            .O(N__54366),
            .I(N__53928));
    ClkMux I__13250 (
            .O(N__54365),
            .I(N__53928));
    ClkMux I__13249 (
            .O(N__54364),
            .I(N__53928));
    ClkMux I__13248 (
            .O(N__54363),
            .I(N__53928));
    ClkMux I__13247 (
            .O(N__54362),
            .I(N__53928));
    ClkMux I__13246 (
            .O(N__54361),
            .I(N__53928));
    ClkMux I__13245 (
            .O(N__54360),
            .I(N__53928));
    ClkMux I__13244 (
            .O(N__54359),
            .I(N__53928));
    ClkMux I__13243 (
            .O(N__54358),
            .I(N__53928));
    ClkMux I__13242 (
            .O(N__54357),
            .I(N__53928));
    ClkMux I__13241 (
            .O(N__54356),
            .I(N__53928));
    ClkMux I__13240 (
            .O(N__54355),
            .I(N__53928));
    ClkMux I__13239 (
            .O(N__54354),
            .I(N__53928));
    ClkMux I__13238 (
            .O(N__54353),
            .I(N__53928));
    ClkMux I__13237 (
            .O(N__54352),
            .I(N__53928));
    ClkMux I__13236 (
            .O(N__54351),
            .I(N__53928));
    ClkMux I__13235 (
            .O(N__54350),
            .I(N__53928));
    ClkMux I__13234 (
            .O(N__54349),
            .I(N__53928));
    ClkMux I__13233 (
            .O(N__54348),
            .I(N__53928));
    ClkMux I__13232 (
            .O(N__54347),
            .I(N__53928));
    ClkMux I__13231 (
            .O(N__54346),
            .I(N__53928));
    ClkMux I__13230 (
            .O(N__54345),
            .I(N__53928));
    ClkMux I__13229 (
            .O(N__54344),
            .I(N__53928));
    ClkMux I__13228 (
            .O(N__54343),
            .I(N__53928));
    ClkMux I__13227 (
            .O(N__54342),
            .I(N__53928));
    ClkMux I__13226 (
            .O(N__54341),
            .I(N__53928));
    ClkMux I__13225 (
            .O(N__54340),
            .I(N__53928));
    ClkMux I__13224 (
            .O(N__54339),
            .I(N__53928));
    ClkMux I__13223 (
            .O(N__54338),
            .I(N__53928));
    ClkMux I__13222 (
            .O(N__54337),
            .I(N__53928));
    ClkMux I__13221 (
            .O(N__54336),
            .I(N__53928));
    ClkMux I__13220 (
            .O(N__54335),
            .I(N__53928));
    ClkMux I__13219 (
            .O(N__54334),
            .I(N__53928));
    ClkMux I__13218 (
            .O(N__54333),
            .I(N__53928));
    ClkMux I__13217 (
            .O(N__54332),
            .I(N__53928));
    ClkMux I__13216 (
            .O(N__54331),
            .I(N__53928));
    ClkMux I__13215 (
            .O(N__54330),
            .I(N__53928));
    ClkMux I__13214 (
            .O(N__54329),
            .I(N__53928));
    ClkMux I__13213 (
            .O(N__54328),
            .I(N__53928));
    ClkMux I__13212 (
            .O(N__54327),
            .I(N__53928));
    ClkMux I__13211 (
            .O(N__54326),
            .I(N__53928));
    ClkMux I__13210 (
            .O(N__54325),
            .I(N__53928));
    ClkMux I__13209 (
            .O(N__54324),
            .I(N__53928));
    ClkMux I__13208 (
            .O(N__54323),
            .I(N__53928));
    ClkMux I__13207 (
            .O(N__54322),
            .I(N__53928));
    ClkMux I__13206 (
            .O(N__54321),
            .I(N__53928));
    ClkMux I__13205 (
            .O(N__54320),
            .I(N__53928));
    ClkMux I__13204 (
            .O(N__54319),
            .I(N__53928));
    ClkMux I__13203 (
            .O(N__54318),
            .I(N__53928));
    ClkMux I__13202 (
            .O(N__54317),
            .I(N__53928));
    ClkMux I__13201 (
            .O(N__54316),
            .I(N__53928));
    ClkMux I__13200 (
            .O(N__54315),
            .I(N__53928));
    ClkMux I__13199 (
            .O(N__54314),
            .I(N__53928));
    ClkMux I__13198 (
            .O(N__54313),
            .I(N__53928));
    ClkMux I__13197 (
            .O(N__54312),
            .I(N__53928));
    ClkMux I__13196 (
            .O(N__54311),
            .I(N__53928));
    ClkMux I__13195 (
            .O(N__54310),
            .I(N__53928));
    ClkMux I__13194 (
            .O(N__54309),
            .I(N__53928));
    ClkMux I__13193 (
            .O(N__54308),
            .I(N__53928));
    ClkMux I__13192 (
            .O(N__54307),
            .I(N__53928));
    ClkMux I__13191 (
            .O(N__54306),
            .I(N__53928));
    ClkMux I__13190 (
            .O(N__54305),
            .I(N__53928));
    ClkMux I__13189 (
            .O(N__54304),
            .I(N__53928));
    ClkMux I__13188 (
            .O(N__54303),
            .I(N__53928));
    ClkMux I__13187 (
            .O(N__54302),
            .I(N__53928));
    ClkMux I__13186 (
            .O(N__54301),
            .I(N__53928));
    ClkMux I__13185 (
            .O(N__54300),
            .I(N__53928));
    ClkMux I__13184 (
            .O(N__54299),
            .I(N__53928));
    ClkMux I__13183 (
            .O(N__54298),
            .I(N__53928));
    ClkMux I__13182 (
            .O(N__54297),
            .I(N__53928));
    ClkMux I__13181 (
            .O(N__54296),
            .I(N__53928));
    ClkMux I__13180 (
            .O(N__54295),
            .I(N__53928));
    ClkMux I__13179 (
            .O(N__54294),
            .I(N__53928));
    ClkMux I__13178 (
            .O(N__54293),
            .I(N__53928));
    ClkMux I__13177 (
            .O(N__54292),
            .I(N__53928));
    ClkMux I__13176 (
            .O(N__54291),
            .I(N__53928));
    ClkMux I__13175 (
            .O(N__54290),
            .I(N__53928));
    ClkMux I__13174 (
            .O(N__54289),
            .I(N__53928));
    ClkMux I__13173 (
            .O(N__54288),
            .I(N__53928));
    ClkMux I__13172 (
            .O(N__54287),
            .I(N__53928));
    ClkMux I__13171 (
            .O(N__54286),
            .I(N__53928));
    ClkMux I__13170 (
            .O(N__54285),
            .I(N__53928));
    ClkMux I__13169 (
            .O(N__54284),
            .I(N__53928));
    ClkMux I__13168 (
            .O(N__54283),
            .I(N__53928));
    ClkMux I__13167 (
            .O(N__54282),
            .I(N__53928));
    ClkMux I__13166 (
            .O(N__54281),
            .I(N__53928));
    ClkMux I__13165 (
            .O(N__54280),
            .I(N__53928));
    ClkMux I__13164 (
            .O(N__54279),
            .I(N__53928));
    ClkMux I__13163 (
            .O(N__54278),
            .I(N__53928));
    ClkMux I__13162 (
            .O(N__54277),
            .I(N__53928));
    ClkMux I__13161 (
            .O(N__54276),
            .I(N__53928));
    ClkMux I__13160 (
            .O(N__54275),
            .I(N__53928));
    ClkMux I__13159 (
            .O(N__54274),
            .I(N__53928));
    ClkMux I__13158 (
            .O(N__54273),
            .I(N__53928));
    ClkMux I__13157 (
            .O(N__54272),
            .I(N__53928));
    ClkMux I__13156 (
            .O(N__54271),
            .I(N__53928));
    ClkMux I__13155 (
            .O(N__54270),
            .I(N__53928));
    ClkMux I__13154 (
            .O(N__54269),
            .I(N__53928));
    GlobalMux I__13153 (
            .O(N__53928),
            .I(clk_32MHz));
    CEMux I__13152 (
            .O(N__53925),
            .I(N__53921));
    InMux I__13151 (
            .O(N__53924),
            .I(N__53918));
    LocalMux I__13150 (
            .O(N__53921),
            .I(N__53914));
    LocalMux I__13149 (
            .O(N__53918),
            .I(N__53911));
    InMux I__13148 (
            .O(N__53917),
            .I(N__53908));
    Odrv4 I__13147 (
            .O(N__53914),
            .I(n11860));
    Odrv4 I__13146 (
            .O(N__53911),
            .I(n11860));
    LocalMux I__13145 (
            .O(N__53908),
            .I(n11860));
    SRMux I__13144 (
            .O(N__53901),
            .I(N__53898));
    LocalMux I__13143 (
            .O(N__53898),
            .I(n14655));
    CascadeMux I__13142 (
            .O(N__53895),
            .I(N__53892));
    InMux I__13141 (
            .O(N__53892),
            .I(N__53889));
    LocalMux I__13140 (
            .O(N__53889),
            .I(N__53886));
    Odrv4 I__13139 (
            .O(N__53886),
            .I(buf_data_iac_12));
    InMux I__13138 (
            .O(N__53883),
            .I(N__53880));
    LocalMux I__13137 (
            .O(N__53880),
            .I(N__53877));
    Odrv4 I__13136 (
            .O(N__53877),
            .I(n21451));
    InMux I__13135 (
            .O(N__53874),
            .I(N__53871));
    LocalMux I__13134 (
            .O(N__53871),
            .I(N__53868));
    Odrv4 I__13133 (
            .O(N__53868),
            .I(buf_data_iac_18));
    CascadeMux I__13132 (
            .O(N__53865),
            .I(N__53862));
    InMux I__13131 (
            .O(N__53862),
            .I(N__53859));
    LocalMux I__13130 (
            .O(N__53859),
            .I(N__53856));
    Span4Mux_h I__13129 (
            .O(N__53856),
            .I(N__53853));
    Odrv4 I__13128 (
            .O(N__53853),
            .I(n21151));
    InMux I__13127 (
            .O(N__53850),
            .I(N__53847));
    LocalMux I__13126 (
            .O(N__53847),
            .I(N__53844));
    Span12Mux_h I__13125 (
            .O(N__53844),
            .I(N__53841));
    Odrv12 I__13124 (
            .O(N__53841),
            .I(n16_adj_1496));
    InMux I__13123 (
            .O(N__53838),
            .I(N__53835));
    LocalMux I__13122 (
            .O(N__53835),
            .I(n22399));
    InMux I__13121 (
            .O(N__53832),
            .I(N__53828));
    CascadeMux I__13120 (
            .O(N__53831),
            .I(N__53825));
    LocalMux I__13119 (
            .O(N__53828),
            .I(N__53822));
    InMux I__13118 (
            .O(N__53825),
            .I(N__53819));
    Span4Mux_h I__13117 (
            .O(N__53822),
            .I(N__53814));
    LocalMux I__13116 (
            .O(N__53819),
            .I(N__53814));
    Span4Mux_v I__13115 (
            .O(N__53814),
            .I(N__53810));
    InMux I__13114 (
            .O(N__53813),
            .I(N__53807));
    Span4Mux_h I__13113 (
            .O(N__53810),
            .I(N__53804));
    LocalMux I__13112 (
            .O(N__53807),
            .I(buf_adcdata_iac_13));
    Odrv4 I__13111 (
            .O(N__53804),
            .I(buf_adcdata_iac_13));
    InMux I__13110 (
            .O(N__53799),
            .I(N__53772));
    InMux I__13109 (
            .O(N__53798),
            .I(N__53772));
    InMux I__13108 (
            .O(N__53797),
            .I(N__53768));
    CascadeMux I__13107 (
            .O(N__53796),
            .I(N__53758));
    CascadeMux I__13106 (
            .O(N__53795),
            .I(N__53751));
    InMux I__13105 (
            .O(N__53794),
            .I(N__53746));
    InMux I__13104 (
            .O(N__53793),
            .I(N__53739));
    InMux I__13103 (
            .O(N__53792),
            .I(N__53739));
    InMux I__13102 (
            .O(N__53791),
            .I(N__53739));
    InMux I__13101 (
            .O(N__53790),
            .I(N__53730));
    InMux I__13100 (
            .O(N__53789),
            .I(N__53730));
    InMux I__13099 (
            .O(N__53788),
            .I(N__53730));
    InMux I__13098 (
            .O(N__53787),
            .I(N__53730));
    InMux I__13097 (
            .O(N__53786),
            .I(N__53724));
    InMux I__13096 (
            .O(N__53785),
            .I(N__53717));
    InMux I__13095 (
            .O(N__53784),
            .I(N__53710));
    InMux I__13094 (
            .O(N__53783),
            .I(N__53710));
    InMux I__13093 (
            .O(N__53782),
            .I(N__53710));
    InMux I__13092 (
            .O(N__53781),
            .I(N__53707));
    InMux I__13091 (
            .O(N__53780),
            .I(N__53704));
    InMux I__13090 (
            .O(N__53779),
            .I(N__53699));
    InMux I__13089 (
            .O(N__53778),
            .I(N__53699));
    InMux I__13088 (
            .O(N__53777),
            .I(N__53696));
    LocalMux I__13087 (
            .O(N__53772),
            .I(N__53693));
    InMux I__13086 (
            .O(N__53771),
            .I(N__53690));
    LocalMux I__13085 (
            .O(N__53768),
            .I(N__53687));
    InMux I__13084 (
            .O(N__53767),
            .I(N__53684));
    InMux I__13083 (
            .O(N__53766),
            .I(N__53676));
    InMux I__13082 (
            .O(N__53765),
            .I(N__53673));
    InMux I__13081 (
            .O(N__53764),
            .I(N__53659));
    InMux I__13080 (
            .O(N__53763),
            .I(N__53659));
    InMux I__13079 (
            .O(N__53762),
            .I(N__53659));
    InMux I__13078 (
            .O(N__53761),
            .I(N__53654));
    InMux I__13077 (
            .O(N__53758),
            .I(N__53654));
    InMux I__13076 (
            .O(N__53757),
            .I(N__53645));
    InMux I__13075 (
            .O(N__53756),
            .I(N__53645));
    InMux I__13074 (
            .O(N__53755),
            .I(N__53645));
    InMux I__13073 (
            .O(N__53754),
            .I(N__53645));
    InMux I__13072 (
            .O(N__53751),
            .I(N__53642));
    InMux I__13071 (
            .O(N__53750),
            .I(N__53637));
    InMux I__13070 (
            .O(N__53749),
            .I(N__53637));
    LocalMux I__13069 (
            .O(N__53746),
            .I(N__53634));
    LocalMux I__13068 (
            .O(N__53739),
            .I(N__53631));
    LocalMux I__13067 (
            .O(N__53730),
            .I(N__53628));
    InMux I__13066 (
            .O(N__53729),
            .I(N__53621));
    InMux I__13065 (
            .O(N__53728),
            .I(N__53621));
    InMux I__13064 (
            .O(N__53727),
            .I(N__53621));
    LocalMux I__13063 (
            .O(N__53724),
            .I(N__53618));
    InMux I__13062 (
            .O(N__53723),
            .I(N__53615));
    InMux I__13061 (
            .O(N__53722),
            .I(N__53608));
    InMux I__13060 (
            .O(N__53721),
            .I(N__53605));
    InMux I__13059 (
            .O(N__53720),
            .I(N__53602));
    LocalMux I__13058 (
            .O(N__53717),
            .I(N__53597));
    LocalMux I__13057 (
            .O(N__53710),
            .I(N__53597));
    LocalMux I__13056 (
            .O(N__53707),
            .I(N__53590));
    LocalMux I__13055 (
            .O(N__53704),
            .I(N__53590));
    LocalMux I__13054 (
            .O(N__53699),
            .I(N__53590));
    LocalMux I__13053 (
            .O(N__53696),
            .I(N__53585));
    Span4Mux_v I__13052 (
            .O(N__53693),
            .I(N__53585));
    LocalMux I__13051 (
            .O(N__53690),
            .I(N__53580));
    Span4Mux_h I__13050 (
            .O(N__53687),
            .I(N__53580));
    LocalMux I__13049 (
            .O(N__53684),
            .I(N__53577));
    InMux I__13048 (
            .O(N__53683),
            .I(N__53568));
    InMux I__13047 (
            .O(N__53682),
            .I(N__53568));
    InMux I__13046 (
            .O(N__53681),
            .I(N__53568));
    InMux I__13045 (
            .O(N__53680),
            .I(N__53568));
    InMux I__13044 (
            .O(N__53679),
            .I(N__53565));
    LocalMux I__13043 (
            .O(N__53676),
            .I(N__53562));
    LocalMux I__13042 (
            .O(N__53673),
            .I(N__53559));
    InMux I__13041 (
            .O(N__53672),
            .I(N__53556));
    InMux I__13040 (
            .O(N__53671),
            .I(N__53549));
    InMux I__13039 (
            .O(N__53670),
            .I(N__53545));
    InMux I__13038 (
            .O(N__53669),
            .I(N__53536));
    InMux I__13037 (
            .O(N__53668),
            .I(N__53536));
    InMux I__13036 (
            .O(N__53667),
            .I(N__53536));
    InMux I__13035 (
            .O(N__53666),
            .I(N__53536));
    LocalMux I__13034 (
            .O(N__53659),
            .I(N__53529));
    LocalMux I__13033 (
            .O(N__53654),
            .I(N__53529));
    LocalMux I__13032 (
            .O(N__53645),
            .I(N__53529));
    LocalMux I__13031 (
            .O(N__53642),
            .I(N__53526));
    LocalMux I__13030 (
            .O(N__53637),
            .I(N__53523));
    Span4Mux_h I__13029 (
            .O(N__53634),
            .I(N__53520));
    Span4Mux_h I__13028 (
            .O(N__53631),
            .I(N__53513));
    Span4Mux_v I__13027 (
            .O(N__53628),
            .I(N__53513));
    LocalMux I__13026 (
            .O(N__53621),
            .I(N__53513));
    Span4Mux_h I__13025 (
            .O(N__53618),
            .I(N__53510));
    LocalMux I__13024 (
            .O(N__53615),
            .I(N__53507));
    InMux I__13023 (
            .O(N__53614),
            .I(N__53502));
    InMux I__13022 (
            .O(N__53613),
            .I(N__53502));
    InMux I__13021 (
            .O(N__53612),
            .I(N__53499));
    InMux I__13020 (
            .O(N__53611),
            .I(N__53496));
    LocalMux I__13019 (
            .O(N__53608),
            .I(N__53493));
    LocalMux I__13018 (
            .O(N__53605),
            .I(N__53490));
    LocalMux I__13017 (
            .O(N__53602),
            .I(N__53486));
    Span4Mux_h I__13016 (
            .O(N__53597),
            .I(N__53483));
    Span4Mux_h I__13015 (
            .O(N__53590),
            .I(N__53480));
    Span4Mux_h I__13014 (
            .O(N__53585),
            .I(N__53475));
    Span4Mux_v I__13013 (
            .O(N__53580),
            .I(N__53475));
    Span4Mux_h I__13012 (
            .O(N__53577),
            .I(N__53472));
    LocalMux I__13011 (
            .O(N__53568),
            .I(N__53469));
    LocalMux I__13010 (
            .O(N__53565),
            .I(N__53466));
    Span4Mux_h I__13009 (
            .O(N__53562),
            .I(N__53459));
    Span4Mux_v I__13008 (
            .O(N__53559),
            .I(N__53459));
    LocalMux I__13007 (
            .O(N__53556),
            .I(N__53459));
    InMux I__13006 (
            .O(N__53555),
            .I(N__53454));
    InMux I__13005 (
            .O(N__53554),
            .I(N__53447));
    InMux I__13004 (
            .O(N__53553),
            .I(N__53447));
    InMux I__13003 (
            .O(N__53552),
            .I(N__53447));
    LocalMux I__13002 (
            .O(N__53549),
            .I(N__53444));
    InMux I__13001 (
            .O(N__53548),
            .I(N__53441));
    LocalMux I__13000 (
            .O(N__53545),
            .I(N__53430));
    LocalMux I__12999 (
            .O(N__53536),
            .I(N__53430));
    Span4Mux_v I__12998 (
            .O(N__53529),
            .I(N__53430));
    Span4Mux_v I__12997 (
            .O(N__53526),
            .I(N__53430));
    Span4Mux_v I__12996 (
            .O(N__53523),
            .I(N__53430));
    Span4Mux_h I__12995 (
            .O(N__53520),
            .I(N__53423));
    Span4Mux_h I__12994 (
            .O(N__53513),
            .I(N__53423));
    Span4Mux_h I__12993 (
            .O(N__53510),
            .I(N__53423));
    Span4Mux_v I__12992 (
            .O(N__53507),
            .I(N__53420));
    LocalMux I__12991 (
            .O(N__53502),
            .I(N__53409));
    LocalMux I__12990 (
            .O(N__53499),
            .I(N__53409));
    LocalMux I__12989 (
            .O(N__53496),
            .I(N__53409));
    Span12Mux_v I__12988 (
            .O(N__53493),
            .I(N__53409));
    Span12Mux_v I__12987 (
            .O(N__53490),
            .I(N__53409));
    InMux I__12986 (
            .O(N__53489),
            .I(N__53406));
    Span4Mux_v I__12985 (
            .O(N__53486),
            .I(N__53397));
    Span4Mux_h I__12984 (
            .O(N__53483),
            .I(N__53397));
    Span4Mux_h I__12983 (
            .O(N__53480),
            .I(N__53397));
    Span4Mux_h I__12982 (
            .O(N__53475),
            .I(N__53397));
    Span4Mux_h I__12981 (
            .O(N__53472),
            .I(N__53388));
    Span4Mux_h I__12980 (
            .O(N__53469),
            .I(N__53388));
    Span4Mux_v I__12979 (
            .O(N__53466),
            .I(N__53388));
    Span4Mux_h I__12978 (
            .O(N__53459),
            .I(N__53388));
    InMux I__12977 (
            .O(N__53458),
            .I(N__53383));
    InMux I__12976 (
            .O(N__53457),
            .I(N__53383));
    LocalMux I__12975 (
            .O(N__53454),
            .I(comm_cmd_2));
    LocalMux I__12974 (
            .O(N__53447),
            .I(comm_cmd_2));
    Odrv4 I__12973 (
            .O(N__53444),
            .I(comm_cmd_2));
    LocalMux I__12972 (
            .O(N__53441),
            .I(comm_cmd_2));
    Odrv4 I__12971 (
            .O(N__53430),
            .I(comm_cmd_2));
    Odrv4 I__12970 (
            .O(N__53423),
            .I(comm_cmd_2));
    Odrv4 I__12969 (
            .O(N__53420),
            .I(comm_cmd_2));
    Odrv12 I__12968 (
            .O(N__53409),
            .I(comm_cmd_2));
    LocalMux I__12967 (
            .O(N__53406),
            .I(comm_cmd_2));
    Odrv4 I__12966 (
            .O(N__53397),
            .I(comm_cmd_2));
    Odrv4 I__12965 (
            .O(N__53388),
            .I(comm_cmd_2));
    LocalMux I__12964 (
            .O(N__53383),
            .I(comm_cmd_2));
    InMux I__12963 (
            .O(N__53358),
            .I(N__53355));
    LocalMux I__12962 (
            .O(N__53355),
            .I(n22402));
    InMux I__12961 (
            .O(N__53352),
            .I(N__53348));
    InMux I__12960 (
            .O(N__53351),
            .I(N__53345));
    LocalMux I__12959 (
            .O(N__53348),
            .I(N__53342));
    LocalMux I__12958 (
            .O(N__53345),
            .I(N__53339));
    Odrv4 I__12957 (
            .O(N__53342),
            .I(\ADC_VDC.genclk.n21444 ));
    Odrv4 I__12956 (
            .O(N__53339),
            .I(\ADC_VDC.genclk.n21444 ));
    SRMux I__12955 (
            .O(N__53334),
            .I(N__53331));
    LocalMux I__12954 (
            .O(N__53331),
            .I(N__53328));
    Odrv12 I__12953 (
            .O(N__53328),
            .I(\comm_spi.DOUT_7__N_747 ));
    ClkMux I__12952 (
            .O(N__53325),
            .I(N__53321));
    IoInMux I__12951 (
            .O(N__53324),
            .I(N__53315));
    LocalMux I__12950 (
            .O(N__53321),
            .I(N__53312));
    ClkMux I__12949 (
            .O(N__53320),
            .I(N__53309));
    ClkMux I__12948 (
            .O(N__53319),
            .I(N__53306));
    ClkMux I__12947 (
            .O(N__53318),
            .I(N__53303));
    LocalMux I__12946 (
            .O(N__53315),
            .I(N__53295));
    Span4Mux_v I__12945 (
            .O(N__53312),
            .I(N__53288));
    LocalMux I__12944 (
            .O(N__53309),
            .I(N__53288));
    LocalMux I__12943 (
            .O(N__53306),
            .I(N__53285));
    LocalMux I__12942 (
            .O(N__53303),
            .I(N__53282));
    ClkMux I__12941 (
            .O(N__53302),
            .I(N__53279));
    ClkMux I__12940 (
            .O(N__53301),
            .I(N__53272));
    ClkMux I__12939 (
            .O(N__53300),
            .I(N__53269));
    ClkMux I__12938 (
            .O(N__53299),
            .I(N__53266));
    ClkMux I__12937 (
            .O(N__53298),
            .I(N__53262));
    Span4Mux_s3_h I__12936 (
            .O(N__53295),
            .I(N__53257));
    ClkMux I__12935 (
            .O(N__53294),
            .I(N__53250));
    ClkMux I__12934 (
            .O(N__53293),
            .I(N__53247));
    Span4Mux_v I__12933 (
            .O(N__53288),
            .I(N__53244));
    Span4Mux_h I__12932 (
            .O(N__53285),
            .I(N__53237));
    Span4Mux_v I__12931 (
            .O(N__53282),
            .I(N__53237));
    LocalMux I__12930 (
            .O(N__53279),
            .I(N__53237));
    ClkMux I__12929 (
            .O(N__53278),
            .I(N__53234));
    ClkMux I__12928 (
            .O(N__53277),
            .I(N__53231));
    ClkMux I__12927 (
            .O(N__53276),
            .I(N__53228));
    ClkMux I__12926 (
            .O(N__53275),
            .I(N__53225));
    LocalMux I__12925 (
            .O(N__53272),
            .I(N__53220));
    LocalMux I__12924 (
            .O(N__53269),
            .I(N__53220));
    LocalMux I__12923 (
            .O(N__53266),
            .I(N__53217));
    ClkMux I__12922 (
            .O(N__53265),
            .I(N__53214));
    LocalMux I__12921 (
            .O(N__53262),
            .I(N__53211));
    ClkMux I__12920 (
            .O(N__53261),
            .I(N__53208));
    ClkMux I__12919 (
            .O(N__53260),
            .I(N__53204));
    Span4Mux_h I__12918 (
            .O(N__53257),
            .I(N__53201));
    ClkMux I__12917 (
            .O(N__53256),
            .I(N__53198));
    ClkMux I__12916 (
            .O(N__53255),
            .I(N__53195));
    ClkMux I__12915 (
            .O(N__53254),
            .I(N__53191));
    ClkMux I__12914 (
            .O(N__53253),
            .I(N__53188));
    LocalMux I__12913 (
            .O(N__53250),
            .I(N__53183));
    LocalMux I__12912 (
            .O(N__53247),
            .I(N__53183));
    Span4Mux_v I__12911 (
            .O(N__53244),
            .I(N__53176));
    Span4Mux_v I__12910 (
            .O(N__53237),
            .I(N__53176));
    LocalMux I__12909 (
            .O(N__53234),
            .I(N__53176));
    LocalMux I__12908 (
            .O(N__53231),
            .I(N__53173));
    LocalMux I__12907 (
            .O(N__53228),
            .I(N__53168));
    LocalMux I__12906 (
            .O(N__53225),
            .I(N__53168));
    Span4Mux_v I__12905 (
            .O(N__53220),
            .I(N__53163));
    Span4Mux_v I__12904 (
            .O(N__53217),
            .I(N__53163));
    LocalMux I__12903 (
            .O(N__53214),
            .I(N__53160));
    Span4Mux_v I__12902 (
            .O(N__53211),
            .I(N__53155));
    LocalMux I__12901 (
            .O(N__53208),
            .I(N__53155));
    ClkMux I__12900 (
            .O(N__53207),
            .I(N__53152));
    LocalMux I__12899 (
            .O(N__53204),
            .I(N__53149));
    Span4Mux_h I__12898 (
            .O(N__53201),
            .I(N__53142));
    LocalMux I__12897 (
            .O(N__53198),
            .I(N__53142));
    LocalMux I__12896 (
            .O(N__53195),
            .I(N__53142));
    ClkMux I__12895 (
            .O(N__53194),
            .I(N__53139));
    LocalMux I__12894 (
            .O(N__53191),
            .I(N__53132));
    LocalMux I__12893 (
            .O(N__53188),
            .I(N__53132));
    Span4Mux_v I__12892 (
            .O(N__53183),
            .I(N__53132));
    Span4Mux_h I__12891 (
            .O(N__53176),
            .I(N__53129));
    Span4Mux_h I__12890 (
            .O(N__53173),
            .I(N__53124));
    Span4Mux_v I__12889 (
            .O(N__53168),
            .I(N__53124));
    Span4Mux_h I__12888 (
            .O(N__53163),
            .I(N__53119));
    Span4Mux_v I__12887 (
            .O(N__53160),
            .I(N__53119));
    Span4Mux_h I__12886 (
            .O(N__53155),
            .I(N__53114));
    LocalMux I__12885 (
            .O(N__53152),
            .I(N__53114));
    Span4Mux_h I__12884 (
            .O(N__53149),
            .I(N__53109));
    Span4Mux_h I__12883 (
            .O(N__53142),
            .I(N__53109));
    LocalMux I__12882 (
            .O(N__53139),
            .I(N__53106));
    Sp12to4 I__12881 (
            .O(N__53132),
            .I(N__53103));
    Span4Mux_h I__12880 (
            .O(N__53129),
            .I(N__53100));
    Span4Mux_h I__12879 (
            .O(N__53124),
            .I(N__53093));
    Span4Mux_v I__12878 (
            .O(N__53119),
            .I(N__53093));
    Span4Mux_v I__12877 (
            .O(N__53114),
            .I(N__53093));
    Span4Mux_h I__12876 (
            .O(N__53109),
            .I(N__53088));
    Span4Mux_v I__12875 (
            .O(N__53106),
            .I(N__53088));
    Span12Mux_h I__12874 (
            .O(N__53103),
            .I(N__53085));
    Span4Mux_h I__12873 (
            .O(N__53100),
            .I(N__53082));
    Sp12to4 I__12872 (
            .O(N__53093),
            .I(N__53079));
    Span4Mux_h I__12871 (
            .O(N__53088),
            .I(N__53076));
    Odrv12 I__12870 (
            .O(N__53085),
            .I(VDC_CLK));
    Odrv4 I__12869 (
            .O(N__53082),
            .I(VDC_CLK));
    Odrv12 I__12868 (
            .O(N__53079),
            .I(VDC_CLK));
    Odrv4 I__12867 (
            .O(N__53076),
            .I(VDC_CLK));
    InMux I__12866 (
            .O(N__53067),
            .I(N__53064));
    LocalMux I__12865 (
            .O(N__53064),
            .I(\comm_spi.n14614 ));
    InMux I__12864 (
            .O(N__53061),
            .I(N__53058));
    LocalMux I__12863 (
            .O(N__53058),
            .I(\comm_spi.n14615 ));
    InMux I__12862 (
            .O(N__53055),
            .I(N__53052));
    LocalMux I__12861 (
            .O(N__53052),
            .I(N__53047));
    InMux I__12860 (
            .O(N__53051),
            .I(N__53044));
    InMux I__12859 (
            .O(N__53050),
            .I(N__53041));
    Span4Mux_v I__12858 (
            .O(N__53047),
            .I(N__53030));
    LocalMux I__12857 (
            .O(N__53044),
            .I(N__53030));
    LocalMux I__12856 (
            .O(N__53041),
            .I(N__53027));
    InMux I__12855 (
            .O(N__53040),
            .I(N__53022));
    InMux I__12854 (
            .O(N__53039),
            .I(N__53022));
    InMux I__12853 (
            .O(N__53038),
            .I(N__53019));
    InMux I__12852 (
            .O(N__53037),
            .I(N__53016));
    InMux I__12851 (
            .O(N__53036),
            .I(N__53013));
    InMux I__12850 (
            .O(N__53035),
            .I(N__53010));
    Span4Mux_v I__12849 (
            .O(N__53030),
            .I(N__53007));
    Sp12to4 I__12848 (
            .O(N__53027),
            .I(N__53000));
    LocalMux I__12847 (
            .O(N__53022),
            .I(N__53000));
    LocalMux I__12846 (
            .O(N__53019),
            .I(N__53000));
    LocalMux I__12845 (
            .O(N__53016),
            .I(N__52995));
    LocalMux I__12844 (
            .O(N__53013),
            .I(N__52995));
    LocalMux I__12843 (
            .O(N__53010),
            .I(N__52992));
    Span4Mux_h I__12842 (
            .O(N__53007),
            .I(N__52989));
    Span12Mux_v I__12841 (
            .O(N__53000),
            .I(N__52986));
    Span4Mux_h I__12840 (
            .O(N__52995),
            .I(N__52983));
    Span4Mux_v I__12839 (
            .O(N__52992),
            .I(N__52980));
    Odrv4 I__12838 (
            .O(N__52989),
            .I(comm_rx_buf_0));
    Odrv12 I__12837 (
            .O(N__52986),
            .I(comm_rx_buf_0));
    Odrv4 I__12836 (
            .O(N__52983),
            .I(comm_rx_buf_0));
    Odrv4 I__12835 (
            .O(N__52980),
            .I(comm_rx_buf_0));
    InMux I__12834 (
            .O(N__52971),
            .I(N__52966));
    InMux I__12833 (
            .O(N__52970),
            .I(N__52963));
    InMux I__12832 (
            .O(N__52969),
            .I(N__52960));
    LocalMux I__12831 (
            .O(N__52966),
            .I(\comm_spi.n22866 ));
    LocalMux I__12830 (
            .O(N__52963),
            .I(\comm_spi.n22866 ));
    LocalMux I__12829 (
            .O(N__52960),
            .I(\comm_spi.n22866 ));
    CascadeMux I__12828 (
            .O(N__52953),
            .I(\comm_spi.n22866_cascade_ ));
    InMux I__12827 (
            .O(N__52950),
            .I(N__52945));
    InMux I__12826 (
            .O(N__52949),
            .I(N__52942));
    InMux I__12825 (
            .O(N__52948),
            .I(N__52939));
    LocalMux I__12824 (
            .O(N__52945),
            .I(N__52934));
    LocalMux I__12823 (
            .O(N__52942),
            .I(N__52934));
    LocalMux I__12822 (
            .O(N__52939),
            .I(N__52931));
    Span4Mux_v I__12821 (
            .O(N__52934),
            .I(N__52928));
    Odrv4 I__12820 (
            .O(N__52931),
            .I(\comm_spi.n14601 ));
    Odrv4 I__12819 (
            .O(N__52928),
            .I(\comm_spi.n14601 ));
    CascadeMux I__12818 (
            .O(N__52923),
            .I(\comm_spi.imosi_cascade_ ));
    SRMux I__12817 (
            .O(N__52920),
            .I(N__52917));
    LocalMux I__12816 (
            .O(N__52917),
            .I(N__52914));
    Span4Mux_v I__12815 (
            .O(N__52914),
            .I(N__52911));
    Odrv4 I__12814 (
            .O(N__52911),
            .I(\comm_spi.DOUT_7__N_746 ));
    InMux I__12813 (
            .O(N__52908),
            .I(N__52901));
    InMux I__12812 (
            .O(N__52907),
            .I(N__52901));
    InMux I__12811 (
            .O(N__52906),
            .I(N__52898));
    LocalMux I__12810 (
            .O(N__52901),
            .I(N__52895));
    LocalMux I__12809 (
            .O(N__52898),
            .I(N__52890));
    Span4Mux_h I__12808 (
            .O(N__52895),
            .I(N__52887));
    InMux I__12807 (
            .O(N__52894),
            .I(N__52882));
    InMux I__12806 (
            .O(N__52893),
            .I(N__52882));
    Odrv12 I__12805 (
            .O(N__52890),
            .I(\ADC_VDC.genclk.div_state_0 ));
    Odrv4 I__12804 (
            .O(N__52887),
            .I(\ADC_VDC.genclk.div_state_0 ));
    LocalMux I__12803 (
            .O(N__52882),
            .I(\ADC_VDC.genclk.div_state_0 ));
    InMux I__12802 (
            .O(N__52875),
            .I(N__52871));
    InMux I__12801 (
            .O(N__52874),
            .I(N__52868));
    LocalMux I__12800 (
            .O(N__52871),
            .I(\comm_spi.imosi ));
    LocalMux I__12799 (
            .O(N__52868),
            .I(\comm_spi.imosi ));
    InMux I__12798 (
            .O(N__52863),
            .I(N__52859));
    InMux I__12797 (
            .O(N__52862),
            .I(N__52856));
    LocalMux I__12796 (
            .O(N__52859),
            .I(\comm_spi.n22863 ));
    LocalMux I__12795 (
            .O(N__52856),
            .I(\comm_spi.n22863 ));
    InMux I__12794 (
            .O(N__52851),
            .I(N__52848));
    LocalMux I__12793 (
            .O(N__52848),
            .I(N__52845));
    Span4Mux_h I__12792 (
            .O(N__52845),
            .I(N__52841));
    InMux I__12791 (
            .O(N__52844),
            .I(N__52837));
    Span4Mux_h I__12790 (
            .O(N__52841),
            .I(N__52834));
    InMux I__12789 (
            .O(N__52840),
            .I(N__52831));
    LocalMux I__12788 (
            .O(N__52837),
            .I(req_data_cnt_5));
    Odrv4 I__12787 (
            .O(N__52834),
            .I(req_data_cnt_5));
    LocalMux I__12786 (
            .O(N__52831),
            .I(req_data_cnt_5));
    CascadeMux I__12785 (
            .O(N__52824),
            .I(n22345_cascade_));
    InMux I__12784 (
            .O(N__52821),
            .I(N__52818));
    LocalMux I__12783 (
            .O(N__52818),
            .I(N__52815));
    Span4Mux_h I__12782 (
            .O(N__52815),
            .I(N__52812));
    Span4Mux_h I__12781 (
            .O(N__52812),
            .I(N__52807));
    InMux I__12780 (
            .O(N__52811),
            .I(N__52802));
    InMux I__12779 (
            .O(N__52810),
            .I(N__52802));
    Odrv4 I__12778 (
            .O(N__52807),
            .I(acadc_skipCount_5));
    LocalMux I__12777 (
            .O(N__52802),
            .I(acadc_skipCount_5));
    CascadeMux I__12776 (
            .O(N__52797),
            .I(n22348_cascade_));
    InMux I__12775 (
            .O(N__52794),
            .I(N__52791));
    LocalMux I__12774 (
            .O(N__52791),
            .I(n30_adj_1500));
    InMux I__12773 (
            .O(N__52788),
            .I(N__52784));
    InMux I__12772 (
            .O(N__52787),
            .I(N__52781));
    LocalMux I__12771 (
            .O(N__52784),
            .I(N__52778));
    LocalMux I__12770 (
            .O(N__52781),
            .I(N__52775));
    Span4Mux_v I__12769 (
            .O(N__52778),
            .I(N__52771));
    Span4Mux_h I__12768 (
            .O(N__52775),
            .I(N__52768));
    InMux I__12767 (
            .O(N__52774),
            .I(N__52765));
    Sp12to4 I__12766 (
            .O(N__52771),
            .I(N__52762));
    Span4Mux_h I__12765 (
            .O(N__52768),
            .I(N__52759));
    LocalMux I__12764 (
            .O(N__52765),
            .I(buf_adcdata_iac_11));
    Odrv12 I__12763 (
            .O(N__52762),
            .I(buf_adcdata_iac_11));
    Odrv4 I__12762 (
            .O(N__52759),
            .I(buf_adcdata_iac_11));
    InMux I__12761 (
            .O(N__52752),
            .I(N__52749));
    LocalMux I__12760 (
            .O(N__52749),
            .I(n16_adj_1514));
    InMux I__12759 (
            .O(N__52746),
            .I(N__52743));
    LocalMux I__12758 (
            .O(N__52743),
            .I(N__52740));
    Span4Mux_h I__12757 (
            .O(N__52740),
            .I(N__52737));
    Odrv4 I__12756 (
            .O(N__52737),
            .I(n21126));
    InMux I__12755 (
            .O(N__52734),
            .I(N__52731));
    LocalMux I__12754 (
            .O(N__52731),
            .I(N__52728));
    Span4Mux_h I__12753 (
            .O(N__52728),
            .I(N__52725));
    Odrv4 I__12752 (
            .O(N__52725),
            .I(buf_data_iac_10));
    CascadeMux I__12751 (
            .O(N__52722),
            .I(N__52719));
    InMux I__12750 (
            .O(N__52719),
            .I(N__52716));
    LocalMux I__12749 (
            .O(N__52716),
            .I(N__52713));
    Span4Mux_v I__12748 (
            .O(N__52713),
            .I(N__52710));
    Odrv4 I__12747 (
            .O(N__52710),
            .I(n21564));
    InMux I__12746 (
            .O(N__52707),
            .I(N__52704));
    LocalMux I__12745 (
            .O(N__52704),
            .I(N__52701));
    Span4Mux_v I__12744 (
            .O(N__52701),
            .I(N__52698));
    Odrv4 I__12743 (
            .O(N__52698),
            .I(buf_data_iac_8));
    InMux I__12742 (
            .O(N__52695),
            .I(N__52692));
    LocalMux I__12741 (
            .O(N__52692),
            .I(N__52689));
    Span4Mux_h I__12740 (
            .O(N__52689),
            .I(N__52686));
    Span4Mux_v I__12739 (
            .O(N__52686),
            .I(N__52683));
    Odrv4 I__12738 (
            .O(N__52683),
            .I(n21218));
    InMux I__12737 (
            .O(N__52680),
            .I(N__52677));
    LocalMux I__12736 (
            .O(N__52677),
            .I(N__52674));
    Odrv4 I__12735 (
            .O(N__52674),
            .I(buf_data_iac_23));
    CascadeMux I__12734 (
            .O(N__52671),
            .I(N__52668));
    InMux I__12733 (
            .O(N__52668),
            .I(N__52665));
    LocalMux I__12732 (
            .O(N__52665),
            .I(N__52662));
    Span12Mux_h I__12731 (
            .O(N__52662),
            .I(N__52659));
    Span12Mux_h I__12730 (
            .O(N__52659),
            .I(N__52656));
    Span12Mux_v I__12729 (
            .O(N__52656),
            .I(N__52653));
    Odrv12 I__12728 (
            .O(N__52653),
            .I(n21364));
    CEMux I__12727 (
            .O(N__52650),
            .I(N__52647));
    LocalMux I__12726 (
            .O(N__52647),
            .I(N__52644));
    Odrv12 I__12725 (
            .O(N__52644),
            .I(\ADC_VDC.genclk.n6 ));
    ClkMux I__12724 (
            .O(N__52641),
            .I(N__52635));
    ClkMux I__12723 (
            .O(N__52640),
            .I(N__52632));
    ClkMux I__12722 (
            .O(N__52639),
            .I(N__52629));
    ClkMux I__12721 (
            .O(N__52638),
            .I(N__52623));
    LocalMux I__12720 (
            .O(N__52635),
            .I(N__52620));
    LocalMux I__12719 (
            .O(N__52632),
            .I(N__52617));
    LocalMux I__12718 (
            .O(N__52629),
            .I(N__52614));
    ClkMux I__12717 (
            .O(N__52628),
            .I(N__52611));
    ClkMux I__12716 (
            .O(N__52627),
            .I(N__52606));
    ClkMux I__12715 (
            .O(N__52626),
            .I(N__52603));
    LocalMux I__12714 (
            .O(N__52623),
            .I(N__52598));
    Span4Mux_v I__12713 (
            .O(N__52620),
            .I(N__52589));
    Span4Mux_h I__12712 (
            .O(N__52617),
            .I(N__52589));
    Span4Mux_v I__12711 (
            .O(N__52614),
            .I(N__52589));
    LocalMux I__12710 (
            .O(N__52611),
            .I(N__52589));
    ClkMux I__12709 (
            .O(N__52610),
            .I(N__52583));
    ClkMux I__12708 (
            .O(N__52609),
            .I(N__52580));
    LocalMux I__12707 (
            .O(N__52606),
            .I(N__52577));
    LocalMux I__12706 (
            .O(N__52603),
            .I(N__52574));
    ClkMux I__12705 (
            .O(N__52602),
            .I(N__52571));
    ClkMux I__12704 (
            .O(N__52601),
            .I(N__52567));
    Span4Mux_v I__12703 (
            .O(N__52598),
            .I(N__52562));
    Span4Mux_v I__12702 (
            .O(N__52589),
            .I(N__52562));
    ClkMux I__12701 (
            .O(N__52588),
            .I(N__52559));
    ClkMux I__12700 (
            .O(N__52587),
            .I(N__52556));
    ClkMux I__12699 (
            .O(N__52586),
            .I(N__52553));
    LocalMux I__12698 (
            .O(N__52583),
            .I(N__52549));
    LocalMux I__12697 (
            .O(N__52580),
            .I(N__52543));
    Span4Mux_h I__12696 (
            .O(N__52577),
            .I(N__52538));
    Span4Mux_v I__12695 (
            .O(N__52574),
            .I(N__52538));
    LocalMux I__12694 (
            .O(N__52571),
            .I(N__52535));
    ClkMux I__12693 (
            .O(N__52570),
            .I(N__52532));
    LocalMux I__12692 (
            .O(N__52567),
            .I(N__52528));
    Span4Mux_h I__12691 (
            .O(N__52562),
            .I(N__52523));
    LocalMux I__12690 (
            .O(N__52559),
            .I(N__52523));
    LocalMux I__12689 (
            .O(N__52556),
            .I(N__52518));
    LocalMux I__12688 (
            .O(N__52553),
            .I(N__52518));
    ClkMux I__12687 (
            .O(N__52552),
            .I(N__52515));
    Span4Mux_h I__12686 (
            .O(N__52549),
            .I(N__52512));
    ClkMux I__12685 (
            .O(N__52548),
            .I(N__52509));
    ClkMux I__12684 (
            .O(N__52547),
            .I(N__52506));
    ClkMux I__12683 (
            .O(N__52546),
            .I(N__52503));
    Span4Mux_h I__12682 (
            .O(N__52543),
            .I(N__52499));
    Span4Mux_h I__12681 (
            .O(N__52538),
            .I(N__52495));
    Span4Mux_v I__12680 (
            .O(N__52535),
            .I(N__52490));
    LocalMux I__12679 (
            .O(N__52532),
            .I(N__52490));
    ClkMux I__12678 (
            .O(N__52531),
            .I(N__52487));
    Span4Mux_h I__12677 (
            .O(N__52528),
            .I(N__52482));
    Span4Mux_h I__12676 (
            .O(N__52523),
            .I(N__52482));
    Span4Mux_v I__12675 (
            .O(N__52518),
            .I(N__52473));
    LocalMux I__12674 (
            .O(N__52515),
            .I(N__52473));
    Span4Mux_v I__12673 (
            .O(N__52512),
            .I(N__52473));
    LocalMux I__12672 (
            .O(N__52509),
            .I(N__52473));
    LocalMux I__12671 (
            .O(N__52506),
            .I(N__52468));
    LocalMux I__12670 (
            .O(N__52503),
            .I(N__52468));
    ClkMux I__12669 (
            .O(N__52502),
            .I(N__52465));
    Span4Mux_h I__12668 (
            .O(N__52499),
            .I(N__52462));
    ClkMux I__12667 (
            .O(N__52498),
            .I(N__52459));
    Sp12to4 I__12666 (
            .O(N__52495),
            .I(N__52452));
    Sp12to4 I__12665 (
            .O(N__52490),
            .I(N__52452));
    LocalMux I__12664 (
            .O(N__52487),
            .I(N__52452));
    Span4Mux_v I__12663 (
            .O(N__52482),
            .I(N__52449));
    Span4Mux_h I__12662 (
            .O(N__52473),
            .I(N__52442));
    Span4Mux_v I__12661 (
            .O(N__52468),
            .I(N__52442));
    LocalMux I__12660 (
            .O(N__52465),
            .I(N__52442));
    Span4Mux_v I__12659 (
            .O(N__52462),
            .I(N__52437));
    LocalMux I__12658 (
            .O(N__52459),
            .I(N__52437));
    Odrv12 I__12657 (
            .O(N__52452),
            .I(\comm_spi.iclk ));
    Odrv4 I__12656 (
            .O(N__52449),
            .I(\comm_spi.iclk ));
    Odrv4 I__12655 (
            .O(N__52442),
            .I(\comm_spi.iclk ));
    Odrv4 I__12654 (
            .O(N__52437),
            .I(\comm_spi.iclk ));
    InMux I__12653 (
            .O(N__52428),
            .I(N__52425));
    LocalMux I__12652 (
            .O(N__52425),
            .I(N__52422));
    Span4Mux_h I__12651 (
            .O(N__52422),
            .I(N__52419));
    Odrv4 I__12650 (
            .O(N__52419),
            .I(n4_adj_1600));
    CascadeMux I__12649 (
            .O(N__52416),
            .I(n4_adj_1600_cascade_));
    InMux I__12648 (
            .O(N__52413),
            .I(N__52401));
    InMux I__12647 (
            .O(N__52412),
            .I(N__52398));
    InMux I__12646 (
            .O(N__52411),
            .I(N__52395));
    InMux I__12645 (
            .O(N__52410),
            .I(N__52392));
    InMux I__12644 (
            .O(N__52409),
            .I(N__52389));
    InMux I__12643 (
            .O(N__52408),
            .I(N__52383));
    InMux I__12642 (
            .O(N__52407),
            .I(N__52374));
    InMux I__12641 (
            .O(N__52406),
            .I(N__52374));
    InMux I__12640 (
            .O(N__52405),
            .I(N__52374));
    InMux I__12639 (
            .O(N__52404),
            .I(N__52374));
    LocalMux I__12638 (
            .O(N__52401),
            .I(N__52371));
    LocalMux I__12637 (
            .O(N__52398),
            .I(N__52367));
    LocalMux I__12636 (
            .O(N__52395),
            .I(N__52362));
    LocalMux I__12635 (
            .O(N__52392),
            .I(N__52362));
    LocalMux I__12634 (
            .O(N__52389),
            .I(N__52359));
    InMux I__12633 (
            .O(N__52388),
            .I(N__52356));
    InMux I__12632 (
            .O(N__52387),
            .I(N__52351));
    InMux I__12631 (
            .O(N__52386),
            .I(N__52348));
    LocalMux I__12630 (
            .O(N__52383),
            .I(N__52339));
    LocalMux I__12629 (
            .O(N__52374),
            .I(N__52339));
    Span4Mux_v I__12628 (
            .O(N__52371),
            .I(N__52336));
    InMux I__12627 (
            .O(N__52370),
            .I(N__52333));
    Span4Mux_v I__12626 (
            .O(N__52367),
            .I(N__52321));
    Span4Mux_v I__12625 (
            .O(N__52362),
            .I(N__52321));
    Span4Mux_h I__12624 (
            .O(N__52359),
            .I(N__52321));
    LocalMux I__12623 (
            .O(N__52356),
            .I(N__52321));
    InMux I__12622 (
            .O(N__52355),
            .I(N__52316));
    InMux I__12621 (
            .O(N__52354),
            .I(N__52316));
    LocalMux I__12620 (
            .O(N__52351),
            .I(N__52311));
    LocalMux I__12619 (
            .O(N__52348),
            .I(N__52311));
    InMux I__12618 (
            .O(N__52347),
            .I(N__52302));
    InMux I__12617 (
            .O(N__52346),
            .I(N__52302));
    InMux I__12616 (
            .O(N__52345),
            .I(N__52302));
    InMux I__12615 (
            .O(N__52344),
            .I(N__52302));
    Span4Mux_h I__12614 (
            .O(N__52339),
            .I(N__52299));
    Span4Mux_v I__12613 (
            .O(N__52336),
            .I(N__52294));
    LocalMux I__12612 (
            .O(N__52333),
            .I(N__52294));
    InMux I__12611 (
            .O(N__52332),
            .I(N__52287));
    InMux I__12610 (
            .O(N__52331),
            .I(N__52287));
    InMux I__12609 (
            .O(N__52330),
            .I(N__52287));
    Span4Mux_h I__12608 (
            .O(N__52321),
            .I(N__52284));
    LocalMux I__12607 (
            .O(N__52316),
            .I(comm_index_1));
    Odrv4 I__12606 (
            .O(N__52311),
            .I(comm_index_1));
    LocalMux I__12605 (
            .O(N__52302),
            .I(comm_index_1));
    Odrv4 I__12604 (
            .O(N__52299),
            .I(comm_index_1));
    Odrv4 I__12603 (
            .O(N__52294),
            .I(comm_index_1));
    LocalMux I__12602 (
            .O(N__52287),
            .I(comm_index_1));
    Odrv4 I__12601 (
            .O(N__52284),
            .I(comm_index_1));
    CascadeMux I__12600 (
            .O(N__52269),
            .I(n5_cascade_));
    InMux I__12599 (
            .O(N__52266),
            .I(N__52262));
    InMux I__12598 (
            .O(N__52265),
            .I(N__52259));
    LocalMux I__12597 (
            .O(N__52262),
            .I(N__52255));
    LocalMux I__12596 (
            .O(N__52259),
            .I(N__52251));
    InMux I__12595 (
            .O(N__52258),
            .I(N__52248));
    Span4Mux_h I__12594 (
            .O(N__52255),
            .I(N__52245));
    InMux I__12593 (
            .O(N__52254),
            .I(N__52240));
    Span4Mux_h I__12592 (
            .O(N__52251),
            .I(N__52237));
    LocalMux I__12591 (
            .O(N__52248),
            .I(N__52234));
    Span4Mux_h I__12590 (
            .O(N__52245),
            .I(N__52231));
    InMux I__12589 (
            .O(N__52244),
            .I(N__52228));
    InMux I__12588 (
            .O(N__52243),
            .I(N__52225));
    LocalMux I__12587 (
            .O(N__52240),
            .I(comm_cmd_7));
    Odrv4 I__12586 (
            .O(N__52237),
            .I(comm_cmd_7));
    Odrv4 I__12585 (
            .O(N__52234),
            .I(comm_cmd_7));
    Odrv4 I__12584 (
            .O(N__52231),
            .I(comm_cmd_7));
    LocalMux I__12583 (
            .O(N__52228),
            .I(comm_cmd_7));
    LocalMux I__12582 (
            .O(N__52225),
            .I(comm_cmd_7));
    InMux I__12581 (
            .O(N__52212),
            .I(N__52209));
    LocalMux I__12580 (
            .O(N__52209),
            .I(N__52206));
    Span4Mux_h I__12579 (
            .O(N__52206),
            .I(N__52203));
    Span4Mux_h I__12578 (
            .O(N__52203),
            .I(N__52200));
    Odrv4 I__12577 (
            .O(N__52200),
            .I(n21888));
    CascadeMux I__12576 (
            .O(N__52197),
            .I(N__52194));
    InMux I__12575 (
            .O(N__52194),
            .I(N__52191));
    LocalMux I__12574 (
            .O(N__52191),
            .I(n21317));
    InMux I__12573 (
            .O(N__52188),
            .I(N__52184));
    InMux I__12572 (
            .O(N__52187),
            .I(N__52181));
    LocalMux I__12571 (
            .O(N__52184),
            .I(N__52178));
    LocalMux I__12570 (
            .O(N__52181),
            .I(N__52174));
    Span4Mux_v I__12569 (
            .O(N__52178),
            .I(N__52171));
    CascadeMux I__12568 (
            .O(N__52177),
            .I(N__52168));
    Span12Mux_v I__12567 (
            .O(N__52174),
            .I(N__52165));
    Sp12to4 I__12566 (
            .O(N__52171),
            .I(N__52162));
    InMux I__12565 (
            .O(N__52168),
            .I(N__52159));
    Span12Mux_h I__12564 (
            .O(N__52165),
            .I(N__52156));
    Span12Mux_h I__12563 (
            .O(N__52162),
            .I(N__52153));
    LocalMux I__12562 (
            .O(N__52159),
            .I(buf_adcdata_iac_15));
    Odrv12 I__12561 (
            .O(N__52156),
            .I(buf_adcdata_iac_15));
    Odrv12 I__12560 (
            .O(N__52153),
            .I(buf_adcdata_iac_15));
    InMux I__12559 (
            .O(N__52146),
            .I(N__52143));
    LocalMux I__12558 (
            .O(N__52143),
            .I(N__52140));
    Sp12to4 I__12557 (
            .O(N__52140),
            .I(N__52137));
    Odrv12 I__12556 (
            .O(N__52137),
            .I(n16_adj_1504));
    InMux I__12555 (
            .O(N__52134),
            .I(N__52131));
    LocalMux I__12554 (
            .O(N__52131),
            .I(N__52128));
    Odrv4 I__12553 (
            .O(N__52128),
            .I(n21048));
    CascadeMux I__12552 (
            .O(N__52125),
            .I(N__52121));
    InMux I__12551 (
            .O(N__52124),
            .I(N__52118));
    InMux I__12550 (
            .O(N__52121),
            .I(N__52114));
    LocalMux I__12549 (
            .O(N__52118),
            .I(N__52108));
    InMux I__12548 (
            .O(N__52117),
            .I(N__52105));
    LocalMux I__12547 (
            .O(N__52114),
            .I(N__52102));
    InMux I__12546 (
            .O(N__52113),
            .I(N__52099));
    InMux I__12545 (
            .O(N__52112),
            .I(N__52096));
    InMux I__12544 (
            .O(N__52111),
            .I(N__52093));
    Span4Mux_h I__12543 (
            .O(N__52108),
            .I(N__52087));
    LocalMux I__12542 (
            .O(N__52105),
            .I(N__52087));
    Span4Mux_h I__12541 (
            .O(N__52102),
            .I(N__52084));
    LocalMux I__12540 (
            .O(N__52099),
            .I(N__52079));
    LocalMux I__12539 (
            .O(N__52096),
            .I(N__52079));
    LocalMux I__12538 (
            .O(N__52093),
            .I(N__52076));
    InMux I__12537 (
            .O(N__52092),
            .I(N__52073));
    Sp12to4 I__12536 (
            .O(N__52087),
            .I(N__52066));
    Sp12to4 I__12535 (
            .O(N__52084),
            .I(N__52066));
    Sp12to4 I__12534 (
            .O(N__52079),
            .I(N__52066));
    Span4Mux_v I__12533 (
            .O(N__52076),
            .I(N__52063));
    LocalMux I__12532 (
            .O(N__52073),
            .I(N__52060));
    Span12Mux_v I__12531 (
            .O(N__52066),
            .I(N__52055));
    Span4Mux_h I__12530 (
            .O(N__52063),
            .I(N__52052));
    Span4Mux_v I__12529 (
            .O(N__52060),
            .I(N__52049));
    InMux I__12528 (
            .O(N__52059),
            .I(N__52046));
    InMux I__12527 (
            .O(N__52058),
            .I(N__52043));
    Odrv12 I__12526 (
            .O(N__52055),
            .I(comm_rx_buf_5));
    Odrv4 I__12525 (
            .O(N__52052),
            .I(comm_rx_buf_5));
    Odrv4 I__12524 (
            .O(N__52049),
            .I(comm_rx_buf_5));
    LocalMux I__12523 (
            .O(N__52046),
            .I(comm_rx_buf_5));
    LocalMux I__12522 (
            .O(N__52043),
            .I(comm_rx_buf_5));
    InMux I__12521 (
            .O(N__52032),
            .I(N__52029));
    LocalMux I__12520 (
            .O(N__52029),
            .I(N__52023));
    InMux I__12519 (
            .O(N__52028),
            .I(N__52004));
    InMux I__12518 (
            .O(N__52027),
            .I(N__52001));
    InMux I__12517 (
            .O(N__52026),
            .I(N__51989));
    Span4Mux_v I__12516 (
            .O(N__52023),
            .I(N__51986));
    InMux I__12515 (
            .O(N__52022),
            .I(N__51983));
    InMux I__12514 (
            .O(N__52021),
            .I(N__51978));
    InMux I__12513 (
            .O(N__52020),
            .I(N__51978));
    InMux I__12512 (
            .O(N__52019),
            .I(N__51961));
    InMux I__12511 (
            .O(N__52018),
            .I(N__51961));
    InMux I__12510 (
            .O(N__52017),
            .I(N__51961));
    InMux I__12509 (
            .O(N__52016),
            .I(N__51961));
    InMux I__12508 (
            .O(N__52015),
            .I(N__51961));
    InMux I__12507 (
            .O(N__52014),
            .I(N__51961));
    InMux I__12506 (
            .O(N__52013),
            .I(N__51961));
    InMux I__12505 (
            .O(N__52012),
            .I(N__51961));
    InMux I__12504 (
            .O(N__52011),
            .I(N__51951));
    InMux I__12503 (
            .O(N__52010),
            .I(N__51951));
    InMux I__12502 (
            .O(N__52009),
            .I(N__51951));
    InMux I__12501 (
            .O(N__52008),
            .I(N__51940));
    InMux I__12500 (
            .O(N__52007),
            .I(N__51937));
    LocalMux I__12499 (
            .O(N__52004),
            .I(N__51932));
    LocalMux I__12498 (
            .O(N__52001),
            .I(N__51932));
    InMux I__12497 (
            .O(N__52000),
            .I(N__51929));
    InMux I__12496 (
            .O(N__51999),
            .I(N__51926));
    InMux I__12495 (
            .O(N__51998),
            .I(N__51921));
    InMux I__12494 (
            .O(N__51997),
            .I(N__51918));
    CascadeMux I__12493 (
            .O(N__51996),
            .I(N__51913));
    CascadeMux I__12492 (
            .O(N__51995),
            .I(N__51910));
    InMux I__12491 (
            .O(N__51994),
            .I(N__51906));
    InMux I__12490 (
            .O(N__51993),
            .I(N__51901));
    InMux I__12489 (
            .O(N__51992),
            .I(N__51898));
    LocalMux I__12488 (
            .O(N__51989),
            .I(N__51887));
    Span4Mux_h I__12487 (
            .O(N__51986),
            .I(N__51887));
    LocalMux I__12486 (
            .O(N__51983),
            .I(N__51887));
    LocalMux I__12485 (
            .O(N__51978),
            .I(N__51887));
    LocalMux I__12484 (
            .O(N__51961),
            .I(N__51887));
    InMux I__12483 (
            .O(N__51960),
            .I(N__51884));
    InMux I__12482 (
            .O(N__51959),
            .I(N__51881));
    CascadeMux I__12481 (
            .O(N__51958),
            .I(N__51873));
    LocalMux I__12480 (
            .O(N__51951),
            .I(N__51855));
    InMux I__12479 (
            .O(N__51950),
            .I(N__51838));
    InMux I__12478 (
            .O(N__51949),
            .I(N__51838));
    InMux I__12477 (
            .O(N__51948),
            .I(N__51838));
    InMux I__12476 (
            .O(N__51947),
            .I(N__51838));
    InMux I__12475 (
            .O(N__51946),
            .I(N__51838));
    InMux I__12474 (
            .O(N__51945),
            .I(N__51838));
    InMux I__12473 (
            .O(N__51944),
            .I(N__51838));
    InMux I__12472 (
            .O(N__51943),
            .I(N__51838));
    LocalMux I__12471 (
            .O(N__51940),
            .I(N__51827));
    LocalMux I__12470 (
            .O(N__51937),
            .I(N__51827));
    Span4Mux_v I__12469 (
            .O(N__51932),
            .I(N__51827));
    LocalMux I__12468 (
            .O(N__51929),
            .I(N__51827));
    LocalMux I__12467 (
            .O(N__51926),
            .I(N__51827));
    InMux I__12466 (
            .O(N__51925),
            .I(N__51821));
    InMux I__12465 (
            .O(N__51924),
            .I(N__51818));
    LocalMux I__12464 (
            .O(N__51921),
            .I(N__51813));
    LocalMux I__12463 (
            .O(N__51918),
            .I(N__51813));
    InMux I__12462 (
            .O(N__51917),
            .I(N__51808));
    InMux I__12461 (
            .O(N__51916),
            .I(N__51808));
    InMux I__12460 (
            .O(N__51913),
            .I(N__51801));
    InMux I__12459 (
            .O(N__51910),
            .I(N__51801));
    InMux I__12458 (
            .O(N__51909),
            .I(N__51801));
    LocalMux I__12457 (
            .O(N__51906),
            .I(N__51796));
    InMux I__12456 (
            .O(N__51905),
            .I(N__51793));
    InMux I__12455 (
            .O(N__51904),
            .I(N__51789));
    LocalMux I__12454 (
            .O(N__51901),
            .I(N__51778));
    LocalMux I__12453 (
            .O(N__51898),
            .I(N__51778));
    Span4Mux_v I__12452 (
            .O(N__51887),
            .I(N__51778));
    LocalMux I__12451 (
            .O(N__51884),
            .I(N__51778));
    LocalMux I__12450 (
            .O(N__51881),
            .I(N__51778));
    InMux I__12449 (
            .O(N__51880),
            .I(N__51775));
    InMux I__12448 (
            .O(N__51879),
            .I(N__51772));
    InMux I__12447 (
            .O(N__51878),
            .I(N__51769));
    InMux I__12446 (
            .O(N__51877),
            .I(N__51762));
    InMux I__12445 (
            .O(N__51876),
            .I(N__51762));
    InMux I__12444 (
            .O(N__51873),
            .I(N__51762));
    InMux I__12443 (
            .O(N__51872),
            .I(N__51755));
    InMux I__12442 (
            .O(N__51871),
            .I(N__51740));
    InMux I__12441 (
            .O(N__51870),
            .I(N__51740));
    InMux I__12440 (
            .O(N__51869),
            .I(N__51740));
    InMux I__12439 (
            .O(N__51868),
            .I(N__51740));
    InMux I__12438 (
            .O(N__51867),
            .I(N__51740));
    InMux I__12437 (
            .O(N__51866),
            .I(N__51740));
    InMux I__12436 (
            .O(N__51865),
            .I(N__51740));
    InMux I__12435 (
            .O(N__51864),
            .I(N__51731));
    InMux I__12434 (
            .O(N__51863),
            .I(N__51731));
    InMux I__12433 (
            .O(N__51862),
            .I(N__51731));
    InMux I__12432 (
            .O(N__51861),
            .I(N__51731));
    InMux I__12431 (
            .O(N__51860),
            .I(N__51728));
    CascadeMux I__12430 (
            .O(N__51859),
            .I(N__51715));
    InMux I__12429 (
            .O(N__51858),
            .I(N__51711));
    Span4Mux_v I__12428 (
            .O(N__51855),
            .I(N__51708));
    LocalMux I__12427 (
            .O(N__51838),
            .I(N__51703));
    Span4Mux_v I__12426 (
            .O(N__51827),
            .I(N__51703));
    InMux I__12425 (
            .O(N__51826),
            .I(N__51696));
    InMux I__12424 (
            .O(N__51825),
            .I(N__51696));
    InMux I__12423 (
            .O(N__51824),
            .I(N__51696));
    LocalMux I__12422 (
            .O(N__51821),
            .I(N__51685));
    LocalMux I__12421 (
            .O(N__51818),
            .I(N__51685));
    Span4Mux_v I__12420 (
            .O(N__51813),
            .I(N__51685));
    LocalMux I__12419 (
            .O(N__51808),
            .I(N__51685));
    LocalMux I__12418 (
            .O(N__51801),
            .I(N__51685));
    InMux I__12417 (
            .O(N__51800),
            .I(N__51682));
    InMux I__12416 (
            .O(N__51799),
            .I(N__51679));
    Span4Mux_v I__12415 (
            .O(N__51796),
            .I(N__51674));
    LocalMux I__12414 (
            .O(N__51793),
            .I(N__51674));
    InMux I__12413 (
            .O(N__51792),
            .I(N__51671));
    LocalMux I__12412 (
            .O(N__51789),
            .I(N__51666));
    Span4Mux_v I__12411 (
            .O(N__51778),
            .I(N__51666));
    LocalMux I__12410 (
            .O(N__51775),
            .I(N__51657));
    LocalMux I__12409 (
            .O(N__51772),
            .I(N__51657));
    LocalMux I__12408 (
            .O(N__51769),
            .I(N__51657));
    LocalMux I__12407 (
            .O(N__51762),
            .I(N__51657));
    InMux I__12406 (
            .O(N__51761),
            .I(N__51646));
    CascadeMux I__12405 (
            .O(N__51760),
            .I(N__51638));
    CascadeMux I__12404 (
            .O(N__51759),
            .I(N__51633));
    InMux I__12403 (
            .O(N__51758),
            .I(N__51629));
    LocalMux I__12402 (
            .O(N__51755),
            .I(N__51626));
    LocalMux I__12401 (
            .O(N__51740),
            .I(N__51623));
    LocalMux I__12400 (
            .O(N__51731),
            .I(N__51620));
    LocalMux I__12399 (
            .O(N__51728),
            .I(N__51617));
    InMux I__12398 (
            .O(N__51727),
            .I(N__51614));
    InMux I__12397 (
            .O(N__51726),
            .I(N__51611));
    InMux I__12396 (
            .O(N__51725),
            .I(N__51604));
    InMux I__12395 (
            .O(N__51724),
            .I(N__51604));
    InMux I__12394 (
            .O(N__51723),
            .I(N__51604));
    InMux I__12393 (
            .O(N__51722),
            .I(N__51599));
    InMux I__12392 (
            .O(N__51721),
            .I(N__51599));
    InMux I__12391 (
            .O(N__51720),
            .I(N__51596));
    InMux I__12390 (
            .O(N__51719),
            .I(N__51587));
    InMux I__12389 (
            .O(N__51718),
            .I(N__51587));
    InMux I__12388 (
            .O(N__51715),
            .I(N__51587));
    InMux I__12387 (
            .O(N__51714),
            .I(N__51587));
    LocalMux I__12386 (
            .O(N__51711),
            .I(N__51578));
    Span4Mux_h I__12385 (
            .O(N__51708),
            .I(N__51578));
    Span4Mux_h I__12384 (
            .O(N__51703),
            .I(N__51578));
    LocalMux I__12383 (
            .O(N__51696),
            .I(N__51578));
    Span4Mux_v I__12382 (
            .O(N__51685),
            .I(N__51575));
    LocalMux I__12381 (
            .O(N__51682),
            .I(N__51569));
    LocalMux I__12380 (
            .O(N__51679),
            .I(N__51566));
    Span4Mux_v I__12379 (
            .O(N__51674),
            .I(N__51563));
    LocalMux I__12378 (
            .O(N__51671),
            .I(N__51556));
    Span4Mux_h I__12377 (
            .O(N__51666),
            .I(N__51556));
    Span4Mux_v I__12376 (
            .O(N__51657),
            .I(N__51556));
    InMux I__12375 (
            .O(N__51656),
            .I(N__51539));
    InMux I__12374 (
            .O(N__51655),
            .I(N__51539));
    InMux I__12373 (
            .O(N__51654),
            .I(N__51539));
    InMux I__12372 (
            .O(N__51653),
            .I(N__51539));
    InMux I__12371 (
            .O(N__51652),
            .I(N__51539));
    InMux I__12370 (
            .O(N__51651),
            .I(N__51539));
    InMux I__12369 (
            .O(N__51650),
            .I(N__51539));
    InMux I__12368 (
            .O(N__51649),
            .I(N__51539));
    LocalMux I__12367 (
            .O(N__51646),
            .I(N__51536));
    InMux I__12366 (
            .O(N__51645),
            .I(N__51533));
    InMux I__12365 (
            .O(N__51644),
            .I(N__51526));
    InMux I__12364 (
            .O(N__51643),
            .I(N__51526));
    InMux I__12363 (
            .O(N__51642),
            .I(N__51526));
    InMux I__12362 (
            .O(N__51641),
            .I(N__51519));
    InMux I__12361 (
            .O(N__51638),
            .I(N__51519));
    InMux I__12360 (
            .O(N__51637),
            .I(N__51519));
    InMux I__12359 (
            .O(N__51636),
            .I(N__51512));
    InMux I__12358 (
            .O(N__51633),
            .I(N__51512));
    InMux I__12357 (
            .O(N__51632),
            .I(N__51512));
    LocalMux I__12356 (
            .O(N__51629),
            .I(N__51503));
    Span4Mux_h I__12355 (
            .O(N__51626),
            .I(N__51503));
    Span4Mux_h I__12354 (
            .O(N__51623),
            .I(N__51503));
    Span4Mux_v I__12353 (
            .O(N__51620),
            .I(N__51503));
    Span12Mux_v I__12352 (
            .O(N__51617),
            .I(N__51496));
    LocalMux I__12351 (
            .O(N__51614),
            .I(N__51496));
    LocalMux I__12350 (
            .O(N__51611),
            .I(N__51496));
    LocalMux I__12349 (
            .O(N__51604),
            .I(N__51491));
    LocalMux I__12348 (
            .O(N__51599),
            .I(N__51491));
    LocalMux I__12347 (
            .O(N__51596),
            .I(N__51486));
    LocalMux I__12346 (
            .O(N__51587),
            .I(N__51486));
    Span4Mux_v I__12345 (
            .O(N__51578),
            .I(N__51481));
    Span4Mux_h I__12344 (
            .O(N__51575),
            .I(N__51481));
    InMux I__12343 (
            .O(N__51574),
            .I(N__51474));
    InMux I__12342 (
            .O(N__51573),
            .I(N__51474));
    InMux I__12341 (
            .O(N__51572),
            .I(N__51474));
    Span4Mux_v I__12340 (
            .O(N__51569),
            .I(N__51465));
    Span4Mux_v I__12339 (
            .O(N__51566),
            .I(N__51465));
    Span4Mux_h I__12338 (
            .O(N__51563),
            .I(N__51465));
    Span4Mux_v I__12337 (
            .O(N__51556),
            .I(N__51465));
    LocalMux I__12336 (
            .O(N__51539),
            .I(comm_state_1));
    Odrv4 I__12335 (
            .O(N__51536),
            .I(comm_state_1));
    LocalMux I__12334 (
            .O(N__51533),
            .I(comm_state_1));
    LocalMux I__12333 (
            .O(N__51526),
            .I(comm_state_1));
    LocalMux I__12332 (
            .O(N__51519),
            .I(comm_state_1));
    LocalMux I__12331 (
            .O(N__51512),
            .I(comm_state_1));
    Odrv4 I__12330 (
            .O(N__51503),
            .I(comm_state_1));
    Odrv12 I__12329 (
            .O(N__51496),
            .I(comm_state_1));
    Odrv12 I__12328 (
            .O(N__51491),
            .I(comm_state_1));
    Odrv4 I__12327 (
            .O(N__51486),
            .I(comm_state_1));
    Odrv4 I__12326 (
            .O(N__51481),
            .I(comm_state_1));
    LocalMux I__12325 (
            .O(N__51474),
            .I(comm_state_1));
    Odrv4 I__12324 (
            .O(N__51465),
            .I(comm_state_1));
    InMux I__12323 (
            .O(N__51438),
            .I(N__51432));
    InMux I__12322 (
            .O(N__51437),
            .I(N__51429));
    InMux I__12321 (
            .O(N__51436),
            .I(N__51425));
    InMux I__12320 (
            .O(N__51435),
            .I(N__51422));
    LocalMux I__12319 (
            .O(N__51432),
            .I(N__51419));
    LocalMux I__12318 (
            .O(N__51429),
            .I(N__51416));
    InMux I__12317 (
            .O(N__51428),
            .I(N__51413));
    LocalMux I__12316 (
            .O(N__51425),
            .I(N__51410));
    LocalMux I__12315 (
            .O(N__51422),
            .I(N__51407));
    Span4Mux_v I__12314 (
            .O(N__51419),
            .I(N__51400));
    Span4Mux_h I__12313 (
            .O(N__51416),
            .I(N__51400));
    LocalMux I__12312 (
            .O(N__51413),
            .I(N__51400));
    Span4Mux_v I__12311 (
            .O(N__51410),
            .I(N__51397));
    Span12Mux_v I__12310 (
            .O(N__51407),
            .I(N__51394));
    Span4Mux_h I__12309 (
            .O(N__51400),
            .I(N__51389));
    Span4Mux_v I__12308 (
            .O(N__51397),
            .I(N__51389));
    Odrv12 I__12307 (
            .O(N__51394),
            .I(comm_buf_1_5));
    Odrv4 I__12306 (
            .O(N__51389),
            .I(comm_buf_1_5));
    CEMux I__12305 (
            .O(N__51384),
            .I(N__51378));
    CEMux I__12304 (
            .O(N__51383),
            .I(N__51375));
    CEMux I__12303 (
            .O(N__51382),
            .I(N__51371));
    CEMux I__12302 (
            .O(N__51381),
            .I(N__51368));
    LocalMux I__12301 (
            .O(N__51378),
            .I(N__51365));
    LocalMux I__12300 (
            .O(N__51375),
            .I(N__51362));
    CEMux I__12299 (
            .O(N__51374),
            .I(N__51359));
    LocalMux I__12298 (
            .O(N__51371),
            .I(N__51353));
    LocalMux I__12297 (
            .O(N__51368),
            .I(N__51350));
    Span4Mux_h I__12296 (
            .O(N__51365),
            .I(N__51347));
    Span4Mux_h I__12295 (
            .O(N__51362),
            .I(N__51342));
    LocalMux I__12294 (
            .O(N__51359),
            .I(N__51342));
    CEMux I__12293 (
            .O(N__51358),
            .I(N__51339));
    CEMux I__12292 (
            .O(N__51357),
            .I(N__51336));
    CEMux I__12291 (
            .O(N__51356),
            .I(N__51333));
    Span4Mux_h I__12290 (
            .O(N__51353),
            .I(N__51330));
    Span4Mux_v I__12289 (
            .O(N__51350),
            .I(N__51327));
    Sp12to4 I__12288 (
            .O(N__51347),
            .I(N__51324));
    Span4Mux_v I__12287 (
            .O(N__51342),
            .I(N__51321));
    LocalMux I__12286 (
            .O(N__51339),
            .I(n11991));
    LocalMux I__12285 (
            .O(N__51336),
            .I(n11991));
    LocalMux I__12284 (
            .O(N__51333),
            .I(n11991));
    Odrv4 I__12283 (
            .O(N__51330),
            .I(n11991));
    Odrv4 I__12282 (
            .O(N__51327),
            .I(n11991));
    Odrv12 I__12281 (
            .O(N__51324),
            .I(n11991));
    Odrv4 I__12280 (
            .O(N__51321),
            .I(n11991));
    SRMux I__12279 (
            .O(N__51306),
            .I(N__51303));
    LocalMux I__12278 (
            .O(N__51303),
            .I(N__51296));
    SRMux I__12277 (
            .O(N__51302),
            .I(N__51293));
    SRMux I__12276 (
            .O(N__51301),
            .I(N__51290));
    SRMux I__12275 (
            .O(N__51300),
            .I(N__51287));
    SRMux I__12274 (
            .O(N__51299),
            .I(N__51284));
    Span4Mux_h I__12273 (
            .O(N__51296),
            .I(N__51278));
    LocalMux I__12272 (
            .O(N__51293),
            .I(N__51278));
    LocalMux I__12271 (
            .O(N__51290),
            .I(N__51270));
    LocalMux I__12270 (
            .O(N__51287),
            .I(N__51270));
    LocalMux I__12269 (
            .O(N__51284),
            .I(N__51270));
    SRMux I__12268 (
            .O(N__51283),
            .I(N__51267));
    Span4Mux_h I__12267 (
            .O(N__51278),
            .I(N__51264));
    SRMux I__12266 (
            .O(N__51277),
            .I(N__51261));
    Span4Mux_v I__12265 (
            .O(N__51270),
            .I(N__51258));
    LocalMux I__12264 (
            .O(N__51267),
            .I(N__51250));
    Span4Mux_h I__12263 (
            .O(N__51264),
            .I(N__51250));
    LocalMux I__12262 (
            .O(N__51261),
            .I(N__51250));
    Span4Mux_h I__12261 (
            .O(N__51258),
            .I(N__51247));
    SRMux I__12260 (
            .O(N__51257),
            .I(N__51244));
    Span4Mux_v I__12259 (
            .O(N__51250),
            .I(N__51241));
    Sp12to4 I__12258 (
            .O(N__51247),
            .I(N__51238));
    LocalMux I__12257 (
            .O(N__51244),
            .I(N__51233));
    Sp12to4 I__12256 (
            .O(N__51241),
            .I(N__51233));
    Odrv12 I__12255 (
            .O(N__51238),
            .I(n14757));
    Odrv12 I__12254 (
            .O(N__51233),
            .I(n14757));
    InMux I__12253 (
            .O(N__51228),
            .I(N__51225));
    LocalMux I__12252 (
            .O(N__51225),
            .I(N__51222));
    Span4Mux_v I__12251 (
            .O(N__51222),
            .I(N__51219));
    Span4Mux_h I__12250 (
            .O(N__51219),
            .I(N__51216));
    Span4Mux_h I__12249 (
            .O(N__51216),
            .I(N__51213));
    Odrv4 I__12248 (
            .O(N__51213),
            .I(n19_adj_1497));
    CascadeMux I__12247 (
            .O(N__51210),
            .I(N__51207));
    InMux I__12246 (
            .O(N__51207),
            .I(N__51204));
    LocalMux I__12245 (
            .O(N__51204),
            .I(N__51201));
    Span4Mux_v I__12244 (
            .O(N__51201),
            .I(N__51198));
    Span4Mux_h I__12243 (
            .O(N__51198),
            .I(N__51195));
    Span4Mux_h I__12242 (
            .O(N__51195),
            .I(N__51191));
    CascadeMux I__12241 (
            .O(N__51194),
            .I(N__51188));
    Span4Mux_h I__12240 (
            .O(N__51191),
            .I(N__51185));
    InMux I__12239 (
            .O(N__51188),
            .I(N__51182));
    Odrv4 I__12238 (
            .O(N__51185),
            .I(buf_readRTD_5));
    LocalMux I__12237 (
            .O(N__51182),
            .I(buf_readRTD_5));
    InMux I__12236 (
            .O(N__51177),
            .I(N__51173));
    CascadeMux I__12235 (
            .O(N__51176),
            .I(N__51170));
    LocalMux I__12234 (
            .O(N__51173),
            .I(N__51167));
    InMux I__12233 (
            .O(N__51170),
            .I(N__51164));
    Span4Mux_h I__12232 (
            .O(N__51167),
            .I(N__51161));
    LocalMux I__12231 (
            .O(N__51164),
            .I(data_idxvec_5));
    Odrv4 I__12230 (
            .O(N__51161),
            .I(data_idxvec_5));
    InMux I__12229 (
            .O(N__51156),
            .I(N__51152));
    InMux I__12228 (
            .O(N__51155),
            .I(N__51148));
    LocalMux I__12227 (
            .O(N__51152),
            .I(N__51145));
    InMux I__12226 (
            .O(N__51151),
            .I(N__51142));
    LocalMux I__12225 (
            .O(N__51148),
            .I(N__51139));
    Span4Mux_h I__12224 (
            .O(N__51145),
            .I(N__51136));
    LocalMux I__12223 (
            .O(N__51142),
            .I(data_cntvec_5));
    Odrv4 I__12222 (
            .O(N__51139),
            .I(data_cntvec_5));
    Odrv4 I__12221 (
            .O(N__51136),
            .I(data_cntvec_5));
    CascadeMux I__12220 (
            .O(N__51129),
            .I(n26_adj_1498_cascade_));
    CascadeMux I__12219 (
            .O(N__51126),
            .I(n21132_cascade_));
    InMux I__12218 (
            .O(N__51123),
            .I(N__51120));
    LocalMux I__12217 (
            .O(N__51120),
            .I(n21127));
    CascadeMux I__12216 (
            .O(N__51117),
            .I(n22333_cascade_));
    InMux I__12215 (
            .O(N__51114),
            .I(N__51111));
    LocalMux I__12214 (
            .O(N__51111),
            .I(N__51103));
    InMux I__12213 (
            .O(N__51110),
            .I(N__51100));
    InMux I__12212 (
            .O(N__51109),
            .I(N__51097));
    InMux I__12211 (
            .O(N__51108),
            .I(N__51094));
    InMux I__12210 (
            .O(N__51107),
            .I(N__51091));
    CascadeMux I__12209 (
            .O(N__51106),
            .I(N__51088));
    Span4Mux_v I__12208 (
            .O(N__51103),
            .I(N__51083));
    LocalMux I__12207 (
            .O(N__51100),
            .I(N__51083));
    LocalMux I__12206 (
            .O(N__51097),
            .I(N__51078));
    LocalMux I__12205 (
            .O(N__51094),
            .I(N__51078));
    LocalMux I__12204 (
            .O(N__51091),
            .I(N__51075));
    InMux I__12203 (
            .O(N__51088),
            .I(N__51072));
    Span4Mux_v I__12202 (
            .O(N__51083),
            .I(N__51068));
    Span4Mux_v I__12201 (
            .O(N__51078),
            .I(N__51065));
    Span4Mux_v I__12200 (
            .O(N__51075),
            .I(N__51062));
    LocalMux I__12199 (
            .O(N__51072),
            .I(N__51059));
    InMux I__12198 (
            .O(N__51071),
            .I(N__51056));
    Sp12to4 I__12197 (
            .O(N__51068),
            .I(N__51049));
    Sp12to4 I__12196 (
            .O(N__51065),
            .I(N__51049));
    Span4Mux_h I__12195 (
            .O(N__51062),
            .I(N__51046));
    Span4Mux_v I__12194 (
            .O(N__51059),
            .I(N__51041));
    LocalMux I__12193 (
            .O(N__51056),
            .I(N__51041));
    InMux I__12192 (
            .O(N__51055),
            .I(N__51038));
    InMux I__12191 (
            .O(N__51054),
            .I(N__51035));
    Odrv12 I__12190 (
            .O(N__51049),
            .I(comm_rx_buf_3));
    Odrv4 I__12189 (
            .O(N__51046),
            .I(comm_rx_buf_3));
    Odrv4 I__12188 (
            .O(N__51041),
            .I(comm_rx_buf_3));
    LocalMux I__12187 (
            .O(N__51038),
            .I(comm_rx_buf_3));
    LocalMux I__12186 (
            .O(N__51035),
            .I(comm_rx_buf_3));
    CascadeMux I__12185 (
            .O(N__51024),
            .I(n22336_cascade_));
    CascadeMux I__12184 (
            .O(N__51021),
            .I(N__51016));
    CascadeMux I__12183 (
            .O(N__51020),
            .I(N__51013));
    InMux I__12182 (
            .O(N__51019),
            .I(N__51009));
    InMux I__12181 (
            .O(N__51016),
            .I(N__51006));
    InMux I__12180 (
            .O(N__51013),
            .I(N__51003));
    InMux I__12179 (
            .O(N__51012),
            .I(N__51000));
    LocalMux I__12178 (
            .O(N__51009),
            .I(N__50996));
    LocalMux I__12177 (
            .O(N__51006),
            .I(N__50993));
    LocalMux I__12176 (
            .O(N__51003),
            .I(N__50990));
    LocalMux I__12175 (
            .O(N__51000),
            .I(N__50987));
    InMux I__12174 (
            .O(N__50999),
            .I(N__50984));
    Span4Mux_v I__12173 (
            .O(N__50996),
            .I(N__50981));
    Span4Mux_v I__12172 (
            .O(N__50993),
            .I(N__50978));
    Span4Mux_v I__12171 (
            .O(N__50990),
            .I(N__50973));
    Span4Mux_v I__12170 (
            .O(N__50987),
            .I(N__50973));
    LocalMux I__12169 (
            .O(N__50984),
            .I(N__50970));
    Span4Mux_v I__12168 (
            .O(N__50981),
            .I(N__50967));
    Span4Mux_v I__12167 (
            .O(N__50978),
            .I(N__50962));
    Span4Mux_h I__12166 (
            .O(N__50973),
            .I(N__50962));
    Sp12to4 I__12165 (
            .O(N__50970),
            .I(N__50959));
    Span4Mux_h I__12164 (
            .O(N__50967),
            .I(N__50956));
    Odrv4 I__12163 (
            .O(N__50962),
            .I(comm_buf_1_3));
    Odrv12 I__12162 (
            .O(N__50959),
            .I(comm_buf_1_3));
    Odrv4 I__12161 (
            .O(N__50956),
            .I(comm_buf_1_3));
    InMux I__12160 (
            .O(N__50949),
            .I(N__50946));
    LocalMux I__12159 (
            .O(N__50946),
            .I(N__50943));
    Span4Mux_v I__12158 (
            .O(N__50943),
            .I(N__50940));
    Span4Mux_h I__12157 (
            .O(N__50940),
            .I(N__50936));
    CascadeMux I__12156 (
            .O(N__50939),
            .I(N__50933));
    Span4Mux_h I__12155 (
            .O(N__50936),
            .I(N__50930));
    InMux I__12154 (
            .O(N__50933),
            .I(N__50927));
    Odrv4 I__12153 (
            .O(N__50930),
            .I(buf_adcdata_vdc_11));
    LocalMux I__12152 (
            .O(N__50927),
            .I(buf_adcdata_vdc_11));
    InMux I__12151 (
            .O(N__50922),
            .I(N__50917));
    InMux I__12150 (
            .O(N__50921),
            .I(N__50914));
    CascadeMux I__12149 (
            .O(N__50920),
            .I(N__50911));
    LocalMux I__12148 (
            .O(N__50917),
            .I(N__50908));
    LocalMux I__12147 (
            .O(N__50914),
            .I(N__50905));
    InMux I__12146 (
            .O(N__50911),
            .I(N__50902));
    Span12Mux_v I__12145 (
            .O(N__50908),
            .I(N__50899));
    Span12Mux_h I__12144 (
            .O(N__50905),
            .I(N__50896));
    LocalMux I__12143 (
            .O(N__50902),
            .I(buf_adcdata_vac_11));
    Odrv12 I__12142 (
            .O(N__50899),
            .I(buf_adcdata_vac_11));
    Odrv12 I__12141 (
            .O(N__50896),
            .I(buf_adcdata_vac_11));
    InMux I__12140 (
            .O(N__50889),
            .I(N__50886));
    LocalMux I__12139 (
            .O(N__50886),
            .I(n19_adj_1515));
    InMux I__12138 (
            .O(N__50883),
            .I(N__50879));
    CascadeMux I__12137 (
            .O(N__50882),
            .I(N__50876));
    LocalMux I__12136 (
            .O(N__50879),
            .I(N__50873));
    InMux I__12135 (
            .O(N__50876),
            .I(N__50870));
    Span4Mux_v I__12134 (
            .O(N__50873),
            .I(N__50867));
    LocalMux I__12133 (
            .O(N__50870),
            .I(data_idxvec_3));
    Odrv4 I__12132 (
            .O(N__50867),
            .I(data_idxvec_3));
    InMux I__12131 (
            .O(N__50862),
            .I(N__50858));
    InMux I__12130 (
            .O(N__50861),
            .I(N__50855));
    LocalMux I__12129 (
            .O(N__50858),
            .I(N__50851));
    LocalMux I__12128 (
            .O(N__50855),
            .I(N__50848));
    InMux I__12127 (
            .O(N__50854),
            .I(N__50845));
    Span4Mux_h I__12126 (
            .O(N__50851),
            .I(N__50840));
    Span4Mux_h I__12125 (
            .O(N__50848),
            .I(N__50840));
    LocalMux I__12124 (
            .O(N__50845),
            .I(data_cntvec_3));
    Odrv4 I__12123 (
            .O(N__50840),
            .I(data_cntvec_3));
    InMux I__12122 (
            .O(N__50835),
            .I(N__50832));
    LocalMux I__12121 (
            .O(N__50832),
            .I(N__50829));
    Span4Mux_h I__12120 (
            .O(N__50829),
            .I(N__50826));
    Span4Mux_v I__12119 (
            .O(N__50826),
            .I(N__50823));
    Odrv4 I__12118 (
            .O(N__50823),
            .I(buf_data_iac_11));
    CascadeMux I__12117 (
            .O(N__50820),
            .I(n26_adj_1516_cascade_));
    InMux I__12116 (
            .O(N__50817),
            .I(N__50814));
    LocalMux I__12115 (
            .O(N__50814),
            .I(n21133));
    CascadeMux I__12114 (
            .O(N__50811),
            .I(n21316_cascade_));
    InMux I__12113 (
            .O(N__50808),
            .I(N__50802));
    InMux I__12112 (
            .O(N__50807),
            .I(N__50802));
    LocalMux I__12111 (
            .O(N__50802),
            .I(comm_length_2));
    CascadeMux I__12110 (
            .O(N__50799),
            .I(N__50787));
    CascadeMux I__12109 (
            .O(N__50798),
            .I(N__50783));
    InMux I__12108 (
            .O(N__50797),
            .I(N__50768));
    InMux I__12107 (
            .O(N__50796),
            .I(N__50768));
    InMux I__12106 (
            .O(N__50795),
            .I(N__50768));
    InMux I__12105 (
            .O(N__50794),
            .I(N__50768));
    InMux I__12104 (
            .O(N__50793),
            .I(N__50761));
    InMux I__12103 (
            .O(N__50792),
            .I(N__50761));
    InMux I__12102 (
            .O(N__50791),
            .I(N__50761));
    InMux I__12101 (
            .O(N__50790),
            .I(N__50758));
    InMux I__12100 (
            .O(N__50787),
            .I(N__50748));
    InMux I__12099 (
            .O(N__50786),
            .I(N__50743));
    InMux I__12098 (
            .O(N__50783),
            .I(N__50743));
    InMux I__12097 (
            .O(N__50782),
            .I(N__50740));
    CascadeMux I__12096 (
            .O(N__50781),
            .I(N__50737));
    CascadeMux I__12095 (
            .O(N__50780),
            .I(N__50734));
    InMux I__12094 (
            .O(N__50779),
            .I(N__50726));
    InMux I__12093 (
            .O(N__50778),
            .I(N__50721));
    InMux I__12092 (
            .O(N__50777),
            .I(N__50721));
    LocalMux I__12091 (
            .O(N__50768),
            .I(N__50714));
    LocalMux I__12090 (
            .O(N__50761),
            .I(N__50714));
    LocalMux I__12089 (
            .O(N__50758),
            .I(N__50714));
    InMux I__12088 (
            .O(N__50757),
            .I(N__50705));
    InMux I__12087 (
            .O(N__50756),
            .I(N__50705));
    InMux I__12086 (
            .O(N__50755),
            .I(N__50705));
    InMux I__12085 (
            .O(N__50754),
            .I(N__50705));
    InMux I__12084 (
            .O(N__50753),
            .I(N__50702));
    InMux I__12083 (
            .O(N__50752),
            .I(N__50697));
    InMux I__12082 (
            .O(N__50751),
            .I(N__50697));
    LocalMux I__12081 (
            .O(N__50748),
            .I(N__50694));
    LocalMux I__12080 (
            .O(N__50743),
            .I(N__50689));
    LocalMux I__12079 (
            .O(N__50740),
            .I(N__50689));
    InMux I__12078 (
            .O(N__50737),
            .I(N__50681));
    InMux I__12077 (
            .O(N__50734),
            .I(N__50681));
    InMux I__12076 (
            .O(N__50733),
            .I(N__50681));
    InMux I__12075 (
            .O(N__50732),
            .I(N__50672));
    InMux I__12074 (
            .O(N__50731),
            .I(N__50672));
    InMux I__12073 (
            .O(N__50730),
            .I(N__50672));
    InMux I__12072 (
            .O(N__50729),
            .I(N__50672));
    LocalMux I__12071 (
            .O(N__50726),
            .I(N__50659));
    LocalMux I__12070 (
            .O(N__50721),
            .I(N__50659));
    Span4Mux_v I__12069 (
            .O(N__50714),
            .I(N__50659));
    LocalMux I__12068 (
            .O(N__50705),
            .I(N__50659));
    LocalMux I__12067 (
            .O(N__50702),
            .I(N__50654));
    LocalMux I__12066 (
            .O(N__50697),
            .I(N__50647));
    Span4Mux_h I__12065 (
            .O(N__50694),
            .I(N__50647));
    Span4Mux_v I__12064 (
            .O(N__50689),
            .I(N__50647));
    InMux I__12063 (
            .O(N__50688),
            .I(N__50644));
    LocalMux I__12062 (
            .O(N__50681),
            .I(N__50639));
    LocalMux I__12061 (
            .O(N__50672),
            .I(N__50639));
    InMux I__12060 (
            .O(N__50671),
            .I(N__50630));
    InMux I__12059 (
            .O(N__50670),
            .I(N__50630));
    InMux I__12058 (
            .O(N__50669),
            .I(N__50630));
    InMux I__12057 (
            .O(N__50668),
            .I(N__50630));
    Span4Mux_h I__12056 (
            .O(N__50659),
            .I(N__50627));
    InMux I__12055 (
            .O(N__50658),
            .I(N__50622));
    InMux I__12054 (
            .O(N__50657),
            .I(N__50622));
    Span4Mux_h I__12053 (
            .O(N__50654),
            .I(N__50617));
    Span4Mux_h I__12052 (
            .O(N__50647),
            .I(N__50617));
    LocalMux I__12051 (
            .O(N__50644),
            .I(comm_index_0));
    Odrv4 I__12050 (
            .O(N__50639),
            .I(comm_index_0));
    LocalMux I__12049 (
            .O(N__50630),
            .I(comm_index_0));
    Odrv4 I__12048 (
            .O(N__50627),
            .I(comm_index_0));
    LocalMux I__12047 (
            .O(N__50622),
            .I(comm_index_0));
    Odrv4 I__12046 (
            .O(N__50617),
            .I(comm_index_0));
    InMux I__12045 (
            .O(N__50604),
            .I(N__50588));
    InMux I__12044 (
            .O(N__50603),
            .I(N__50588));
    InMux I__12043 (
            .O(N__50602),
            .I(N__50585));
    InMux I__12042 (
            .O(N__50601),
            .I(N__50581));
    InMux I__12041 (
            .O(N__50600),
            .I(N__50573));
    InMux I__12040 (
            .O(N__50599),
            .I(N__50573));
    InMux I__12039 (
            .O(N__50598),
            .I(N__50566));
    InMux I__12038 (
            .O(N__50597),
            .I(N__50566));
    InMux I__12037 (
            .O(N__50596),
            .I(N__50557));
    InMux I__12036 (
            .O(N__50595),
            .I(N__50557));
    InMux I__12035 (
            .O(N__50594),
            .I(N__50557));
    InMux I__12034 (
            .O(N__50593),
            .I(N__50557));
    LocalMux I__12033 (
            .O(N__50588),
            .I(N__50552));
    LocalMux I__12032 (
            .O(N__50585),
            .I(N__50552));
    InMux I__12031 (
            .O(N__50584),
            .I(N__50549));
    LocalMux I__12030 (
            .O(N__50581),
            .I(N__50546));
    InMux I__12029 (
            .O(N__50580),
            .I(N__50543));
    InMux I__12028 (
            .O(N__50579),
            .I(N__50540));
    InMux I__12027 (
            .O(N__50578),
            .I(N__50535));
    LocalMux I__12026 (
            .O(N__50573),
            .I(N__50532));
    InMux I__12025 (
            .O(N__50572),
            .I(N__50527));
    InMux I__12024 (
            .O(N__50571),
            .I(N__50527));
    LocalMux I__12023 (
            .O(N__50566),
            .I(N__50522));
    LocalMux I__12022 (
            .O(N__50557),
            .I(N__50522));
    Span4Mux_v I__12021 (
            .O(N__50552),
            .I(N__50515));
    LocalMux I__12020 (
            .O(N__50549),
            .I(N__50515));
    Span4Mux_v I__12019 (
            .O(N__50546),
            .I(N__50515));
    LocalMux I__12018 (
            .O(N__50543),
            .I(N__50510));
    LocalMux I__12017 (
            .O(N__50540),
            .I(N__50510));
    InMux I__12016 (
            .O(N__50539),
            .I(N__50505));
    InMux I__12015 (
            .O(N__50538),
            .I(N__50505));
    LocalMux I__12014 (
            .O(N__50535),
            .I(N__50498));
    Span4Mux_h I__12013 (
            .O(N__50532),
            .I(N__50498));
    LocalMux I__12012 (
            .O(N__50527),
            .I(N__50498));
    Span4Mux_h I__12011 (
            .O(N__50522),
            .I(N__50495));
    Span4Mux_h I__12010 (
            .O(N__50515),
            .I(N__50490));
    Span4Mux_v I__12009 (
            .O(N__50510),
            .I(N__50490));
    LocalMux I__12008 (
            .O(N__50505),
            .I(comm_index_2));
    Odrv4 I__12007 (
            .O(N__50498),
            .I(comm_index_2));
    Odrv4 I__12006 (
            .O(N__50495),
            .I(comm_index_2));
    Odrv4 I__12005 (
            .O(N__50490),
            .I(comm_index_2));
    CascadeMux I__12004 (
            .O(N__50481),
            .I(n22267_cascade_));
    InMux I__12003 (
            .O(N__50478),
            .I(N__50474));
    CascadeMux I__12002 (
            .O(N__50477),
            .I(N__50471));
    LocalMux I__12001 (
            .O(N__50474),
            .I(N__50468));
    InMux I__12000 (
            .O(N__50471),
            .I(N__50465));
    Span4Mux_h I__11999 (
            .O(N__50468),
            .I(N__50462));
    LocalMux I__11998 (
            .O(N__50465),
            .I(data_idxvec_7));
    Odrv4 I__11997 (
            .O(N__50462),
            .I(data_idxvec_7));
    InMux I__11996 (
            .O(N__50457),
            .I(N__50454));
    LocalMux I__11995 (
            .O(N__50454),
            .I(N__50449));
    InMux I__11994 (
            .O(N__50453),
            .I(N__50446));
    InMux I__11993 (
            .O(N__50452),
            .I(N__50443));
    Span12Mux_h I__11992 (
            .O(N__50449),
            .I(N__50440));
    LocalMux I__11991 (
            .O(N__50446),
            .I(data_cntvec_7));
    LocalMux I__11990 (
            .O(N__50443),
            .I(data_cntvec_7));
    Odrv12 I__11989 (
            .O(N__50440),
            .I(data_cntvec_7));
    InMux I__11988 (
            .O(N__50433),
            .I(N__50430));
    LocalMux I__11987 (
            .O(N__50430),
            .I(N__50427));
    Span12Mux_h I__11986 (
            .O(N__50427),
            .I(N__50424));
    Odrv12 I__11985 (
            .O(N__50424),
            .I(buf_data_iac_15));
    CascadeMux I__11984 (
            .O(N__50421),
            .I(n26_adj_1502_cascade_));
    InMux I__11983 (
            .O(N__50418),
            .I(N__50415));
    LocalMux I__11982 (
            .O(N__50415),
            .I(n21055));
    CascadeMux I__11981 (
            .O(N__50412),
            .I(N__50405));
    InMux I__11980 (
            .O(N__50411),
            .I(N__50402));
    InMux I__11979 (
            .O(N__50410),
            .I(N__50399));
    InMux I__11978 (
            .O(N__50409),
            .I(N__50396));
    InMux I__11977 (
            .O(N__50408),
            .I(N__50393));
    InMux I__11976 (
            .O(N__50405),
            .I(N__50390));
    LocalMux I__11975 (
            .O(N__50402),
            .I(N__50384));
    LocalMux I__11974 (
            .O(N__50399),
            .I(N__50384));
    LocalMux I__11973 (
            .O(N__50396),
            .I(N__50381));
    LocalMux I__11972 (
            .O(N__50393),
            .I(N__50377));
    LocalMux I__11971 (
            .O(N__50390),
            .I(N__50374));
    InMux I__11970 (
            .O(N__50389),
            .I(N__50371));
    Span4Mux_v I__11969 (
            .O(N__50384),
            .I(N__50366));
    Span4Mux_h I__11968 (
            .O(N__50381),
            .I(N__50366));
    InMux I__11967 (
            .O(N__50380),
            .I(N__50363));
    Span4Mux_v I__11966 (
            .O(N__50377),
            .I(N__50358));
    Span4Mux_v I__11965 (
            .O(N__50374),
            .I(N__50358));
    LocalMux I__11964 (
            .O(N__50371),
            .I(N__50355));
    Span4Mux_h I__11963 (
            .O(N__50366),
            .I(N__50350));
    LocalMux I__11962 (
            .O(N__50363),
            .I(N__50350));
    Sp12to4 I__11961 (
            .O(N__50358),
            .I(N__50346));
    Span4Mux_v I__11960 (
            .O(N__50355),
            .I(N__50343));
    Span4Mux_v I__11959 (
            .O(N__50350),
            .I(N__50340));
    InMux I__11958 (
            .O(N__50349),
            .I(N__50337));
    Odrv12 I__11957 (
            .O(N__50346),
            .I(comm_rx_buf_7));
    Odrv4 I__11956 (
            .O(N__50343),
            .I(comm_rx_buf_7));
    Odrv4 I__11955 (
            .O(N__50340),
            .I(comm_rx_buf_7));
    LocalMux I__11954 (
            .O(N__50337),
            .I(comm_rx_buf_7));
    InMux I__11953 (
            .O(N__50328),
            .I(N__50325));
    LocalMux I__11952 (
            .O(N__50325),
            .I(n22270));
    CascadeMux I__11951 (
            .O(N__50322),
            .I(N__50315));
    CascadeMux I__11950 (
            .O(N__50321),
            .I(N__50312));
    CascadeMux I__11949 (
            .O(N__50320),
            .I(N__50309));
    InMux I__11948 (
            .O(N__50319),
            .I(N__50306));
    InMux I__11947 (
            .O(N__50318),
            .I(N__50303));
    InMux I__11946 (
            .O(N__50315),
            .I(N__50299));
    InMux I__11945 (
            .O(N__50312),
            .I(N__50296));
    InMux I__11944 (
            .O(N__50309),
            .I(N__50293));
    LocalMux I__11943 (
            .O(N__50306),
            .I(N__50290));
    LocalMux I__11942 (
            .O(N__50303),
            .I(N__50287));
    InMux I__11941 (
            .O(N__50302),
            .I(N__50284));
    LocalMux I__11940 (
            .O(N__50299),
            .I(N__50281));
    LocalMux I__11939 (
            .O(N__50296),
            .I(N__50278));
    LocalMux I__11938 (
            .O(N__50293),
            .I(N__50275));
    Span4Mux_v I__11937 (
            .O(N__50290),
            .I(N__50272));
    Span4Mux_h I__11936 (
            .O(N__50287),
            .I(N__50267));
    LocalMux I__11935 (
            .O(N__50284),
            .I(N__50267));
    Span4Mux_h I__11934 (
            .O(N__50281),
            .I(N__50264));
    Span4Mux_v I__11933 (
            .O(N__50278),
            .I(N__50257));
    Span4Mux_v I__11932 (
            .O(N__50275),
            .I(N__50257));
    Span4Mux_h I__11931 (
            .O(N__50272),
            .I(N__50257));
    Span4Mux_h I__11930 (
            .O(N__50267),
            .I(N__50254));
    Span4Mux_v I__11929 (
            .O(N__50264),
            .I(N__50251));
    Sp12to4 I__11928 (
            .O(N__50257),
            .I(N__50248));
    Span4Mux_v I__11927 (
            .O(N__50254),
            .I(N__50245));
    Odrv4 I__11926 (
            .O(N__50251),
            .I(comm_buf_1_7));
    Odrv12 I__11925 (
            .O(N__50248),
            .I(comm_buf_1_7));
    Odrv4 I__11924 (
            .O(N__50245),
            .I(comm_buf_1_7));
    InMux I__11923 (
            .O(N__50238),
            .I(N__50235));
    LocalMux I__11922 (
            .O(N__50235),
            .I(N__50232));
    Span12Mux_h I__11921 (
            .O(N__50232),
            .I(N__50228));
    InMux I__11920 (
            .O(N__50231),
            .I(N__50225));
    Odrv12 I__11919 (
            .O(N__50228),
            .I(buf_adcdata_vdc_15));
    LocalMux I__11918 (
            .O(N__50225),
            .I(buf_adcdata_vdc_15));
    InMux I__11917 (
            .O(N__50220),
            .I(N__50217));
    LocalMux I__11916 (
            .O(N__50217),
            .I(N__50213));
    InMux I__11915 (
            .O(N__50216),
            .I(N__50210));
    Span4Mux_v I__11914 (
            .O(N__50213),
            .I(N__50205));
    LocalMux I__11913 (
            .O(N__50210),
            .I(N__50205));
    Span4Mux_h I__11912 (
            .O(N__50205),
            .I(N__50202));
    Span4Mux_h I__11911 (
            .O(N__50202),
            .I(N__50198));
    InMux I__11910 (
            .O(N__50201),
            .I(N__50195));
    Span4Mux_h I__11909 (
            .O(N__50198),
            .I(N__50192));
    LocalMux I__11908 (
            .O(N__50195),
            .I(buf_adcdata_vac_15));
    Odrv4 I__11907 (
            .O(N__50192),
            .I(buf_adcdata_vac_15));
    CascadeMux I__11906 (
            .O(N__50187),
            .I(n19_adj_1503_cascade_));
    InMux I__11905 (
            .O(N__50184),
            .I(N__50181));
    LocalMux I__11904 (
            .O(N__50181),
            .I(N__50178));
    Span12Mux_s11_h I__11903 (
            .O(N__50178),
            .I(N__50174));
    CascadeMux I__11902 (
            .O(N__50177),
            .I(N__50171));
    Span12Mux_h I__11901 (
            .O(N__50174),
            .I(N__50168));
    InMux I__11900 (
            .O(N__50171),
            .I(N__50165));
    Odrv12 I__11899 (
            .O(N__50168),
            .I(buf_readRTD_7));
    LocalMux I__11898 (
            .O(N__50165),
            .I(buf_readRTD_7));
    InMux I__11897 (
            .O(N__50160),
            .I(N__50157));
    LocalMux I__11896 (
            .O(N__50157),
            .I(n21049));
    InMux I__11895 (
            .O(N__50154),
            .I(N__50151));
    LocalMux I__11894 (
            .O(N__50151),
            .I(N__50148));
    Span4Mux_v I__11893 (
            .O(N__50148),
            .I(N__50145));
    Span4Mux_h I__11892 (
            .O(N__50145),
            .I(N__50142));
    Span4Mux_h I__11891 (
            .O(N__50142),
            .I(N__50138));
    CascadeMux I__11890 (
            .O(N__50141),
            .I(N__50135));
    Span4Mux_h I__11889 (
            .O(N__50138),
            .I(N__50132));
    InMux I__11888 (
            .O(N__50135),
            .I(N__50129));
    Odrv4 I__11887 (
            .O(N__50132),
            .I(buf_readRTD_3));
    LocalMux I__11886 (
            .O(N__50129),
            .I(buf_readRTD_3));
    InMux I__11885 (
            .O(N__50124),
            .I(N__50121));
    LocalMux I__11884 (
            .O(N__50121),
            .I(N__50118));
    Span4Mux_h I__11883 (
            .O(N__50118),
            .I(N__50114));
    CascadeMux I__11882 (
            .O(N__50117),
            .I(N__50110));
    Span4Mux_v I__11881 (
            .O(N__50114),
            .I(N__50107));
    CascadeMux I__11880 (
            .O(N__50113),
            .I(N__50104));
    InMux I__11879 (
            .O(N__50110),
            .I(N__50101));
    Span4Mux_h I__11878 (
            .O(N__50107),
            .I(N__50098));
    InMux I__11877 (
            .O(N__50104),
            .I(N__50095));
    LocalMux I__11876 (
            .O(N__50101),
            .I(req_data_cnt_3));
    Odrv4 I__11875 (
            .O(N__50098),
            .I(req_data_cnt_3));
    LocalMux I__11874 (
            .O(N__50095),
            .I(req_data_cnt_3));
    InMux I__11873 (
            .O(N__50088),
            .I(N__50084));
    CascadeMux I__11872 (
            .O(N__50087),
            .I(N__50081));
    LocalMux I__11871 (
            .O(N__50084),
            .I(N__50077));
    InMux I__11870 (
            .O(N__50081),
            .I(N__50074));
    InMux I__11869 (
            .O(N__50080),
            .I(N__50071));
    Span12Mux_h I__11868 (
            .O(N__50077),
            .I(N__50068));
    LocalMux I__11867 (
            .O(N__50074),
            .I(N__50065));
    LocalMux I__11866 (
            .O(N__50071),
            .I(acadc_skipCount_3));
    Odrv12 I__11865 (
            .O(N__50068),
            .I(acadc_skipCount_3));
    Odrv4 I__11864 (
            .O(N__50065),
            .I(acadc_skipCount_3));
    InMux I__11863 (
            .O(N__50058),
            .I(N__50055));
    LocalMux I__11862 (
            .O(N__50055),
            .I(n12_adj_1548));
    InMux I__11861 (
            .O(N__50052),
            .I(N__50048));
    CascadeMux I__11860 (
            .O(N__50051),
            .I(N__50042));
    LocalMux I__11859 (
            .O(N__50048),
            .I(N__50039));
    CascadeMux I__11858 (
            .O(N__50047),
            .I(N__50032));
    CascadeMux I__11857 (
            .O(N__50046),
            .I(N__50027));
    InMux I__11856 (
            .O(N__50045),
            .I(N__50023));
    InMux I__11855 (
            .O(N__50042),
            .I(N__50020));
    Span4Mux_h I__11854 (
            .O(N__50039),
            .I(N__50017));
    InMux I__11853 (
            .O(N__50038),
            .I(N__50014));
    CascadeMux I__11852 (
            .O(N__50037),
            .I(N__50009));
    InMux I__11851 (
            .O(N__50036),
            .I(N__50001));
    InMux I__11850 (
            .O(N__50035),
            .I(N__50001));
    InMux I__11849 (
            .O(N__50032),
            .I(N__50001));
    CascadeMux I__11848 (
            .O(N__50031),
            .I(N__49998));
    CascadeMux I__11847 (
            .O(N__50030),
            .I(N__49995));
    InMux I__11846 (
            .O(N__50027),
            .I(N__49990));
    InMux I__11845 (
            .O(N__50026),
            .I(N__49987));
    LocalMux I__11844 (
            .O(N__50023),
            .I(N__49984));
    LocalMux I__11843 (
            .O(N__50020),
            .I(N__49981));
    Span4Mux_v I__11842 (
            .O(N__50017),
            .I(N__49976));
    LocalMux I__11841 (
            .O(N__50014),
            .I(N__49976));
    InMux I__11840 (
            .O(N__50013),
            .I(N__49973));
    InMux I__11839 (
            .O(N__50012),
            .I(N__49966));
    InMux I__11838 (
            .O(N__50009),
            .I(N__49966));
    InMux I__11837 (
            .O(N__50008),
            .I(N__49966));
    LocalMux I__11836 (
            .O(N__50001),
            .I(N__49961));
    InMux I__11835 (
            .O(N__49998),
            .I(N__49952));
    InMux I__11834 (
            .O(N__49995),
            .I(N__49952));
    InMux I__11833 (
            .O(N__49994),
            .I(N__49952));
    InMux I__11832 (
            .O(N__49993),
            .I(N__49952));
    LocalMux I__11831 (
            .O(N__49990),
            .I(N__49949));
    LocalMux I__11830 (
            .O(N__49987),
            .I(N__49946));
    Span4Mux_h I__11829 (
            .O(N__49984),
            .I(N__49941));
    Span4Mux_h I__11828 (
            .O(N__49981),
            .I(N__49941));
    Span4Mux_v I__11827 (
            .O(N__49976),
            .I(N__49936));
    LocalMux I__11826 (
            .O(N__49973),
            .I(N__49936));
    LocalMux I__11825 (
            .O(N__49966),
            .I(N__49933));
    InMux I__11824 (
            .O(N__49965),
            .I(N__49928));
    InMux I__11823 (
            .O(N__49964),
            .I(N__49928));
    Span4Mux_v I__11822 (
            .O(N__49961),
            .I(N__49921));
    LocalMux I__11821 (
            .O(N__49952),
            .I(N__49921));
    Span4Mux_v I__11820 (
            .O(N__49949),
            .I(N__49921));
    Span4Mux_v I__11819 (
            .O(N__49946),
            .I(N__49918));
    Span4Mux_v I__11818 (
            .O(N__49941),
            .I(N__49913));
    Span4Mux_h I__11817 (
            .O(N__49936),
            .I(N__49913));
    Span12Mux_v I__11816 (
            .O(N__49933),
            .I(N__49908));
    LocalMux I__11815 (
            .O(N__49928),
            .I(N__49908));
    Sp12to4 I__11814 (
            .O(N__49921),
            .I(N__49905));
    Sp12to4 I__11813 (
            .O(N__49918),
            .I(N__49900));
    Sp12to4 I__11812 (
            .O(N__49913),
            .I(N__49900));
    Span12Mux_v I__11811 (
            .O(N__49908),
            .I(N__49897));
    Span12Mux_h I__11810 (
            .O(N__49905),
            .I(N__49894));
    Span12Mux_v I__11809 (
            .O(N__49900),
            .I(N__49891));
    Span12Mux_h I__11808 (
            .O(N__49897),
            .I(N__49886));
    Span12Mux_v I__11807 (
            .O(N__49894),
            .I(N__49886));
    Odrv12 I__11806 (
            .O(N__49891),
            .I(ICE_SPI_CE0));
    Odrv12 I__11805 (
            .O(N__49886),
            .I(ICE_SPI_CE0));
    InMux I__11804 (
            .O(N__49881),
            .I(N__49878));
    LocalMux I__11803 (
            .O(N__49878),
            .I(N__49868));
    CascadeMux I__11802 (
            .O(N__49877),
            .I(N__49864));
    InMux I__11801 (
            .O(N__49876),
            .I(N__49859));
    InMux I__11800 (
            .O(N__49875),
            .I(N__49859));
    InMux I__11799 (
            .O(N__49874),
            .I(N__49850));
    InMux I__11798 (
            .O(N__49873),
            .I(N__49850));
    InMux I__11797 (
            .O(N__49872),
            .I(N__49850));
    InMux I__11796 (
            .O(N__49871),
            .I(N__49850));
    Span4Mux_v I__11795 (
            .O(N__49868),
            .I(N__49843));
    InMux I__11794 (
            .O(N__49867),
            .I(N__49840));
    InMux I__11793 (
            .O(N__49864),
            .I(N__49837));
    LocalMux I__11792 (
            .O(N__49859),
            .I(N__49832));
    LocalMux I__11791 (
            .O(N__49850),
            .I(N__49832));
    InMux I__11790 (
            .O(N__49849),
            .I(N__49829));
    InMux I__11789 (
            .O(N__49848),
            .I(N__49826));
    InMux I__11788 (
            .O(N__49847),
            .I(N__49823));
    InMux I__11787 (
            .O(N__49846),
            .I(N__49820));
    Sp12to4 I__11786 (
            .O(N__49843),
            .I(N__49813));
    LocalMux I__11785 (
            .O(N__49840),
            .I(N__49813));
    LocalMux I__11784 (
            .O(N__49837),
            .I(N__49813));
    Odrv4 I__11783 (
            .O(N__49832),
            .I(comm_data_vld));
    LocalMux I__11782 (
            .O(N__49829),
            .I(comm_data_vld));
    LocalMux I__11781 (
            .O(N__49826),
            .I(comm_data_vld));
    LocalMux I__11780 (
            .O(N__49823),
            .I(comm_data_vld));
    LocalMux I__11779 (
            .O(N__49820),
            .I(comm_data_vld));
    Odrv12 I__11778 (
            .O(N__49813),
            .I(comm_data_vld));
    InMux I__11777 (
            .O(N__49800),
            .I(N__49797));
    LocalMux I__11776 (
            .O(N__49797),
            .I(n18984));
    InMux I__11775 (
            .O(N__49794),
            .I(N__49790));
    InMux I__11774 (
            .O(N__49793),
            .I(N__49787));
    LocalMux I__11773 (
            .O(N__49790),
            .I(N__49781));
    LocalMux I__11772 (
            .O(N__49787),
            .I(N__49781));
    InMux I__11771 (
            .O(N__49786),
            .I(N__49778));
    Span4Mux_v I__11770 (
            .O(N__49781),
            .I(N__49773));
    LocalMux I__11769 (
            .O(N__49778),
            .I(N__49770));
    InMux I__11768 (
            .O(N__49777),
            .I(N__49767));
    InMux I__11767 (
            .O(N__49776),
            .I(N__49764));
    Span4Mux_h I__11766 (
            .O(N__49773),
            .I(N__49761));
    Sp12to4 I__11765 (
            .O(N__49770),
            .I(N__49756));
    LocalMux I__11764 (
            .O(N__49767),
            .I(N__49756));
    LocalMux I__11763 (
            .O(N__49764),
            .I(comm_cmd_4));
    Odrv4 I__11762 (
            .O(N__49761),
            .I(comm_cmd_4));
    Odrv12 I__11761 (
            .O(N__49756),
            .I(comm_cmd_4));
    InMux I__11760 (
            .O(N__49749),
            .I(N__49745));
    InMux I__11759 (
            .O(N__49748),
            .I(N__49742));
    LocalMux I__11758 (
            .O(N__49745),
            .I(N__49737));
    LocalMux I__11757 (
            .O(N__49742),
            .I(N__49737));
    Span4Mux_h I__11756 (
            .O(N__49737),
            .I(N__49734));
    Span4Mux_h I__11755 (
            .O(N__49734),
            .I(N__49728));
    InMux I__11754 (
            .O(N__49733),
            .I(N__49723));
    InMux I__11753 (
            .O(N__49732),
            .I(N__49723));
    InMux I__11752 (
            .O(N__49731),
            .I(N__49720));
    Odrv4 I__11751 (
            .O(N__49728),
            .I(comm_cmd_6));
    LocalMux I__11750 (
            .O(N__49723),
            .I(comm_cmd_6));
    LocalMux I__11749 (
            .O(N__49720),
            .I(comm_cmd_6));
    InMux I__11748 (
            .O(N__49713),
            .I(N__49709));
    InMux I__11747 (
            .O(N__49712),
            .I(N__49706));
    LocalMux I__11746 (
            .O(N__49709),
            .I(N__49701));
    LocalMux I__11745 (
            .O(N__49706),
            .I(N__49701));
    Span4Mux_h I__11744 (
            .O(N__49701),
            .I(N__49697));
    InMux I__11743 (
            .O(N__49700),
            .I(N__49692));
    Span4Mux_v I__11742 (
            .O(N__49697),
            .I(N__49689));
    InMux I__11741 (
            .O(N__49696),
            .I(N__49686));
    InMux I__11740 (
            .O(N__49695),
            .I(N__49683));
    LocalMux I__11739 (
            .O(N__49692),
            .I(comm_cmd_5));
    Odrv4 I__11738 (
            .O(N__49689),
            .I(comm_cmd_5));
    LocalMux I__11737 (
            .O(N__49686),
            .I(comm_cmd_5));
    LocalMux I__11736 (
            .O(N__49683),
            .I(comm_cmd_5));
    CascadeMux I__11735 (
            .O(N__49674),
            .I(N__49671));
    InMux I__11734 (
            .O(N__49671),
            .I(N__49668));
    LocalMux I__11733 (
            .O(N__49668),
            .I(n21546));
    InMux I__11732 (
            .O(N__49665),
            .I(N__49662));
    LocalMux I__11731 (
            .O(N__49662),
            .I(N__49659));
    Odrv4 I__11730 (
            .O(N__49659),
            .I(n12092));
    InMux I__11729 (
            .O(N__49656),
            .I(N__49650));
    InMux I__11728 (
            .O(N__49655),
            .I(N__49643));
    InMux I__11727 (
            .O(N__49654),
            .I(N__49643));
    InMux I__11726 (
            .O(N__49653),
            .I(N__49643));
    LocalMux I__11725 (
            .O(N__49650),
            .I(N__49640));
    LocalMux I__11724 (
            .O(N__49643),
            .I(N__49637));
    Span4Mux_h I__11723 (
            .O(N__49640),
            .I(N__49634));
    Span4Mux_v I__11722 (
            .O(N__49637),
            .I(N__49629));
    Span4Mux_h I__11721 (
            .O(N__49634),
            .I(N__49629));
    Span4Mux_h I__11720 (
            .O(N__49629),
            .I(N__49626));
    Odrv4 I__11719 (
            .O(N__49626),
            .I(n12219));
    InMux I__11718 (
            .O(N__49623),
            .I(N__49620));
    LocalMux I__11717 (
            .O(N__49620),
            .I(N__49616));
    InMux I__11716 (
            .O(N__49619),
            .I(N__49613));
    Span4Mux_h I__11715 (
            .O(N__49616),
            .I(N__49610));
    LocalMux I__11714 (
            .O(N__49613),
            .I(n9255));
    Odrv4 I__11713 (
            .O(N__49610),
            .I(n9255));
    CascadeMux I__11712 (
            .O(N__49605),
            .I(n11853_cascade_));
    InMux I__11711 (
            .O(N__49602),
            .I(N__49598));
    InMux I__11710 (
            .O(N__49601),
            .I(N__49595));
    LocalMux I__11709 (
            .O(N__49598),
            .I(N__49592));
    LocalMux I__11708 (
            .O(N__49595),
            .I(N__49582));
    Span4Mux_v I__11707 (
            .O(N__49592),
            .I(N__49579));
    CascadeMux I__11706 (
            .O(N__49591),
            .I(N__49576));
    InMux I__11705 (
            .O(N__49590),
            .I(N__49567));
    InMux I__11704 (
            .O(N__49589),
            .I(N__49567));
    InMux I__11703 (
            .O(N__49588),
            .I(N__49567));
    InMux I__11702 (
            .O(N__49587),
            .I(N__49563));
    InMux I__11701 (
            .O(N__49586),
            .I(N__49559));
    InMux I__11700 (
            .O(N__49585),
            .I(N__49556));
    Span4Mux_v I__11699 (
            .O(N__49582),
            .I(N__49553));
    Span4Mux_h I__11698 (
            .O(N__49579),
            .I(N__49550));
    InMux I__11697 (
            .O(N__49576),
            .I(N__49543));
    InMux I__11696 (
            .O(N__49575),
            .I(N__49543));
    InMux I__11695 (
            .O(N__49574),
            .I(N__49543));
    LocalMux I__11694 (
            .O(N__49567),
            .I(N__49540));
    InMux I__11693 (
            .O(N__49566),
            .I(N__49537));
    LocalMux I__11692 (
            .O(N__49563),
            .I(N__49534));
    InMux I__11691 (
            .O(N__49562),
            .I(N__49531));
    LocalMux I__11690 (
            .O(N__49559),
            .I(N__49526));
    LocalMux I__11689 (
            .O(N__49556),
            .I(N__49526));
    Span4Mux_h I__11688 (
            .O(N__49553),
            .I(N__49519));
    Span4Mux_v I__11687 (
            .O(N__49550),
            .I(N__49519));
    LocalMux I__11686 (
            .O(N__49543),
            .I(N__49519));
    Span4Mux_h I__11685 (
            .O(N__49540),
            .I(N__49512));
    LocalMux I__11684 (
            .O(N__49537),
            .I(N__49512));
    Span4Mux_h I__11683 (
            .O(N__49534),
            .I(N__49512));
    LocalMux I__11682 (
            .O(N__49531),
            .I(n12226));
    Odrv12 I__11681 (
            .O(N__49526),
            .I(n12226));
    Odrv4 I__11680 (
            .O(N__49519),
            .I(n12226));
    Odrv4 I__11679 (
            .O(N__49512),
            .I(n12226));
    InMux I__11678 (
            .O(N__49503),
            .I(N__49500));
    LocalMux I__11677 (
            .O(N__49500),
            .I(N__49478));
    InMux I__11676 (
            .O(N__49499),
            .I(N__49471));
    InMux I__11675 (
            .O(N__49498),
            .I(N__49471));
    InMux I__11674 (
            .O(N__49497),
            .I(N__49471));
    CascadeMux I__11673 (
            .O(N__49496),
            .I(N__49468));
    CascadeMux I__11672 (
            .O(N__49495),
            .I(N__49465));
    CascadeMux I__11671 (
            .O(N__49494),
            .I(N__49460));
    InMux I__11670 (
            .O(N__49493),
            .I(N__49457));
    InMux I__11669 (
            .O(N__49492),
            .I(N__49454));
    InMux I__11668 (
            .O(N__49491),
            .I(N__49449));
    InMux I__11667 (
            .O(N__49490),
            .I(N__49449));
    InMux I__11666 (
            .O(N__49489),
            .I(N__49446));
    InMux I__11665 (
            .O(N__49488),
            .I(N__49439));
    InMux I__11664 (
            .O(N__49487),
            .I(N__49439));
    InMux I__11663 (
            .O(N__49486),
            .I(N__49439));
    InMux I__11662 (
            .O(N__49485),
            .I(N__49430));
    InMux I__11661 (
            .O(N__49484),
            .I(N__49430));
    InMux I__11660 (
            .O(N__49483),
            .I(N__49430));
    InMux I__11659 (
            .O(N__49482),
            .I(N__49430));
    InMux I__11658 (
            .O(N__49481),
            .I(N__49427));
    Span4Mux_v I__11657 (
            .O(N__49478),
            .I(N__49420));
    LocalMux I__11656 (
            .O(N__49471),
            .I(N__49420));
    InMux I__11655 (
            .O(N__49468),
            .I(N__49417));
    InMux I__11654 (
            .O(N__49465),
            .I(N__49414));
    InMux I__11653 (
            .O(N__49464),
            .I(N__49394));
    InMux I__11652 (
            .O(N__49463),
            .I(N__49394));
    InMux I__11651 (
            .O(N__49460),
            .I(N__49394));
    LocalMux I__11650 (
            .O(N__49457),
            .I(N__49391));
    LocalMux I__11649 (
            .O(N__49454),
            .I(N__49388));
    LocalMux I__11648 (
            .O(N__49449),
            .I(N__49385));
    LocalMux I__11647 (
            .O(N__49446),
            .I(N__49380));
    LocalMux I__11646 (
            .O(N__49439),
            .I(N__49380));
    LocalMux I__11645 (
            .O(N__49430),
            .I(N__49375));
    LocalMux I__11644 (
            .O(N__49427),
            .I(N__49375));
    InMux I__11643 (
            .O(N__49426),
            .I(N__49372));
    InMux I__11642 (
            .O(N__49425),
            .I(N__49369));
    Span4Mux_h I__11641 (
            .O(N__49420),
            .I(N__49362));
    LocalMux I__11640 (
            .O(N__49417),
            .I(N__49362));
    LocalMux I__11639 (
            .O(N__49414),
            .I(N__49362));
    InMux I__11638 (
            .O(N__49413),
            .I(N__49353));
    InMux I__11637 (
            .O(N__49412),
            .I(N__49353));
    InMux I__11636 (
            .O(N__49411),
            .I(N__49353));
    InMux I__11635 (
            .O(N__49410),
            .I(N__49353));
    InMux I__11634 (
            .O(N__49409),
            .I(N__49348));
    InMux I__11633 (
            .O(N__49408),
            .I(N__49348));
    InMux I__11632 (
            .O(N__49407),
            .I(N__49339));
    InMux I__11631 (
            .O(N__49406),
            .I(N__49339));
    InMux I__11630 (
            .O(N__49405),
            .I(N__49339));
    InMux I__11629 (
            .O(N__49404),
            .I(N__49339));
    InMux I__11628 (
            .O(N__49403),
            .I(N__49332));
    InMux I__11627 (
            .O(N__49402),
            .I(N__49332));
    InMux I__11626 (
            .O(N__49401),
            .I(N__49332));
    LocalMux I__11625 (
            .O(N__49394),
            .I(N__49327));
    Span12Mux_v I__11624 (
            .O(N__49391),
            .I(N__49327));
    Span12Mux_h I__11623 (
            .O(N__49388),
            .I(N__49324));
    Span4Mux_h I__11622 (
            .O(N__49385),
            .I(N__49317));
    Span4Mux_h I__11621 (
            .O(N__49380),
            .I(N__49317));
    Span4Mux_v I__11620 (
            .O(N__49375),
            .I(N__49317));
    LocalMux I__11619 (
            .O(N__49372),
            .I(N__49310));
    LocalMux I__11618 (
            .O(N__49369),
            .I(N__49310));
    Sp12to4 I__11617 (
            .O(N__49362),
            .I(N__49310));
    LocalMux I__11616 (
            .O(N__49353),
            .I(comm_state_0));
    LocalMux I__11615 (
            .O(N__49348),
            .I(comm_state_0));
    LocalMux I__11614 (
            .O(N__49339),
            .I(comm_state_0));
    LocalMux I__11613 (
            .O(N__49332),
            .I(comm_state_0));
    Odrv12 I__11612 (
            .O(N__49327),
            .I(comm_state_0));
    Odrv12 I__11611 (
            .O(N__49324),
            .I(comm_state_0));
    Odrv4 I__11610 (
            .O(N__49317),
            .I(comm_state_0));
    Odrv12 I__11609 (
            .O(N__49310),
            .I(comm_state_0));
    InMux I__11608 (
            .O(N__49293),
            .I(N__49289));
    InMux I__11607 (
            .O(N__49292),
            .I(N__49286));
    LocalMux I__11606 (
            .O(N__49289),
            .I(n18991));
    LocalMux I__11605 (
            .O(N__49286),
            .I(n18991));
    InMux I__11604 (
            .O(N__49281),
            .I(N__49272));
    InMux I__11603 (
            .O(N__49280),
            .I(N__49272));
    InMux I__11602 (
            .O(N__49279),
            .I(N__49272));
    LocalMux I__11601 (
            .O(N__49272),
            .I(N__49268));
    InMux I__11600 (
            .O(N__49271),
            .I(N__49265));
    Span12Mux_h I__11599 (
            .O(N__49268),
            .I(N__49262));
    LocalMux I__11598 (
            .O(N__49265),
            .I(N__49259));
    Odrv12 I__11597 (
            .O(N__49262),
            .I(n20804));
    Odrv4 I__11596 (
            .O(N__49259),
            .I(n20804));
    InMux I__11595 (
            .O(N__49254),
            .I(N__49251));
    LocalMux I__11594 (
            .O(N__49251),
            .I(N__49248));
    Span4Mux_v I__11593 (
            .O(N__49248),
            .I(N__49245));
    Span4Mux_v I__11592 (
            .O(N__49245),
            .I(N__49242));
    Odrv4 I__11591 (
            .O(N__49242),
            .I(n21341));
    CascadeMux I__11590 (
            .O(N__49239),
            .I(n21339_cascade_));
    InMux I__11589 (
            .O(N__49236),
            .I(N__49233));
    LocalMux I__11588 (
            .O(N__49233),
            .I(n38_adj_1608));
    CascadeMux I__11587 (
            .O(N__49230),
            .I(N__49227));
    InMux I__11586 (
            .O(N__49227),
            .I(N__49224));
    LocalMux I__11585 (
            .O(N__49224),
            .I(N__49221));
    Span4Mux_v I__11584 (
            .O(N__49221),
            .I(N__49218));
    Odrv4 I__11583 (
            .O(N__49218),
            .I(n21054));
    InMux I__11582 (
            .O(N__49215),
            .I(\ADC_VDC.genclk.n19723 ));
    InMux I__11581 (
            .O(N__49212),
            .I(N__49208));
    InMux I__11580 (
            .O(N__49211),
            .I(N__49205));
    LocalMux I__11579 (
            .O(N__49208),
            .I(N__49202));
    LocalMux I__11578 (
            .O(N__49205),
            .I(\ADC_VDC.genclk.t0off_15 ));
    Odrv4 I__11577 (
            .O(N__49202),
            .I(\ADC_VDC.genclk.t0off_15 ));
    CEMux I__11576 (
            .O(N__49197),
            .I(N__49193));
    CEMux I__11575 (
            .O(N__49196),
            .I(N__49190));
    LocalMux I__11574 (
            .O(N__49193),
            .I(N__49187));
    LocalMux I__11573 (
            .O(N__49190),
            .I(N__49184));
    Span4Mux_h I__11572 (
            .O(N__49187),
            .I(N__49181));
    Odrv12 I__11571 (
            .O(N__49184),
            .I(\ADC_VDC.genclk.n11735 ));
    Odrv4 I__11570 (
            .O(N__49181),
            .I(\ADC_VDC.genclk.n11735 ));
    InMux I__11569 (
            .O(N__49176),
            .I(N__49173));
    LocalMux I__11568 (
            .O(N__49173),
            .I(N__49168));
    CascadeMux I__11567 (
            .O(N__49172),
            .I(N__49164));
    InMux I__11566 (
            .O(N__49171),
            .I(N__49161));
    Span4Mux_h I__11565 (
            .O(N__49168),
            .I(N__49158));
    InMux I__11564 (
            .O(N__49167),
            .I(N__49155));
    InMux I__11563 (
            .O(N__49164),
            .I(N__49152));
    LocalMux I__11562 (
            .O(N__49161),
            .I(n14529));
    Odrv4 I__11561 (
            .O(N__49158),
            .I(n14529));
    LocalMux I__11560 (
            .O(N__49155),
            .I(n14529));
    LocalMux I__11559 (
            .O(N__49152),
            .I(n14529));
    InMux I__11558 (
            .O(N__49143),
            .I(N__49140));
    LocalMux I__11557 (
            .O(N__49140),
            .I(N__49137));
    Span4Mux_h I__11556 (
            .O(N__49137),
            .I(N__49134));
    Span4Mux_h I__11555 (
            .O(N__49134),
            .I(N__49131));
    Odrv4 I__11554 (
            .O(N__49131),
            .I(n17815));
    InMux I__11553 (
            .O(N__49128),
            .I(N__49125));
    LocalMux I__11552 (
            .O(N__49125),
            .I(N__49122));
    Span4Mux_v I__11551 (
            .O(N__49122),
            .I(N__49119));
    Span4Mux_h I__11550 (
            .O(N__49119),
            .I(N__49116));
    Odrv4 I__11549 (
            .O(N__49116),
            .I(n23_adj_1620));
    CascadeMux I__11548 (
            .O(N__49113),
            .I(n21_adj_1598_cascade_));
    InMux I__11547 (
            .O(N__49110),
            .I(N__49107));
    LocalMux I__11546 (
            .O(N__49107),
            .I(N__49104));
    Span4Mux_h I__11545 (
            .O(N__49104),
            .I(N__49101));
    Span4Mux_h I__11544 (
            .O(N__49101),
            .I(N__49098));
    Span4Mux_h I__11543 (
            .O(N__49098),
            .I(N__49095));
    Odrv4 I__11542 (
            .O(N__49095),
            .I(n17564));
    InMux I__11541 (
            .O(N__49092),
            .I(N__49089));
    LocalMux I__11540 (
            .O(N__49089),
            .I(N__49083));
    InMux I__11539 (
            .O(N__49088),
            .I(N__49080));
    InMux I__11538 (
            .O(N__49087),
            .I(N__49077));
    InMux I__11537 (
            .O(N__49086),
            .I(N__49074));
    Span4Mux_v I__11536 (
            .O(N__49083),
            .I(N__49071));
    LocalMux I__11535 (
            .O(N__49080),
            .I(N__49068));
    LocalMux I__11534 (
            .O(N__49077),
            .I(N__49063));
    LocalMux I__11533 (
            .O(N__49074),
            .I(N__49063));
    Span4Mux_h I__11532 (
            .O(N__49071),
            .I(N__49058));
    Span4Mux_v I__11531 (
            .O(N__49068),
            .I(N__49058));
    Span4Mux_h I__11530 (
            .O(N__49063),
            .I(N__49055));
    Odrv4 I__11529 (
            .O(N__49058),
            .I(n2358));
    Odrv4 I__11528 (
            .O(N__49055),
            .I(n2358));
    InMux I__11527 (
            .O(N__49050),
            .I(N__49047));
    LocalMux I__11526 (
            .O(N__49047),
            .I(N__49044));
    Sp12to4 I__11525 (
            .O(N__49044),
            .I(N__49041));
    Span12Mux_h I__11524 (
            .O(N__49041),
            .I(N__49038));
    Odrv12 I__11523 (
            .O(N__49038),
            .I(n20856));
    CascadeMux I__11522 (
            .O(N__49035),
            .I(n15_cascade_));
    CEMux I__11521 (
            .O(N__49032),
            .I(N__49029));
    LocalMux I__11520 (
            .O(N__49029),
            .I(n18_adj_1619));
    CascadeMux I__11519 (
            .O(N__49026),
            .I(N__49023));
    InMux I__11518 (
            .O(N__49023),
            .I(N__49020));
    LocalMux I__11517 (
            .O(N__49020),
            .I(n14130));
    InMux I__11516 (
            .O(N__49017),
            .I(N__49014));
    LocalMux I__11515 (
            .O(N__49014),
            .I(n20880));
    CascadeMux I__11514 (
            .O(N__49011),
            .I(n20880_cascade_));
    CascadeMux I__11513 (
            .O(N__49008),
            .I(N__49004));
    InMux I__11512 (
            .O(N__49007),
            .I(N__49001));
    InMux I__11511 (
            .O(N__49004),
            .I(N__48998));
    LocalMux I__11510 (
            .O(N__49001),
            .I(\ADC_VDC.genclk.t0off_7 ));
    LocalMux I__11509 (
            .O(N__48998),
            .I(\ADC_VDC.genclk.t0off_7 ));
    InMux I__11508 (
            .O(N__48993),
            .I(\ADC_VDC.genclk.n19715 ));
    InMux I__11507 (
            .O(N__48990),
            .I(N__48986));
    InMux I__11506 (
            .O(N__48989),
            .I(N__48983));
    LocalMux I__11505 (
            .O(N__48986),
            .I(\ADC_VDC.genclk.t0off_8 ));
    LocalMux I__11504 (
            .O(N__48983),
            .I(\ADC_VDC.genclk.t0off_8 ));
    InMux I__11503 (
            .O(N__48978),
            .I(bfn_19_8_0_));
    CascadeMux I__11502 (
            .O(N__48975),
            .I(N__48971));
    CascadeMux I__11501 (
            .O(N__48974),
            .I(N__48968));
    InMux I__11500 (
            .O(N__48971),
            .I(N__48965));
    InMux I__11499 (
            .O(N__48968),
            .I(N__48962));
    LocalMux I__11498 (
            .O(N__48965),
            .I(\ADC_VDC.genclk.t0off_9 ));
    LocalMux I__11497 (
            .O(N__48962),
            .I(\ADC_VDC.genclk.t0off_9 ));
    InMux I__11496 (
            .O(N__48957),
            .I(\ADC_VDC.genclk.n19717 ));
    InMux I__11495 (
            .O(N__48954),
            .I(N__48950));
    InMux I__11494 (
            .O(N__48953),
            .I(N__48947));
    LocalMux I__11493 (
            .O(N__48950),
            .I(\ADC_VDC.genclk.t0off_10 ));
    LocalMux I__11492 (
            .O(N__48947),
            .I(\ADC_VDC.genclk.t0off_10 ));
    InMux I__11491 (
            .O(N__48942),
            .I(\ADC_VDC.genclk.n19718 ));
    CascadeMux I__11490 (
            .O(N__48939),
            .I(N__48936));
    InMux I__11489 (
            .O(N__48936),
            .I(N__48932));
    InMux I__11488 (
            .O(N__48935),
            .I(N__48929));
    LocalMux I__11487 (
            .O(N__48932),
            .I(\ADC_VDC.genclk.t0off_11 ));
    LocalMux I__11486 (
            .O(N__48929),
            .I(\ADC_VDC.genclk.t0off_11 ));
    InMux I__11485 (
            .O(N__48924),
            .I(\ADC_VDC.genclk.n19719 ));
    InMux I__11484 (
            .O(N__48921),
            .I(N__48917));
    InMux I__11483 (
            .O(N__48920),
            .I(N__48914));
    LocalMux I__11482 (
            .O(N__48917),
            .I(\ADC_VDC.genclk.t0off_12 ));
    LocalMux I__11481 (
            .O(N__48914),
            .I(\ADC_VDC.genclk.t0off_12 ));
    InMux I__11480 (
            .O(N__48909),
            .I(\ADC_VDC.genclk.n19720 ));
    CascadeMux I__11479 (
            .O(N__48906),
            .I(N__48903));
    InMux I__11478 (
            .O(N__48903),
            .I(N__48899));
    InMux I__11477 (
            .O(N__48902),
            .I(N__48896));
    LocalMux I__11476 (
            .O(N__48899),
            .I(\ADC_VDC.genclk.t0off_13 ));
    LocalMux I__11475 (
            .O(N__48896),
            .I(\ADC_VDC.genclk.t0off_13 ));
    InMux I__11474 (
            .O(N__48891),
            .I(\ADC_VDC.genclk.n19721 ));
    InMux I__11473 (
            .O(N__48888),
            .I(N__48884));
    InMux I__11472 (
            .O(N__48887),
            .I(N__48881));
    LocalMux I__11471 (
            .O(N__48884),
            .I(\ADC_VDC.genclk.t0off_14 ));
    LocalMux I__11470 (
            .O(N__48881),
            .I(\ADC_VDC.genclk.t0off_14 ));
    InMux I__11469 (
            .O(N__48876),
            .I(\ADC_VDC.genclk.n19722 ));
    CascadeMux I__11468 (
            .O(N__48873),
            .I(N__48859));
    CascadeMux I__11467 (
            .O(N__48872),
            .I(N__48856));
    CascadeMux I__11466 (
            .O(N__48871),
            .I(N__48848));
    CascadeMux I__11465 (
            .O(N__48870),
            .I(N__48840));
    CascadeMux I__11464 (
            .O(N__48869),
            .I(N__48837));
    InMux I__11463 (
            .O(N__48868),
            .I(N__48817));
    InMux I__11462 (
            .O(N__48867),
            .I(N__48817));
    InMux I__11461 (
            .O(N__48866),
            .I(N__48817));
    InMux I__11460 (
            .O(N__48865),
            .I(N__48817));
    InMux I__11459 (
            .O(N__48864),
            .I(N__48817));
    InMux I__11458 (
            .O(N__48863),
            .I(N__48817));
    InMux I__11457 (
            .O(N__48862),
            .I(N__48817));
    InMux I__11456 (
            .O(N__48859),
            .I(N__48806));
    InMux I__11455 (
            .O(N__48856),
            .I(N__48806));
    InMux I__11454 (
            .O(N__48855),
            .I(N__48806));
    InMux I__11453 (
            .O(N__48854),
            .I(N__48806));
    InMux I__11452 (
            .O(N__48853),
            .I(N__48806));
    CascadeMux I__11451 (
            .O(N__48852),
            .I(N__48801));
    CascadeMux I__11450 (
            .O(N__48851),
            .I(N__48793));
    InMux I__11449 (
            .O(N__48848),
            .I(N__48787));
    InMux I__11448 (
            .O(N__48847),
            .I(N__48787));
    InMux I__11447 (
            .O(N__48846),
            .I(N__48779));
    InMux I__11446 (
            .O(N__48845),
            .I(N__48779));
    CascadeMux I__11445 (
            .O(N__48844),
            .I(N__48775));
    InMux I__11444 (
            .O(N__48843),
            .I(N__48769));
    InMux I__11443 (
            .O(N__48840),
            .I(N__48764));
    InMux I__11442 (
            .O(N__48837),
            .I(N__48764));
    CascadeMux I__11441 (
            .O(N__48836),
            .I(N__48761));
    CascadeMux I__11440 (
            .O(N__48835),
            .I(N__48755));
    InMux I__11439 (
            .O(N__48834),
            .I(N__48747));
    InMux I__11438 (
            .O(N__48833),
            .I(N__48747));
    InMux I__11437 (
            .O(N__48832),
            .I(N__48747));
    LocalMux I__11436 (
            .O(N__48817),
            .I(N__48742));
    LocalMux I__11435 (
            .O(N__48806),
            .I(N__48742));
    InMux I__11434 (
            .O(N__48805),
            .I(N__48735));
    InMux I__11433 (
            .O(N__48804),
            .I(N__48735));
    InMux I__11432 (
            .O(N__48801),
            .I(N__48735));
    InMux I__11431 (
            .O(N__48800),
            .I(N__48728));
    InMux I__11430 (
            .O(N__48799),
            .I(N__48728));
    InMux I__11429 (
            .O(N__48798),
            .I(N__48728));
    InMux I__11428 (
            .O(N__48797),
            .I(N__48721));
    InMux I__11427 (
            .O(N__48796),
            .I(N__48721));
    InMux I__11426 (
            .O(N__48793),
            .I(N__48721));
    InMux I__11425 (
            .O(N__48792),
            .I(N__48718));
    LocalMux I__11424 (
            .O(N__48787),
            .I(N__48715));
    InMux I__11423 (
            .O(N__48786),
            .I(N__48710));
    InMux I__11422 (
            .O(N__48785),
            .I(N__48710));
    InMux I__11421 (
            .O(N__48784),
            .I(N__48706));
    LocalMux I__11420 (
            .O(N__48779),
            .I(N__48703));
    InMux I__11419 (
            .O(N__48778),
            .I(N__48696));
    InMux I__11418 (
            .O(N__48775),
            .I(N__48696));
    InMux I__11417 (
            .O(N__48774),
            .I(N__48696));
    CascadeMux I__11416 (
            .O(N__48773),
            .I(N__48693));
    CascadeMux I__11415 (
            .O(N__48772),
            .I(N__48690));
    LocalMux I__11414 (
            .O(N__48769),
            .I(N__48684));
    LocalMux I__11413 (
            .O(N__48764),
            .I(N__48684));
    InMux I__11412 (
            .O(N__48761),
            .I(N__48681));
    InMux I__11411 (
            .O(N__48760),
            .I(N__48678));
    InMux I__11410 (
            .O(N__48759),
            .I(N__48675));
    InMux I__11409 (
            .O(N__48758),
            .I(N__48668));
    InMux I__11408 (
            .O(N__48755),
            .I(N__48668));
    InMux I__11407 (
            .O(N__48754),
            .I(N__48668));
    LocalMux I__11406 (
            .O(N__48747),
            .I(N__48657));
    Span4Mux_v I__11405 (
            .O(N__48742),
            .I(N__48657));
    LocalMux I__11404 (
            .O(N__48735),
            .I(N__48657));
    LocalMux I__11403 (
            .O(N__48728),
            .I(N__48657));
    LocalMux I__11402 (
            .O(N__48721),
            .I(N__48657));
    LocalMux I__11401 (
            .O(N__48718),
            .I(N__48654));
    Span4Mux_v I__11400 (
            .O(N__48715),
            .I(N__48651));
    LocalMux I__11399 (
            .O(N__48710),
            .I(N__48648));
    InMux I__11398 (
            .O(N__48709),
            .I(N__48645));
    LocalMux I__11397 (
            .O(N__48706),
            .I(N__48640));
    Span4Mux_h I__11396 (
            .O(N__48703),
            .I(N__48640));
    LocalMux I__11395 (
            .O(N__48696),
            .I(N__48637));
    InMux I__11394 (
            .O(N__48693),
            .I(N__48634));
    InMux I__11393 (
            .O(N__48690),
            .I(N__48629));
    InMux I__11392 (
            .O(N__48689),
            .I(N__48629));
    Span12Mux_h I__11391 (
            .O(N__48684),
            .I(N__48626));
    LocalMux I__11390 (
            .O(N__48681),
            .I(N__48613));
    LocalMux I__11389 (
            .O(N__48678),
            .I(N__48613));
    LocalMux I__11388 (
            .O(N__48675),
            .I(N__48613));
    LocalMux I__11387 (
            .O(N__48668),
            .I(N__48613));
    Span4Mux_v I__11386 (
            .O(N__48657),
            .I(N__48613));
    Span4Mux_v I__11385 (
            .O(N__48654),
            .I(N__48613));
    Sp12to4 I__11384 (
            .O(N__48651),
            .I(N__48608));
    Span12Mux_v I__11383 (
            .O(N__48648),
            .I(N__48608));
    LocalMux I__11382 (
            .O(N__48645),
            .I(adc_state_2));
    Odrv4 I__11381 (
            .O(N__48640),
            .I(adc_state_2));
    Odrv4 I__11380 (
            .O(N__48637),
            .I(adc_state_2));
    LocalMux I__11379 (
            .O(N__48634),
            .I(adc_state_2));
    LocalMux I__11378 (
            .O(N__48629),
            .I(adc_state_2));
    Odrv12 I__11377 (
            .O(N__48626),
            .I(adc_state_2));
    Odrv4 I__11376 (
            .O(N__48613),
            .I(adc_state_2));
    Odrv12 I__11375 (
            .O(N__48608),
            .I(adc_state_2));
    InMux I__11374 (
            .O(N__48591),
            .I(N__48570));
    InMux I__11373 (
            .O(N__48590),
            .I(N__48570));
    InMux I__11372 (
            .O(N__48589),
            .I(N__48539));
    InMux I__11371 (
            .O(N__48588),
            .I(N__48539));
    InMux I__11370 (
            .O(N__48587),
            .I(N__48539));
    InMux I__11369 (
            .O(N__48586),
            .I(N__48539));
    InMux I__11368 (
            .O(N__48585),
            .I(N__48539));
    InMux I__11367 (
            .O(N__48584),
            .I(N__48539));
    InMux I__11366 (
            .O(N__48583),
            .I(N__48539));
    InMux I__11365 (
            .O(N__48582),
            .I(N__48539));
    InMux I__11364 (
            .O(N__48581),
            .I(N__48531));
    InMux I__11363 (
            .O(N__48580),
            .I(N__48531));
    InMux I__11362 (
            .O(N__48579),
            .I(N__48517));
    InMux I__11361 (
            .O(N__48578),
            .I(N__48517));
    InMux I__11360 (
            .O(N__48577),
            .I(N__48517));
    InMux I__11359 (
            .O(N__48576),
            .I(N__48517));
    InMux I__11358 (
            .O(N__48575),
            .I(N__48517));
    LocalMux I__11357 (
            .O(N__48570),
            .I(N__48514));
    InMux I__11356 (
            .O(N__48569),
            .I(N__48509));
    InMux I__11355 (
            .O(N__48568),
            .I(N__48509));
    InMux I__11354 (
            .O(N__48567),
            .I(N__48502));
    InMux I__11353 (
            .O(N__48566),
            .I(N__48502));
    InMux I__11352 (
            .O(N__48565),
            .I(N__48502));
    InMux I__11351 (
            .O(N__48564),
            .I(N__48497));
    InMux I__11350 (
            .O(N__48563),
            .I(N__48497));
    InMux I__11349 (
            .O(N__48562),
            .I(N__48482));
    InMux I__11348 (
            .O(N__48561),
            .I(N__48482));
    InMux I__11347 (
            .O(N__48560),
            .I(N__48482));
    InMux I__11346 (
            .O(N__48559),
            .I(N__48482));
    InMux I__11345 (
            .O(N__48558),
            .I(N__48482));
    InMux I__11344 (
            .O(N__48557),
            .I(N__48482));
    InMux I__11343 (
            .O(N__48556),
            .I(N__48482));
    LocalMux I__11342 (
            .O(N__48539),
            .I(N__48476));
    InMux I__11341 (
            .O(N__48538),
            .I(N__48473));
    InMux I__11340 (
            .O(N__48537),
            .I(N__48470));
    InMux I__11339 (
            .O(N__48536),
            .I(N__48467));
    LocalMux I__11338 (
            .O(N__48531),
            .I(N__48461));
    InMux I__11337 (
            .O(N__48530),
            .I(N__48458));
    CascadeMux I__11336 (
            .O(N__48529),
            .I(N__48452));
    InMux I__11335 (
            .O(N__48528),
            .I(N__48449));
    LocalMux I__11334 (
            .O(N__48517),
            .I(N__48444));
    Span4Mux_v I__11333 (
            .O(N__48514),
            .I(N__48444));
    LocalMux I__11332 (
            .O(N__48509),
            .I(N__48441));
    LocalMux I__11331 (
            .O(N__48502),
            .I(N__48434));
    LocalMux I__11330 (
            .O(N__48497),
            .I(N__48434));
    LocalMux I__11329 (
            .O(N__48482),
            .I(N__48434));
    InMux I__11328 (
            .O(N__48481),
            .I(N__48431));
    InMux I__11327 (
            .O(N__48480),
            .I(N__48426));
    InMux I__11326 (
            .O(N__48479),
            .I(N__48426));
    Span4Mux_h I__11325 (
            .O(N__48476),
            .I(N__48419));
    LocalMux I__11324 (
            .O(N__48473),
            .I(N__48419));
    LocalMux I__11323 (
            .O(N__48470),
            .I(N__48419));
    LocalMux I__11322 (
            .O(N__48467),
            .I(N__48416));
    InMux I__11321 (
            .O(N__48466),
            .I(N__48409));
    InMux I__11320 (
            .O(N__48465),
            .I(N__48409));
    InMux I__11319 (
            .O(N__48464),
            .I(N__48409));
    Span4Mux_v I__11318 (
            .O(N__48461),
            .I(N__48406));
    LocalMux I__11317 (
            .O(N__48458),
            .I(N__48403));
    InMux I__11316 (
            .O(N__48457),
            .I(N__48400));
    InMux I__11315 (
            .O(N__48456),
            .I(N__48393));
    InMux I__11314 (
            .O(N__48455),
            .I(N__48393));
    InMux I__11313 (
            .O(N__48452),
            .I(N__48393));
    LocalMux I__11312 (
            .O(N__48449),
            .I(N__48384));
    Span4Mux_v I__11311 (
            .O(N__48444),
            .I(N__48384));
    Span4Mux_v I__11310 (
            .O(N__48441),
            .I(N__48384));
    Span4Mux_v I__11309 (
            .O(N__48434),
            .I(N__48384));
    LocalMux I__11308 (
            .O(N__48431),
            .I(N__48371));
    LocalMux I__11307 (
            .O(N__48426),
            .I(N__48371));
    Span4Mux_v I__11306 (
            .O(N__48419),
            .I(N__48371));
    Span4Mux_v I__11305 (
            .O(N__48416),
            .I(N__48371));
    LocalMux I__11304 (
            .O(N__48409),
            .I(N__48371));
    Span4Mux_h I__11303 (
            .O(N__48406),
            .I(N__48371));
    Odrv4 I__11302 (
            .O(N__48403),
            .I(adc_state_3));
    LocalMux I__11301 (
            .O(N__48400),
            .I(adc_state_3));
    LocalMux I__11300 (
            .O(N__48393),
            .I(adc_state_3));
    Odrv4 I__11299 (
            .O(N__48384),
            .I(adc_state_3));
    Odrv4 I__11298 (
            .O(N__48371),
            .I(adc_state_3));
    CascadeMux I__11297 (
            .O(N__48360),
            .I(\ADC_VDC.n62_cascade_ ));
    CascadeMux I__11296 (
            .O(N__48357),
            .I(N__48351));
    InMux I__11295 (
            .O(N__48356),
            .I(N__48340));
    InMux I__11294 (
            .O(N__48355),
            .I(N__48340));
    InMux I__11293 (
            .O(N__48354),
            .I(N__48331));
    InMux I__11292 (
            .O(N__48351),
            .I(N__48331));
    InMux I__11291 (
            .O(N__48350),
            .I(N__48331));
    InMux I__11290 (
            .O(N__48349),
            .I(N__48328));
    InMux I__11289 (
            .O(N__48348),
            .I(N__48323));
    InMux I__11288 (
            .O(N__48347),
            .I(N__48323));
    InMux I__11287 (
            .O(N__48346),
            .I(N__48320));
    InMux I__11286 (
            .O(N__48345),
            .I(N__48317));
    LocalMux I__11285 (
            .O(N__48340),
            .I(N__48314));
    InMux I__11284 (
            .O(N__48339),
            .I(N__48309));
    InMux I__11283 (
            .O(N__48338),
            .I(N__48309));
    LocalMux I__11282 (
            .O(N__48331),
            .I(N__48306));
    LocalMux I__11281 (
            .O(N__48328),
            .I(N__48301));
    LocalMux I__11280 (
            .O(N__48323),
            .I(N__48301));
    LocalMux I__11279 (
            .O(N__48320),
            .I(N__48292));
    LocalMux I__11278 (
            .O(N__48317),
            .I(N__48292));
    Span4Mux_v I__11277 (
            .O(N__48314),
            .I(N__48289));
    LocalMux I__11276 (
            .O(N__48309),
            .I(N__48280));
    Span4Mux_v I__11275 (
            .O(N__48306),
            .I(N__48280));
    Span4Mux_v I__11274 (
            .O(N__48301),
            .I(N__48280));
    InMux I__11273 (
            .O(N__48300),
            .I(N__48272));
    InMux I__11272 (
            .O(N__48299),
            .I(N__48269));
    InMux I__11271 (
            .O(N__48298),
            .I(N__48266));
    InMux I__11270 (
            .O(N__48297),
            .I(N__48263));
    Span4Mux_v I__11269 (
            .O(N__48292),
            .I(N__48258));
    Span4Mux_h I__11268 (
            .O(N__48289),
            .I(N__48258));
    InMux I__11267 (
            .O(N__48288),
            .I(N__48253));
    InMux I__11266 (
            .O(N__48287),
            .I(N__48253));
    Span4Mux_h I__11265 (
            .O(N__48280),
            .I(N__48250));
    InMux I__11264 (
            .O(N__48279),
            .I(N__48245));
    InMux I__11263 (
            .O(N__48278),
            .I(N__48245));
    InMux I__11262 (
            .O(N__48277),
            .I(N__48238));
    InMux I__11261 (
            .O(N__48276),
            .I(N__48238));
    InMux I__11260 (
            .O(N__48275),
            .I(N__48238));
    LocalMux I__11259 (
            .O(N__48272),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__11258 (
            .O(N__48269),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__11257 (
            .O(N__48266),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__11256 (
            .O(N__48263),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__11255 (
            .O(N__48258),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__11254 (
            .O(N__48253),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__11253 (
            .O(N__48250),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__11252 (
            .O(N__48245),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__11251 (
            .O(N__48238),
            .I(\ADC_VDC.adc_state_1 ));
    InMux I__11250 (
            .O(N__48219),
            .I(N__48216));
    LocalMux I__11249 (
            .O(N__48216),
            .I(N__48213));
    Span4Mux_h I__11248 (
            .O(N__48213),
            .I(N__48210));
    Odrv4 I__11247 (
            .O(N__48210),
            .I(\ADC_VDC.n11 ));
    InMux I__11246 (
            .O(N__48207),
            .I(N__48203));
    InMux I__11245 (
            .O(N__48206),
            .I(N__48200));
    LocalMux I__11244 (
            .O(N__48203),
            .I(\ADC_VDC.genclk.t0off_0 ));
    LocalMux I__11243 (
            .O(N__48200),
            .I(\ADC_VDC.genclk.t0off_0 ));
    InMux I__11242 (
            .O(N__48195),
            .I(bfn_19_7_0_));
    InMux I__11241 (
            .O(N__48192),
            .I(N__48188));
    InMux I__11240 (
            .O(N__48191),
            .I(N__48185));
    LocalMux I__11239 (
            .O(N__48188),
            .I(\ADC_VDC.genclk.t0off_1 ));
    LocalMux I__11238 (
            .O(N__48185),
            .I(\ADC_VDC.genclk.t0off_1 ));
    InMux I__11237 (
            .O(N__48180),
            .I(\ADC_VDC.genclk.n19709 ));
    CascadeMux I__11236 (
            .O(N__48177),
            .I(N__48174));
    InMux I__11235 (
            .O(N__48174),
            .I(N__48170));
    InMux I__11234 (
            .O(N__48173),
            .I(N__48167));
    LocalMux I__11233 (
            .O(N__48170),
            .I(\ADC_VDC.genclk.t0off_2 ));
    LocalMux I__11232 (
            .O(N__48167),
            .I(\ADC_VDC.genclk.t0off_2 ));
    InMux I__11231 (
            .O(N__48162),
            .I(\ADC_VDC.genclk.n19710 ));
    InMux I__11230 (
            .O(N__48159),
            .I(N__48155));
    InMux I__11229 (
            .O(N__48158),
            .I(N__48152));
    LocalMux I__11228 (
            .O(N__48155),
            .I(\ADC_VDC.genclk.t0off_3 ));
    LocalMux I__11227 (
            .O(N__48152),
            .I(\ADC_VDC.genclk.t0off_3 ));
    InMux I__11226 (
            .O(N__48147),
            .I(\ADC_VDC.genclk.n19711 ));
    CascadeMux I__11225 (
            .O(N__48144),
            .I(N__48140));
    CascadeMux I__11224 (
            .O(N__48143),
            .I(N__48137));
    InMux I__11223 (
            .O(N__48140),
            .I(N__48134));
    InMux I__11222 (
            .O(N__48137),
            .I(N__48131));
    LocalMux I__11221 (
            .O(N__48134),
            .I(N__48128));
    LocalMux I__11220 (
            .O(N__48131),
            .I(\ADC_VDC.genclk.t0off_4 ));
    Odrv4 I__11219 (
            .O(N__48128),
            .I(\ADC_VDC.genclk.t0off_4 ));
    InMux I__11218 (
            .O(N__48123),
            .I(\ADC_VDC.genclk.n19712 ));
    CascadeMux I__11217 (
            .O(N__48120),
            .I(N__48116));
    InMux I__11216 (
            .O(N__48119),
            .I(N__48113));
    InMux I__11215 (
            .O(N__48116),
            .I(N__48110));
    LocalMux I__11214 (
            .O(N__48113),
            .I(\ADC_VDC.genclk.t0off_5 ));
    LocalMux I__11213 (
            .O(N__48110),
            .I(\ADC_VDC.genclk.t0off_5 ));
    InMux I__11212 (
            .O(N__48105),
            .I(\ADC_VDC.genclk.n19713 ));
    CascadeMux I__11211 (
            .O(N__48102),
            .I(N__48099));
    InMux I__11210 (
            .O(N__48099),
            .I(N__48095));
    InMux I__11209 (
            .O(N__48098),
            .I(N__48092));
    LocalMux I__11208 (
            .O(N__48095),
            .I(\ADC_VDC.genclk.t0off_6 ));
    LocalMux I__11207 (
            .O(N__48092),
            .I(\ADC_VDC.genclk.t0off_6 ));
    InMux I__11206 (
            .O(N__48087),
            .I(\ADC_VDC.genclk.n19714 ));
    InMux I__11205 (
            .O(N__48084),
            .I(N__48081));
    LocalMux I__11204 (
            .O(N__48081),
            .I(N__48077));
    InMux I__11203 (
            .O(N__48080),
            .I(N__48074));
    Span4Mux_v I__11202 (
            .O(N__48077),
            .I(N__48069));
    LocalMux I__11201 (
            .O(N__48074),
            .I(N__48069));
    Span4Mux_h I__11200 (
            .O(N__48069),
            .I(N__48063));
    InMux I__11199 (
            .O(N__48068),
            .I(N__48060));
    CascadeMux I__11198 (
            .O(N__48067),
            .I(N__48056));
    InMux I__11197 (
            .O(N__48066),
            .I(N__48053));
    Span4Mux_v I__11196 (
            .O(N__48063),
            .I(N__48048));
    LocalMux I__11195 (
            .O(N__48060),
            .I(N__48048));
    InMux I__11194 (
            .O(N__48059),
            .I(N__48045));
    InMux I__11193 (
            .O(N__48056),
            .I(N__48042));
    LocalMux I__11192 (
            .O(N__48053),
            .I(N__48035));
    Span4Mux_v I__11191 (
            .O(N__48048),
            .I(N__48035));
    LocalMux I__11190 (
            .O(N__48045),
            .I(N__48035));
    LocalMux I__11189 (
            .O(N__48042),
            .I(N__48030));
    Span4Mux_h I__11188 (
            .O(N__48035),
            .I(N__48030));
    Odrv4 I__11187 (
            .O(N__48030),
            .I(comm_buf_1_2));
    InMux I__11186 (
            .O(N__48027),
            .I(N__48021));
    InMux I__11185 (
            .O(N__48026),
            .I(N__48018));
    InMux I__11184 (
            .O(N__48025),
            .I(N__48013));
    InMux I__11183 (
            .O(N__48024),
            .I(N__48013));
    LocalMux I__11182 (
            .O(N__48021),
            .I(N__48006));
    LocalMux I__11181 (
            .O(N__48018),
            .I(N__48001));
    LocalMux I__11180 (
            .O(N__48013),
            .I(N__48001));
    InMux I__11179 (
            .O(N__48012),
            .I(N__47998));
    InMux I__11178 (
            .O(N__48011),
            .I(N__47992));
    InMux I__11177 (
            .O(N__48010),
            .I(N__47987));
    InMux I__11176 (
            .O(N__48009),
            .I(N__47987));
    Span4Mux_v I__11175 (
            .O(N__48006),
            .I(N__47981));
    Span4Mux_v I__11174 (
            .O(N__48001),
            .I(N__47981));
    LocalMux I__11173 (
            .O(N__47998),
            .I(N__47978));
    InMux I__11172 (
            .O(N__47997),
            .I(N__47975));
    InMux I__11171 (
            .O(N__47996),
            .I(N__47970));
    InMux I__11170 (
            .O(N__47995),
            .I(N__47970));
    LocalMux I__11169 (
            .O(N__47992),
            .I(N__47964));
    LocalMux I__11168 (
            .O(N__47987),
            .I(N__47961));
    InMux I__11167 (
            .O(N__47986),
            .I(N__47958));
    Span4Mux_h I__11166 (
            .O(N__47981),
            .I(N__47951));
    Span4Mux_v I__11165 (
            .O(N__47978),
            .I(N__47951));
    LocalMux I__11164 (
            .O(N__47975),
            .I(N__47951));
    LocalMux I__11163 (
            .O(N__47970),
            .I(N__47948));
    InMux I__11162 (
            .O(N__47969),
            .I(N__47941));
    InMux I__11161 (
            .O(N__47968),
            .I(N__47941));
    InMux I__11160 (
            .O(N__47967),
            .I(N__47941));
    Odrv12 I__11159 (
            .O(N__47964),
            .I(n12367));
    Odrv12 I__11158 (
            .O(N__47961),
            .I(n12367));
    LocalMux I__11157 (
            .O(N__47958),
            .I(n12367));
    Odrv4 I__11156 (
            .O(N__47951),
            .I(n12367));
    Odrv4 I__11155 (
            .O(N__47948),
            .I(n12367));
    LocalMux I__11154 (
            .O(N__47941),
            .I(n12367));
    CascadeMux I__11153 (
            .O(N__47928),
            .I(N__47925));
    InMux I__11152 (
            .O(N__47925),
            .I(N__47922));
    LocalMux I__11151 (
            .O(N__47922),
            .I(N__47919));
    Span4Mux_v I__11150 (
            .O(N__47919),
            .I(N__47916));
    Span4Mux_h I__11149 (
            .O(N__47916),
            .I(N__47911));
    InMux I__11148 (
            .O(N__47915),
            .I(N__47906));
    InMux I__11147 (
            .O(N__47914),
            .I(N__47906));
    Odrv4 I__11146 (
            .O(N__47911),
            .I(buf_dds0_2));
    LocalMux I__11145 (
            .O(N__47906),
            .I(buf_dds0_2));
    CascadeMux I__11144 (
            .O(N__47901),
            .I(N__47898));
    InMux I__11143 (
            .O(N__47898),
            .I(N__47892));
    CascadeMux I__11142 (
            .O(N__47897),
            .I(N__47888));
    CascadeMux I__11141 (
            .O(N__47896),
            .I(N__47885));
    InMux I__11140 (
            .O(N__47895),
            .I(N__47882));
    LocalMux I__11139 (
            .O(N__47892),
            .I(N__47879));
    InMux I__11138 (
            .O(N__47891),
            .I(N__47875));
    InMux I__11137 (
            .O(N__47888),
            .I(N__47872));
    InMux I__11136 (
            .O(N__47885),
            .I(N__47869));
    LocalMux I__11135 (
            .O(N__47882),
            .I(N__47866));
    Span4Mux_h I__11134 (
            .O(N__47879),
            .I(N__47863));
    InMux I__11133 (
            .O(N__47878),
            .I(N__47860));
    LocalMux I__11132 (
            .O(N__47875),
            .I(N__47857));
    LocalMux I__11131 (
            .O(N__47872),
            .I(N__47850));
    LocalMux I__11130 (
            .O(N__47869),
            .I(N__47850));
    Span4Mux_v I__11129 (
            .O(N__47866),
            .I(N__47850));
    Span4Mux_v I__11128 (
            .O(N__47863),
            .I(N__47847));
    LocalMux I__11127 (
            .O(N__47860),
            .I(N__47844));
    Span4Mux_v I__11126 (
            .O(N__47857),
            .I(N__47839));
    Span4Mux_h I__11125 (
            .O(N__47850),
            .I(N__47839));
    Odrv4 I__11124 (
            .O(N__47847),
            .I(comm_buf_1_6));
    Odrv12 I__11123 (
            .O(N__47844),
            .I(comm_buf_1_6));
    Odrv4 I__11122 (
            .O(N__47839),
            .I(comm_buf_1_6));
    InMux I__11121 (
            .O(N__47832),
            .I(N__47829));
    LocalMux I__11120 (
            .O(N__47829),
            .I(N__47825));
    InMux I__11119 (
            .O(N__47828),
            .I(N__47822));
    Span4Mux_v I__11118 (
            .O(N__47825),
            .I(N__47819));
    LocalMux I__11117 (
            .O(N__47822),
            .I(N__47816));
    Span4Mux_h I__11116 (
            .O(N__47819),
            .I(N__47813));
    Span4Mux_h I__11115 (
            .O(N__47816),
            .I(N__47810));
    Odrv4 I__11114 (
            .O(N__47813),
            .I(n14_adj_1552));
    Odrv4 I__11113 (
            .O(N__47810),
            .I(n14_adj_1552));
    CascadeMux I__11112 (
            .O(N__47805),
            .I(N__47802));
    InMux I__11111 (
            .O(N__47802),
            .I(N__47798));
    CascadeMux I__11110 (
            .O(N__47801),
            .I(N__47795));
    LocalMux I__11109 (
            .O(N__47798),
            .I(N__47791));
    InMux I__11108 (
            .O(N__47795),
            .I(N__47788));
    InMux I__11107 (
            .O(N__47794),
            .I(N__47785));
    Span4Mux_h I__11106 (
            .O(N__47791),
            .I(N__47778));
    LocalMux I__11105 (
            .O(N__47788),
            .I(N__47778));
    LocalMux I__11104 (
            .O(N__47785),
            .I(N__47775));
    CascadeMux I__11103 (
            .O(N__47784),
            .I(N__47772));
    InMux I__11102 (
            .O(N__47783),
            .I(N__47769));
    Span4Mux_v I__11101 (
            .O(N__47778),
            .I(N__47764));
    Span4Mux_h I__11100 (
            .O(N__47775),
            .I(N__47764));
    InMux I__11099 (
            .O(N__47772),
            .I(N__47760));
    LocalMux I__11098 (
            .O(N__47769),
            .I(N__47757));
    Span4Mux_h I__11097 (
            .O(N__47764),
            .I(N__47754));
    InMux I__11096 (
            .O(N__47763),
            .I(N__47751));
    LocalMux I__11095 (
            .O(N__47760),
            .I(N__47748));
    Span4Mux_h I__11094 (
            .O(N__47757),
            .I(N__47745));
    Span4Mux_h I__11093 (
            .O(N__47754),
            .I(N__47740));
    LocalMux I__11092 (
            .O(N__47751),
            .I(N__47740));
    Span4Mux_h I__11091 (
            .O(N__47748),
            .I(N__47737));
    Span4Mux_v I__11090 (
            .O(N__47745),
            .I(N__47732));
    Span4Mux_v I__11089 (
            .O(N__47740),
            .I(N__47732));
    Odrv4 I__11088 (
            .O(N__47737),
            .I(comm_buf_1_4));
    Odrv4 I__11087 (
            .O(N__47732),
            .I(comm_buf_1_4));
    InMux I__11086 (
            .O(N__47727),
            .I(N__47724));
    LocalMux I__11085 (
            .O(N__47724),
            .I(N__47719));
    InMux I__11084 (
            .O(N__47723),
            .I(N__47716));
    InMux I__11083 (
            .O(N__47722),
            .I(N__47713));
    Span12Mux_s10_h I__11082 (
            .O(N__47719),
            .I(N__47706));
    LocalMux I__11081 (
            .O(N__47716),
            .I(N__47706));
    LocalMux I__11080 (
            .O(N__47713),
            .I(N__47706));
    Odrv12 I__11079 (
            .O(N__47706),
            .I(data_index_4));
    InMux I__11078 (
            .O(N__47703),
            .I(N__47698));
    InMux I__11077 (
            .O(N__47702),
            .I(N__47695));
    InMux I__11076 (
            .O(N__47701),
            .I(N__47692));
    LocalMux I__11075 (
            .O(N__47698),
            .I(N__47684));
    LocalMux I__11074 (
            .O(N__47695),
            .I(N__47684));
    LocalMux I__11073 (
            .O(N__47692),
            .I(N__47677));
    InMux I__11072 (
            .O(N__47691),
            .I(N__47674));
    InMux I__11071 (
            .O(N__47690),
            .I(N__47669));
    InMux I__11070 (
            .O(N__47689),
            .I(N__47669));
    Span4Mux_h I__11069 (
            .O(N__47684),
            .I(N__47666));
    InMux I__11068 (
            .O(N__47683),
            .I(N__47663));
    InMux I__11067 (
            .O(N__47682),
            .I(N__47656));
    InMux I__11066 (
            .O(N__47681),
            .I(N__47656));
    InMux I__11065 (
            .O(N__47680),
            .I(N__47656));
    Span4Mux_v I__11064 (
            .O(N__47677),
            .I(N__47651));
    LocalMux I__11063 (
            .O(N__47674),
            .I(N__47651));
    LocalMux I__11062 (
            .O(N__47669),
            .I(n8813));
    Odrv4 I__11061 (
            .O(N__47666),
            .I(n8813));
    LocalMux I__11060 (
            .O(N__47663),
            .I(n8813));
    LocalMux I__11059 (
            .O(N__47656),
            .I(n8813));
    Odrv4 I__11058 (
            .O(N__47651),
            .I(n8813));
    InMux I__11057 (
            .O(N__47640),
            .I(N__47637));
    LocalMux I__11056 (
            .O(N__47637),
            .I(N__47634));
    Span12Mux_h I__11055 (
            .O(N__47634),
            .I(N__47630));
    InMux I__11054 (
            .O(N__47633),
            .I(N__47627));
    Odrv12 I__11053 (
            .O(N__47630),
            .I(n8_adj_1567));
    LocalMux I__11052 (
            .O(N__47627),
            .I(n8_adj_1567));
    InMux I__11051 (
            .O(N__47622),
            .I(N__47618));
    InMux I__11050 (
            .O(N__47621),
            .I(N__47615));
    LocalMux I__11049 (
            .O(N__47618),
            .I(N__47612));
    LocalMux I__11048 (
            .O(N__47615),
            .I(N__47609));
    Span4Mux_h I__11047 (
            .O(N__47612),
            .I(N__47604));
    Span4Mux_v I__11046 (
            .O(N__47609),
            .I(N__47604));
    Odrv4 I__11045 (
            .O(N__47604),
            .I(n7_adj_1566));
    CascadeMux I__11044 (
            .O(N__47601),
            .I(N__47598));
    CascadeBuf I__11043 (
            .O(N__47598),
            .I(N__47595));
    CascadeMux I__11042 (
            .O(N__47595),
            .I(N__47592));
    CascadeBuf I__11041 (
            .O(N__47592),
            .I(N__47589));
    CascadeMux I__11040 (
            .O(N__47589),
            .I(N__47586));
    CascadeBuf I__11039 (
            .O(N__47586),
            .I(N__47583));
    CascadeMux I__11038 (
            .O(N__47583),
            .I(N__47580));
    CascadeBuf I__11037 (
            .O(N__47580),
            .I(N__47577));
    CascadeMux I__11036 (
            .O(N__47577),
            .I(N__47574));
    CascadeBuf I__11035 (
            .O(N__47574),
            .I(N__47571));
    CascadeMux I__11034 (
            .O(N__47571),
            .I(N__47568));
    CascadeBuf I__11033 (
            .O(N__47568),
            .I(N__47565));
    CascadeMux I__11032 (
            .O(N__47565),
            .I(N__47561));
    CascadeMux I__11031 (
            .O(N__47564),
            .I(N__47558));
    CascadeBuf I__11030 (
            .O(N__47561),
            .I(N__47555));
    CascadeBuf I__11029 (
            .O(N__47558),
            .I(N__47552));
    CascadeMux I__11028 (
            .O(N__47555),
            .I(N__47549));
    CascadeMux I__11027 (
            .O(N__47552),
            .I(N__47546));
    CascadeBuf I__11026 (
            .O(N__47549),
            .I(N__47543));
    InMux I__11025 (
            .O(N__47546),
            .I(N__47540));
    CascadeMux I__11024 (
            .O(N__47543),
            .I(N__47537));
    LocalMux I__11023 (
            .O(N__47540),
            .I(N__47534));
    CascadeBuf I__11022 (
            .O(N__47537),
            .I(N__47531));
    Sp12to4 I__11021 (
            .O(N__47534),
            .I(N__47528));
    CascadeMux I__11020 (
            .O(N__47531),
            .I(N__47525));
    Span12Mux_v I__11019 (
            .O(N__47528),
            .I(N__47522));
    InMux I__11018 (
            .O(N__47525),
            .I(N__47519));
    Span12Mux_h I__11017 (
            .O(N__47522),
            .I(N__47516));
    LocalMux I__11016 (
            .O(N__47519),
            .I(N__47513));
    Odrv12 I__11015 (
            .O(N__47516),
            .I(data_index_9_N_216_4));
    Odrv4 I__11014 (
            .O(N__47513),
            .I(data_index_9_N_216_4));
    CEMux I__11013 (
            .O(N__47508),
            .I(N__47505));
    LocalMux I__11012 (
            .O(N__47505),
            .I(N__47502));
    Span4Mux_h I__11011 (
            .O(N__47502),
            .I(N__47499));
    Span4Mux_h I__11010 (
            .O(N__47499),
            .I(N__47496));
    Odrv4 I__11009 (
            .O(N__47496),
            .I(\ADC_VDC.n11750 ));
    InMux I__11008 (
            .O(N__47493),
            .I(N__47486));
    CascadeMux I__11007 (
            .O(N__47492),
            .I(N__47483));
    CascadeMux I__11006 (
            .O(N__47491),
            .I(N__47477));
    CascadeMux I__11005 (
            .O(N__47490),
            .I(N__47474));
    CascadeMux I__11004 (
            .O(N__47489),
            .I(N__47470));
    LocalMux I__11003 (
            .O(N__47486),
            .I(N__47467));
    InMux I__11002 (
            .O(N__47483),
            .I(N__47464));
    InMux I__11001 (
            .O(N__47482),
            .I(N__47461));
    InMux I__11000 (
            .O(N__47481),
            .I(N__47456));
    InMux I__10999 (
            .O(N__47480),
            .I(N__47456));
    InMux I__10998 (
            .O(N__47477),
            .I(N__47453));
    InMux I__10997 (
            .O(N__47474),
            .I(N__47448));
    InMux I__10996 (
            .O(N__47473),
            .I(N__47448));
    InMux I__10995 (
            .O(N__47470),
            .I(N__47445));
    Span4Mux_v I__10994 (
            .O(N__47467),
            .I(N__47442));
    LocalMux I__10993 (
            .O(N__47464),
            .I(N__47439));
    LocalMux I__10992 (
            .O(N__47461),
            .I(N__47436));
    LocalMux I__10991 (
            .O(N__47456),
            .I(N__47427));
    LocalMux I__10990 (
            .O(N__47453),
            .I(N__47427));
    LocalMux I__10989 (
            .O(N__47448),
            .I(N__47427));
    LocalMux I__10988 (
            .O(N__47445),
            .I(N__47427));
    Span4Mux_h I__10987 (
            .O(N__47442),
            .I(N__47419));
    Span4Mux_v I__10986 (
            .O(N__47439),
            .I(N__47419));
    Span4Mux_v I__10985 (
            .O(N__47436),
            .I(N__47419));
    Span4Mux_v I__10984 (
            .O(N__47427),
            .I(N__47416));
    CascadeMux I__10983 (
            .O(N__47426),
            .I(N__47413));
    Span4Mux_v I__10982 (
            .O(N__47419),
            .I(N__47410));
    Span4Mux_v I__10981 (
            .O(N__47416),
            .I(N__47407));
    InMux I__10980 (
            .O(N__47413),
            .I(N__47404));
    Sp12to4 I__10979 (
            .O(N__47410),
            .I(N__47401));
    Span4Mux_h I__10978 (
            .O(N__47407),
            .I(N__47398));
    LocalMux I__10977 (
            .O(N__47404),
            .I(N__47395));
    Span12Mux_h I__10976 (
            .O(N__47401),
            .I(N__47388));
    Sp12to4 I__10975 (
            .O(N__47398),
            .I(N__47388));
    Span12Mux_v I__10974 (
            .O(N__47395),
            .I(N__47388));
    Odrv12 I__10973 (
            .O(N__47388),
            .I(VDC_SDO));
    InMux I__10972 (
            .O(N__47385),
            .I(N__47378));
    InMux I__10971 (
            .O(N__47384),
            .I(N__47378));
    InMux I__10970 (
            .O(N__47383),
            .I(N__47374));
    LocalMux I__10969 (
            .O(N__47378),
            .I(N__47371));
    InMux I__10968 (
            .O(N__47377),
            .I(N__47368));
    LocalMux I__10967 (
            .O(N__47374),
            .I(N__47352));
    Span4Mux_v I__10966 (
            .O(N__47371),
            .I(N__47352));
    LocalMux I__10965 (
            .O(N__47368),
            .I(N__47349));
    InMux I__10964 (
            .O(N__47367),
            .I(N__47344));
    InMux I__10963 (
            .O(N__47366),
            .I(N__47341));
    InMux I__10962 (
            .O(N__47365),
            .I(N__47336));
    InMux I__10961 (
            .O(N__47364),
            .I(N__47336));
    InMux I__10960 (
            .O(N__47363),
            .I(N__47329));
    InMux I__10959 (
            .O(N__47362),
            .I(N__47322));
    InMux I__10958 (
            .O(N__47361),
            .I(N__47322));
    InMux I__10957 (
            .O(N__47360),
            .I(N__47322));
    InMux I__10956 (
            .O(N__47359),
            .I(N__47317));
    InMux I__10955 (
            .O(N__47358),
            .I(N__47317));
    InMux I__10954 (
            .O(N__47357),
            .I(N__47314));
    Span4Mux_h I__10953 (
            .O(N__47352),
            .I(N__47309));
    Span4Mux_h I__10952 (
            .O(N__47349),
            .I(N__47309));
    InMux I__10951 (
            .O(N__47348),
            .I(N__47304));
    InMux I__10950 (
            .O(N__47347),
            .I(N__47304));
    LocalMux I__10949 (
            .O(N__47344),
            .I(N__47297));
    LocalMux I__10948 (
            .O(N__47341),
            .I(N__47297));
    LocalMux I__10947 (
            .O(N__47336),
            .I(N__47297));
    InMux I__10946 (
            .O(N__47335),
            .I(N__47290));
    InMux I__10945 (
            .O(N__47334),
            .I(N__47290));
    InMux I__10944 (
            .O(N__47333),
            .I(N__47290));
    InMux I__10943 (
            .O(N__47332),
            .I(N__47287));
    LocalMux I__10942 (
            .O(N__47329),
            .I(N__47284));
    LocalMux I__10941 (
            .O(N__47322),
            .I(N__47279));
    LocalMux I__10940 (
            .O(N__47317),
            .I(N__47279));
    LocalMux I__10939 (
            .O(N__47314),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__10938 (
            .O(N__47309),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__10937 (
            .O(N__47304),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv12 I__10936 (
            .O(N__47297),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__10935 (
            .O(N__47290),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__10934 (
            .O(N__47287),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv12 I__10933 (
            .O(N__47284),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__10932 (
            .O(N__47279),
            .I(\ADC_VDC.adc_state_0 ));
    CascadeMux I__10931 (
            .O(N__47262),
            .I(N__47259));
    InMux I__10930 (
            .O(N__47259),
            .I(N__47256));
    LocalMux I__10929 (
            .O(N__47256),
            .I(\ADC_VDC.n62 ));
    InMux I__10928 (
            .O(N__47253),
            .I(N__47250));
    LocalMux I__10927 (
            .O(N__47250),
            .I(n22210));
    CascadeMux I__10926 (
            .O(N__47247),
            .I(n22432_cascade_));
    InMux I__10925 (
            .O(N__47244),
            .I(N__47240));
    InMux I__10924 (
            .O(N__47243),
            .I(N__47237));
    LocalMux I__10923 (
            .O(N__47240),
            .I(N__47233));
    LocalMux I__10922 (
            .O(N__47237),
            .I(N__47228));
    InMux I__10921 (
            .O(N__47236),
            .I(N__47225));
    Span4Mux_v I__10920 (
            .O(N__47233),
            .I(N__47220));
    InMux I__10919 (
            .O(N__47232),
            .I(N__47217));
    InMux I__10918 (
            .O(N__47231),
            .I(N__47214));
    Span4Mux_v I__10917 (
            .O(N__47228),
            .I(N__47209));
    LocalMux I__10916 (
            .O(N__47225),
            .I(N__47209));
    CascadeMux I__10915 (
            .O(N__47224),
            .I(N__47206));
    CascadeMux I__10914 (
            .O(N__47223),
            .I(N__47203));
    Span4Mux_h I__10913 (
            .O(N__47220),
            .I(N__47196));
    LocalMux I__10912 (
            .O(N__47217),
            .I(N__47196));
    LocalMux I__10911 (
            .O(N__47214),
            .I(N__47196));
    Span4Mux_v I__10910 (
            .O(N__47209),
            .I(N__47193));
    InMux I__10909 (
            .O(N__47206),
            .I(N__47190));
    InMux I__10908 (
            .O(N__47203),
            .I(N__47187));
    Span4Mux_v I__10907 (
            .O(N__47196),
            .I(N__47184));
    Span4Mux_h I__10906 (
            .O(N__47193),
            .I(N__47179));
    LocalMux I__10905 (
            .O(N__47190),
            .I(N__47179));
    LocalMux I__10904 (
            .O(N__47187),
            .I(N__47176));
    Sp12to4 I__10903 (
            .O(N__47184),
            .I(N__47171));
    Span4Mux_v I__10902 (
            .O(N__47179),
            .I(N__47166));
    Span4Mux_v I__10901 (
            .O(N__47176),
            .I(N__47166));
    InMux I__10900 (
            .O(N__47175),
            .I(N__47163));
    InMux I__10899 (
            .O(N__47174),
            .I(N__47160));
    Odrv12 I__10898 (
            .O(N__47171),
            .I(comm_rx_buf_2));
    Odrv4 I__10897 (
            .O(N__47166),
            .I(comm_rx_buf_2));
    LocalMux I__10896 (
            .O(N__47163),
            .I(comm_rx_buf_2));
    LocalMux I__10895 (
            .O(N__47160),
            .I(comm_rx_buf_2));
    CascadeMux I__10894 (
            .O(N__47151),
            .I(n30_adj_1520_cascade_));
    InMux I__10893 (
            .O(N__47148),
            .I(N__47144));
    CascadeMux I__10892 (
            .O(N__47147),
            .I(N__47141));
    LocalMux I__10891 (
            .O(N__47144),
            .I(N__47138));
    InMux I__10890 (
            .O(N__47141),
            .I(N__47135));
    Span4Mux_h I__10889 (
            .O(N__47138),
            .I(N__47132));
    LocalMux I__10888 (
            .O(N__47135),
            .I(data_idxvec_2));
    Odrv4 I__10887 (
            .O(N__47132),
            .I(data_idxvec_2));
    InMux I__10886 (
            .O(N__47127),
            .I(N__47124));
    LocalMux I__10885 (
            .O(N__47124),
            .I(N__47119));
    InMux I__10884 (
            .O(N__47123),
            .I(N__47116));
    InMux I__10883 (
            .O(N__47122),
            .I(N__47113));
    Span4Mux_h I__10882 (
            .O(N__47119),
            .I(N__47110));
    LocalMux I__10881 (
            .O(N__47116),
            .I(data_cntvec_2));
    LocalMux I__10880 (
            .O(N__47113),
            .I(data_cntvec_2));
    Odrv4 I__10879 (
            .O(N__47110),
            .I(data_cntvec_2));
    InMux I__10878 (
            .O(N__47103),
            .I(N__47100));
    LocalMux I__10877 (
            .O(N__47100),
            .I(n26_adj_1519));
    InMux I__10876 (
            .O(N__47097),
            .I(N__47093));
    InMux I__10875 (
            .O(N__47096),
            .I(N__47089));
    LocalMux I__10874 (
            .O(N__47093),
            .I(N__47086));
    InMux I__10873 (
            .O(N__47092),
            .I(N__47083));
    LocalMux I__10872 (
            .O(N__47089),
            .I(N__47080));
    Span4Mux_v I__10871 (
            .O(N__47086),
            .I(N__47077));
    LocalMux I__10870 (
            .O(N__47083),
            .I(N__47074));
    Span4Mux_h I__10869 (
            .O(N__47080),
            .I(N__47071));
    Span4Mux_h I__10868 (
            .O(N__47077),
            .I(N__47068));
    Span4Mux_v I__10867 (
            .O(N__47074),
            .I(N__47063));
    Span4Mux_h I__10866 (
            .O(N__47071),
            .I(N__47063));
    Odrv4 I__10865 (
            .O(N__47068),
            .I(n14_adj_1585));
    Odrv4 I__10864 (
            .O(N__47063),
            .I(n14_adj_1585));
    InMux I__10863 (
            .O(N__47058),
            .I(N__47055));
    LocalMux I__10862 (
            .O(N__47055),
            .I(N__47052));
    Span4Mux_h I__10861 (
            .O(N__47052),
            .I(N__47049));
    Odrv4 I__10860 (
            .O(N__47049),
            .I(n8));
    InMux I__10859 (
            .O(N__47046),
            .I(N__47043));
    LocalMux I__10858 (
            .O(N__47043),
            .I(N__47040));
    Span4Mux_v I__10857 (
            .O(N__47040),
            .I(N__47036));
    InMux I__10856 (
            .O(N__47039),
            .I(N__47033));
    Sp12to4 I__10855 (
            .O(N__47036),
            .I(N__47027));
    LocalMux I__10854 (
            .O(N__47033),
            .I(N__47027));
    InMux I__10853 (
            .O(N__47032),
            .I(N__47024));
    Span12Mux_h I__10852 (
            .O(N__47027),
            .I(N__47021));
    LocalMux I__10851 (
            .O(N__47024),
            .I(buf_adcdata_iac_14));
    Odrv12 I__10850 (
            .O(N__47021),
            .I(buf_adcdata_iac_14));
    InMux I__10849 (
            .O(N__47016),
            .I(N__47013));
    LocalMux I__10848 (
            .O(N__47013),
            .I(N__47010));
    Odrv4 I__10847 (
            .O(N__47010),
            .I(n16));
    InMux I__10846 (
            .O(N__47007),
            .I(N__47004));
    LocalMux I__10845 (
            .O(N__47004),
            .I(N__47001));
    Odrv4 I__10844 (
            .O(N__47001),
            .I(n21045));
    InMux I__10843 (
            .O(N__46998),
            .I(N__46994));
    CascadeMux I__10842 (
            .O(N__46997),
            .I(N__46990));
    LocalMux I__10841 (
            .O(N__46994),
            .I(N__46987));
    InMux I__10840 (
            .O(N__46993),
            .I(N__46982));
    InMux I__10839 (
            .O(N__46990),
            .I(N__46982));
    Odrv12 I__10838 (
            .O(N__46987),
            .I(req_data_cnt_7));
    LocalMux I__10837 (
            .O(N__46982),
            .I(req_data_cnt_7));
    InMux I__10836 (
            .O(N__46977),
            .I(N__46973));
    InMux I__10835 (
            .O(N__46976),
            .I(N__46969));
    LocalMux I__10834 (
            .O(N__46973),
            .I(N__46966));
    InMux I__10833 (
            .O(N__46972),
            .I(N__46963));
    LocalMux I__10832 (
            .O(N__46969),
            .I(acadc_skipCount_7));
    Odrv4 I__10831 (
            .O(N__46966),
            .I(acadc_skipCount_7));
    LocalMux I__10830 (
            .O(N__46963),
            .I(acadc_skipCount_7));
    InMux I__10829 (
            .O(N__46956),
            .I(N__46953));
    LocalMux I__10828 (
            .O(N__46953),
            .I(N__46949));
    CascadeMux I__10827 (
            .O(N__46952),
            .I(N__46946));
    Sp12to4 I__10826 (
            .O(N__46949),
            .I(N__46942));
    InMux I__10825 (
            .O(N__46946),
            .I(N__46939));
    InMux I__10824 (
            .O(N__46945),
            .I(N__46936));
    Span12Mux_v I__10823 (
            .O(N__46942),
            .I(N__46933));
    LocalMux I__10822 (
            .O(N__46939),
            .I(N__46930));
    LocalMux I__10821 (
            .O(N__46936),
            .I(buf_dds1_3));
    Odrv12 I__10820 (
            .O(N__46933),
            .I(buf_dds1_3));
    Odrv4 I__10819 (
            .O(N__46930),
            .I(buf_dds1_3));
    InMux I__10818 (
            .O(N__46923),
            .I(N__46920));
    LocalMux I__10817 (
            .O(N__46920),
            .I(N__46917));
    Span4Mux_h I__10816 (
            .O(N__46917),
            .I(N__46912));
    InMux I__10815 (
            .O(N__46916),
            .I(N__46909));
    InMux I__10814 (
            .O(N__46915),
            .I(N__46906));
    Span4Mux_h I__10813 (
            .O(N__46912),
            .I(N__46903));
    LocalMux I__10812 (
            .O(N__46909),
            .I(N__46900));
    LocalMux I__10811 (
            .O(N__46906),
            .I(buf_dds0_3));
    Odrv4 I__10810 (
            .O(N__46903),
            .I(buf_dds0_3));
    Odrv4 I__10809 (
            .O(N__46900),
            .I(buf_dds0_3));
    InMux I__10808 (
            .O(N__46893),
            .I(N__46888));
    InMux I__10807 (
            .O(N__46892),
            .I(N__46885));
    CascadeMux I__10806 (
            .O(N__46891),
            .I(N__46882));
    LocalMux I__10805 (
            .O(N__46888),
            .I(N__46879));
    LocalMux I__10804 (
            .O(N__46885),
            .I(N__46876));
    InMux I__10803 (
            .O(N__46882),
            .I(N__46873));
    Span4Mux_h I__10802 (
            .O(N__46879),
            .I(N__46868));
    Span4Mux_v I__10801 (
            .O(N__46876),
            .I(N__46868));
    LocalMux I__10800 (
            .O(N__46873),
            .I(buf_dds1_2));
    Odrv4 I__10799 (
            .O(N__46868),
            .I(buf_dds1_2));
    InMux I__10798 (
            .O(N__46863),
            .I(N__46860));
    LocalMux I__10797 (
            .O(N__46860),
            .I(N__46857));
    Odrv4 I__10796 (
            .O(N__46857),
            .I(n16_adj_1517));
    CascadeMux I__10795 (
            .O(N__46854),
            .I(n26_adj_1512_cascade_));
    InMux I__10794 (
            .O(N__46851),
            .I(N__46848));
    LocalMux I__10793 (
            .O(N__46848),
            .I(N__46845));
    Span4Mux_h I__10792 (
            .O(N__46845),
            .I(N__46842));
    Span4Mux_v I__10791 (
            .O(N__46842),
            .I(N__46839));
    Span4Mux_h I__10790 (
            .O(N__46839),
            .I(N__46834));
    InMux I__10789 (
            .O(N__46838),
            .I(N__46829));
    InMux I__10788 (
            .O(N__46837),
            .I(N__46829));
    Odrv4 I__10787 (
            .O(N__46834),
            .I(acadc_skipCount_4));
    LocalMux I__10786 (
            .O(N__46829),
            .I(acadc_skipCount_4));
    CascadeMux I__10785 (
            .O(N__46824),
            .I(n22351_cascade_));
    InMux I__10784 (
            .O(N__46821),
            .I(N__46818));
    LocalMux I__10783 (
            .O(N__46818),
            .I(N__46814));
    CascadeMux I__10782 (
            .O(N__46817),
            .I(N__46810));
    Span4Mux_v I__10781 (
            .O(N__46814),
            .I(N__46807));
    InMux I__10780 (
            .O(N__46813),
            .I(N__46802));
    InMux I__10779 (
            .O(N__46810),
            .I(N__46802));
    Odrv4 I__10778 (
            .O(N__46807),
            .I(req_data_cnt_4));
    LocalMux I__10777 (
            .O(N__46802),
            .I(req_data_cnt_4));
    InMux I__10776 (
            .O(N__46797),
            .I(N__46794));
    LocalMux I__10775 (
            .O(N__46794),
            .I(n22234));
    CascadeMux I__10774 (
            .O(N__46791),
            .I(n22354_cascade_));
    InMux I__10773 (
            .O(N__46788),
            .I(N__46783));
    InMux I__10772 (
            .O(N__46787),
            .I(N__46780));
    InMux I__10771 (
            .O(N__46786),
            .I(N__46777));
    LocalMux I__10770 (
            .O(N__46783),
            .I(N__46773));
    LocalMux I__10769 (
            .O(N__46780),
            .I(N__46769));
    LocalMux I__10768 (
            .O(N__46777),
            .I(N__46766));
    InMux I__10767 (
            .O(N__46776),
            .I(N__46763));
    Span4Mux_h I__10766 (
            .O(N__46773),
            .I(N__46759));
    InMux I__10765 (
            .O(N__46772),
            .I(N__46756));
    Span4Mux_v I__10764 (
            .O(N__46769),
            .I(N__46748));
    Span4Mux_h I__10763 (
            .O(N__46766),
            .I(N__46748));
    LocalMux I__10762 (
            .O(N__46763),
            .I(N__46748));
    InMux I__10761 (
            .O(N__46762),
            .I(N__46745));
    Span4Mux_v I__10760 (
            .O(N__46759),
            .I(N__46740));
    LocalMux I__10759 (
            .O(N__46756),
            .I(N__46740));
    CascadeMux I__10758 (
            .O(N__46755),
            .I(N__46737));
    Span4Mux_v I__10757 (
            .O(N__46748),
            .I(N__46734));
    LocalMux I__10756 (
            .O(N__46745),
            .I(N__46731));
    Span4Mux_h I__10755 (
            .O(N__46740),
            .I(N__46727));
    InMux I__10754 (
            .O(N__46737),
            .I(N__46724));
    Span4Mux_h I__10753 (
            .O(N__46734),
            .I(N__46719));
    Span4Mux_h I__10752 (
            .O(N__46731),
            .I(N__46719));
    InMux I__10751 (
            .O(N__46730),
            .I(N__46716));
    Span4Mux_h I__10750 (
            .O(N__46727),
            .I(N__46712));
    LocalMux I__10749 (
            .O(N__46724),
            .I(N__46709));
    Sp12to4 I__10748 (
            .O(N__46719),
            .I(N__46706));
    LocalMux I__10747 (
            .O(N__46716),
            .I(N__46703));
    InMux I__10746 (
            .O(N__46715),
            .I(N__46700));
    Odrv4 I__10745 (
            .O(N__46712),
            .I(comm_rx_buf_4));
    Odrv4 I__10744 (
            .O(N__46709),
            .I(comm_rx_buf_4));
    Odrv12 I__10743 (
            .O(N__46706),
            .I(comm_rx_buf_4));
    Odrv4 I__10742 (
            .O(N__46703),
            .I(comm_rx_buf_4));
    LocalMux I__10741 (
            .O(N__46700),
            .I(comm_rx_buf_4));
    CascadeMux I__10740 (
            .O(N__46689),
            .I(n30_adj_1513_cascade_));
    InMux I__10739 (
            .O(N__46686),
            .I(N__46683));
    LocalMux I__10738 (
            .O(N__46683),
            .I(N__46680));
    Span4Mux_h I__10737 (
            .O(N__46680),
            .I(N__46677));
    Odrv4 I__10736 (
            .O(N__46677),
            .I(n19_adj_1518));
    CascadeMux I__10735 (
            .O(N__46674),
            .I(N__46671));
    InMux I__10734 (
            .O(N__46671),
            .I(N__46668));
    LocalMux I__10733 (
            .O(N__46668),
            .I(N__46665));
    Span12Mux_h I__10732 (
            .O(N__46665),
            .I(N__46661));
    CascadeMux I__10731 (
            .O(N__46664),
            .I(N__46658));
    Span12Mux_h I__10730 (
            .O(N__46661),
            .I(N__46655));
    InMux I__10729 (
            .O(N__46658),
            .I(N__46652));
    Odrv12 I__10728 (
            .O(N__46655),
            .I(buf_readRTD_2));
    LocalMux I__10727 (
            .O(N__46652),
            .I(buf_readRTD_2));
    InMux I__10726 (
            .O(N__46647),
            .I(N__46644));
    LocalMux I__10725 (
            .O(N__46644),
            .I(N__46641));
    Span4Mux_v I__10724 (
            .O(N__46641),
            .I(N__46637));
    InMux I__10723 (
            .O(N__46640),
            .I(N__46634));
    Sp12to4 I__10722 (
            .O(N__46637),
            .I(N__46628));
    LocalMux I__10721 (
            .O(N__46634),
            .I(N__46628));
    InMux I__10720 (
            .O(N__46633),
            .I(N__46625));
    Span12Mux_h I__10719 (
            .O(N__46628),
            .I(N__46622));
    LocalMux I__10718 (
            .O(N__46625),
            .I(buf_adcdata_iac_10));
    Odrv12 I__10717 (
            .O(N__46622),
            .I(buf_adcdata_iac_10));
    CascadeMux I__10716 (
            .O(N__46617),
            .I(n22207_cascade_));
    InMux I__10715 (
            .O(N__46614),
            .I(N__46611));
    LocalMux I__10714 (
            .O(N__46611),
            .I(N__46608));
    Span4Mux_v I__10713 (
            .O(N__46608),
            .I(N__46604));
    InMux I__10712 (
            .O(N__46607),
            .I(N__46600));
    Span4Mux_h I__10711 (
            .O(N__46604),
            .I(N__46597));
    InMux I__10710 (
            .O(N__46603),
            .I(N__46594));
    LocalMux I__10709 (
            .O(N__46600),
            .I(req_data_cnt_2));
    Odrv4 I__10708 (
            .O(N__46597),
            .I(req_data_cnt_2));
    LocalMux I__10707 (
            .O(N__46594),
            .I(req_data_cnt_2));
    CascadeMux I__10706 (
            .O(N__46587),
            .I(n22429_cascade_));
    InMux I__10705 (
            .O(N__46584),
            .I(N__46581));
    LocalMux I__10704 (
            .O(N__46581),
            .I(N__46576));
    CascadeMux I__10703 (
            .O(N__46580),
            .I(N__46573));
    InMux I__10702 (
            .O(N__46579),
            .I(N__46570));
    Span4Mux_h I__10701 (
            .O(N__46576),
            .I(N__46567));
    InMux I__10700 (
            .O(N__46573),
            .I(N__46564));
    LocalMux I__10699 (
            .O(N__46570),
            .I(acadc_skipCount_2));
    Odrv4 I__10698 (
            .O(N__46567),
            .I(acadc_skipCount_2));
    LocalMux I__10697 (
            .O(N__46564),
            .I(acadc_skipCount_2));
    CascadeMux I__10696 (
            .O(N__46557),
            .I(N__46554));
    InMux I__10695 (
            .O(N__46554),
            .I(N__46551));
    LocalMux I__10694 (
            .O(N__46551),
            .I(N__46548));
    Span4Mux_v I__10693 (
            .O(N__46548),
            .I(N__46545));
    Span4Mux_h I__10692 (
            .O(N__46545),
            .I(N__46542));
    Odrv4 I__10691 (
            .O(N__46542),
            .I(n21177));
    CascadeMux I__10690 (
            .O(N__46539),
            .I(n22225_cascade_));
    InMux I__10689 (
            .O(N__46536),
            .I(N__46532));
    CascadeMux I__10688 (
            .O(N__46535),
            .I(N__46529));
    LocalMux I__10687 (
            .O(N__46532),
            .I(N__46526));
    InMux I__10686 (
            .O(N__46529),
            .I(N__46523));
    Span4Mux_h I__10685 (
            .O(N__46526),
            .I(N__46520));
    LocalMux I__10684 (
            .O(N__46523),
            .I(data_idxvec_6));
    Odrv4 I__10683 (
            .O(N__46520),
            .I(data_idxvec_6));
    InMux I__10682 (
            .O(N__46515),
            .I(N__46512));
    LocalMux I__10681 (
            .O(N__46512),
            .I(N__46508));
    InMux I__10680 (
            .O(N__46511),
            .I(N__46504));
    Span4Mux_v I__10679 (
            .O(N__46508),
            .I(N__46501));
    InMux I__10678 (
            .O(N__46507),
            .I(N__46498));
    LocalMux I__10677 (
            .O(N__46504),
            .I(N__46495));
    Span4Mux_h I__10676 (
            .O(N__46501),
            .I(N__46492));
    LocalMux I__10675 (
            .O(N__46498),
            .I(data_cntvec_6));
    Odrv4 I__10674 (
            .O(N__46495),
            .I(data_cntvec_6));
    Odrv4 I__10673 (
            .O(N__46492),
            .I(data_cntvec_6));
    InMux I__10672 (
            .O(N__46485),
            .I(N__46482));
    LocalMux I__10671 (
            .O(N__46482),
            .I(N__46479));
    Span12Mux_h I__10670 (
            .O(N__46479),
            .I(N__46476));
    Odrv12 I__10669 (
            .O(N__46476),
            .I(buf_data_iac_14));
    CascadeMux I__10668 (
            .O(N__46473),
            .I(n26_adj_1507_cascade_));
    InMux I__10667 (
            .O(N__46470),
            .I(N__46467));
    LocalMux I__10666 (
            .O(N__46467),
            .I(n21178));
    CascadeMux I__10665 (
            .O(N__46464),
            .I(N__46458));
    InMux I__10664 (
            .O(N__46463),
            .I(N__46455));
    InMux I__10663 (
            .O(N__46462),
            .I(N__46452));
    InMux I__10662 (
            .O(N__46461),
            .I(N__46449));
    InMux I__10661 (
            .O(N__46458),
            .I(N__46443));
    LocalMux I__10660 (
            .O(N__46455),
            .I(N__46436));
    LocalMux I__10659 (
            .O(N__46452),
            .I(N__46436));
    LocalMux I__10658 (
            .O(N__46449),
            .I(N__46436));
    CascadeMux I__10657 (
            .O(N__46448),
            .I(N__46433));
    InMux I__10656 (
            .O(N__46447),
            .I(N__46430));
    InMux I__10655 (
            .O(N__46446),
            .I(N__46427));
    LocalMux I__10654 (
            .O(N__46443),
            .I(N__46424));
    Span4Mux_v I__10653 (
            .O(N__46436),
            .I(N__46421));
    InMux I__10652 (
            .O(N__46433),
            .I(N__46418));
    LocalMux I__10651 (
            .O(N__46430),
            .I(N__46413));
    LocalMux I__10650 (
            .O(N__46427),
            .I(N__46413));
    Span4Mux_v I__10649 (
            .O(N__46424),
            .I(N__46406));
    Span4Mux_h I__10648 (
            .O(N__46421),
            .I(N__46406));
    LocalMux I__10647 (
            .O(N__46418),
            .I(N__46406));
    Span4Mux_v I__10646 (
            .O(N__46413),
            .I(N__46401));
    Span4Mux_v I__10645 (
            .O(N__46406),
            .I(N__46398));
    InMux I__10644 (
            .O(N__46405),
            .I(N__46395));
    InMux I__10643 (
            .O(N__46404),
            .I(N__46392));
    Odrv4 I__10642 (
            .O(N__46401),
            .I(comm_rx_buf_6));
    Odrv4 I__10641 (
            .O(N__46398),
            .I(comm_rx_buf_6));
    LocalMux I__10640 (
            .O(N__46395),
            .I(comm_rx_buf_6));
    LocalMux I__10639 (
            .O(N__46392),
            .I(comm_rx_buf_6));
    InMux I__10638 (
            .O(N__46383),
            .I(N__46380));
    LocalMux I__10637 (
            .O(N__46380),
            .I(n22228));
    InMux I__10636 (
            .O(N__46377),
            .I(N__46374));
    LocalMux I__10635 (
            .O(N__46374),
            .I(N__46371));
    Span4Mux_h I__10634 (
            .O(N__46371),
            .I(N__46368));
    Span4Mux_h I__10633 (
            .O(N__46368),
            .I(N__46365));
    Span4Mux_v I__10632 (
            .O(N__46365),
            .I(N__46361));
    InMux I__10631 (
            .O(N__46364),
            .I(N__46358));
    Odrv4 I__10630 (
            .O(N__46361),
            .I(buf_adcdata_vdc_14));
    LocalMux I__10629 (
            .O(N__46358),
            .I(buf_adcdata_vdc_14));
    InMux I__10628 (
            .O(N__46353),
            .I(N__46350));
    LocalMux I__10627 (
            .O(N__46350),
            .I(N__46346));
    InMux I__10626 (
            .O(N__46349),
            .I(N__46343));
    Span12Mux_v I__10625 (
            .O(N__46346),
            .I(N__46339));
    LocalMux I__10624 (
            .O(N__46343),
            .I(N__46336));
    InMux I__10623 (
            .O(N__46342),
            .I(N__46333));
    Span12Mux_h I__10622 (
            .O(N__46339),
            .I(N__46330));
    Span12Mux_s10_h I__10621 (
            .O(N__46336),
            .I(N__46327));
    LocalMux I__10620 (
            .O(N__46333),
            .I(buf_adcdata_vac_14));
    Odrv12 I__10619 (
            .O(N__46330),
            .I(buf_adcdata_vac_14));
    Odrv12 I__10618 (
            .O(N__46327),
            .I(buf_adcdata_vac_14));
    CascadeMux I__10617 (
            .O(N__46320),
            .I(n19_cascade_));
    InMux I__10616 (
            .O(N__46317),
            .I(N__46314));
    LocalMux I__10615 (
            .O(N__46314),
            .I(N__46311));
    Span4Mux_v I__10614 (
            .O(N__46311),
            .I(N__46308));
    Span4Mux_h I__10613 (
            .O(N__46308),
            .I(N__46305));
    Span4Mux_h I__10612 (
            .O(N__46305),
            .I(N__46301));
    CascadeMux I__10611 (
            .O(N__46304),
            .I(N__46298));
    Span4Mux_h I__10610 (
            .O(N__46301),
            .I(N__46295));
    InMux I__10609 (
            .O(N__46298),
            .I(N__46292));
    Odrv4 I__10608 (
            .O(N__46295),
            .I(buf_readRTD_6));
    LocalMux I__10607 (
            .O(N__46292),
            .I(buf_readRTD_6));
    InMux I__10606 (
            .O(N__46287),
            .I(N__46284));
    LocalMux I__10605 (
            .O(N__46284),
            .I(n21046));
    InMux I__10604 (
            .O(N__46281),
            .I(N__46278));
    LocalMux I__10603 (
            .O(N__46278),
            .I(N__46275));
    Sp12to4 I__10602 (
            .O(N__46275),
            .I(N__46272));
    Odrv12 I__10601 (
            .O(N__46272),
            .I(n16_adj_1510));
    CascadeMux I__10600 (
            .O(N__46269),
            .I(N__46265));
    InMux I__10599 (
            .O(N__46268),
            .I(N__46262));
    InMux I__10598 (
            .O(N__46265),
            .I(N__46259));
    LocalMux I__10597 (
            .O(N__46262),
            .I(N__46256));
    LocalMux I__10596 (
            .O(N__46259),
            .I(N__46252));
    Span12Mux_v I__10595 (
            .O(N__46256),
            .I(N__46249));
    InMux I__10594 (
            .O(N__46255),
            .I(N__46246));
    Span4Mux_h I__10593 (
            .O(N__46252),
            .I(N__46243));
    Span12Mux_h I__10592 (
            .O(N__46249),
            .I(N__46240));
    LocalMux I__10591 (
            .O(N__46246),
            .I(N__46235));
    Span4Mux_h I__10590 (
            .O(N__46243),
            .I(N__46235));
    Odrv12 I__10589 (
            .O(N__46240),
            .I(buf_adcdata_iac_12));
    Odrv4 I__10588 (
            .O(N__46235),
            .I(buf_adcdata_iac_12));
    InMux I__10587 (
            .O(N__46230),
            .I(N__46227));
    LocalMux I__10586 (
            .O(N__46227),
            .I(N__46224));
    Sp12to4 I__10585 (
            .O(N__46224),
            .I(N__46221));
    Odrv12 I__10584 (
            .O(N__46221),
            .I(n22231));
    InMux I__10583 (
            .O(N__46218),
            .I(N__46214));
    CascadeMux I__10582 (
            .O(N__46217),
            .I(N__46211));
    LocalMux I__10581 (
            .O(N__46214),
            .I(N__46208));
    InMux I__10580 (
            .O(N__46211),
            .I(N__46205));
    Span4Mux_h I__10579 (
            .O(N__46208),
            .I(N__46202));
    LocalMux I__10578 (
            .O(N__46205),
            .I(data_idxvec_4));
    Odrv4 I__10577 (
            .O(N__46202),
            .I(data_idxvec_4));
    InMux I__10576 (
            .O(N__46197),
            .I(N__46194));
    LocalMux I__10575 (
            .O(N__46194),
            .I(N__46189));
    InMux I__10574 (
            .O(N__46193),
            .I(N__46186));
    InMux I__10573 (
            .O(N__46192),
            .I(N__46183));
    Span4Mux_v I__10572 (
            .O(N__46189),
            .I(N__46180));
    LocalMux I__10571 (
            .O(N__46186),
            .I(data_cntvec_4));
    LocalMux I__10570 (
            .O(N__46183),
            .I(data_cntvec_4));
    Odrv4 I__10569 (
            .O(N__46180),
            .I(data_cntvec_4));
    CEMux I__10568 (
            .O(N__46173),
            .I(N__46170));
    LocalMux I__10567 (
            .O(N__46170),
            .I(N__46161));
    CEMux I__10566 (
            .O(N__46169),
            .I(N__46158));
    CEMux I__10565 (
            .O(N__46168),
            .I(N__46155));
    CEMux I__10564 (
            .O(N__46167),
            .I(N__46152));
    CEMux I__10563 (
            .O(N__46166),
            .I(N__46149));
    CEMux I__10562 (
            .O(N__46165),
            .I(N__46146));
    CEMux I__10561 (
            .O(N__46164),
            .I(N__46143));
    Span4Mux_v I__10560 (
            .O(N__46161),
            .I(N__46138));
    LocalMux I__10559 (
            .O(N__46158),
            .I(N__46138));
    LocalMux I__10558 (
            .O(N__46155),
            .I(N__46135));
    LocalMux I__10557 (
            .O(N__46152),
            .I(N__46132));
    LocalMux I__10556 (
            .O(N__46149),
            .I(N__46127));
    LocalMux I__10555 (
            .O(N__46146),
            .I(N__46127));
    LocalMux I__10554 (
            .O(N__46143),
            .I(N__46124));
    Span4Mux_v I__10553 (
            .O(N__46138),
            .I(N__46120));
    Span4Mux_h I__10552 (
            .O(N__46135),
            .I(N__46117));
    Span4Mux_h I__10551 (
            .O(N__46132),
            .I(N__46114));
    Span4Mux_v I__10550 (
            .O(N__46127),
            .I(N__46109));
    Span4Mux_h I__10549 (
            .O(N__46124),
            .I(N__46109));
    InMux I__10548 (
            .O(N__46123),
            .I(N__46106));
    Odrv4 I__10547 (
            .O(N__46120),
            .I(n11961));
    Odrv4 I__10546 (
            .O(N__46117),
            .I(n11961));
    Odrv4 I__10545 (
            .O(N__46114),
            .I(n11961));
    Odrv4 I__10544 (
            .O(N__46109),
            .I(n11961));
    LocalMux I__10543 (
            .O(N__46106),
            .I(n11961));
    CascadeMux I__10542 (
            .O(N__46095),
            .I(n18993_cascade_));
    InMux I__10541 (
            .O(N__46092),
            .I(N__46089));
    LocalMux I__10540 (
            .O(N__46089),
            .I(n12_adj_1605));
    CascadeMux I__10539 (
            .O(N__46086),
            .I(n11991_cascade_));
    InMux I__10538 (
            .O(N__46083),
            .I(N__46075));
    CascadeMux I__10537 (
            .O(N__46082),
            .I(N__46072));
    InMux I__10536 (
            .O(N__46081),
            .I(N__46067));
    InMux I__10535 (
            .O(N__46080),
            .I(N__46064));
    InMux I__10534 (
            .O(N__46079),
            .I(N__46061));
    InMux I__10533 (
            .O(N__46078),
            .I(N__46058));
    LocalMux I__10532 (
            .O(N__46075),
            .I(N__46055));
    InMux I__10531 (
            .O(N__46072),
            .I(N__46050));
    InMux I__10530 (
            .O(N__46071),
            .I(N__46050));
    InMux I__10529 (
            .O(N__46070),
            .I(N__46047));
    LocalMux I__10528 (
            .O(N__46067),
            .I(N__46040));
    LocalMux I__10527 (
            .O(N__46064),
            .I(N__46040));
    LocalMux I__10526 (
            .O(N__46061),
            .I(N__46040));
    LocalMux I__10525 (
            .O(N__46058),
            .I(N__46037));
    Span4Mux_h I__10524 (
            .O(N__46055),
            .I(N__46032));
    LocalMux I__10523 (
            .O(N__46050),
            .I(N__46032));
    LocalMux I__10522 (
            .O(N__46047),
            .I(N__46025));
    Span4Mux_v I__10521 (
            .O(N__46040),
            .I(N__46025));
    Span4Mux_h I__10520 (
            .O(N__46037),
            .I(N__46025));
    Span4Mux_h I__10519 (
            .O(N__46032),
            .I(N__46022));
    Span4Mux_h I__10518 (
            .O(N__46025),
            .I(N__46019));
    Odrv4 I__10517 (
            .O(N__46022),
            .I(n14506));
    Odrv4 I__10516 (
            .O(N__46019),
            .I(n14506));
    InMux I__10515 (
            .O(N__46014),
            .I(N__46009));
    InMux I__10514 (
            .O(N__46013),
            .I(N__46005));
    InMux I__10513 (
            .O(N__46012),
            .I(N__46002));
    LocalMux I__10512 (
            .O(N__46009),
            .I(N__45995));
    InMux I__10511 (
            .O(N__46008),
            .I(N__45992));
    LocalMux I__10510 (
            .O(N__46005),
            .I(N__45987));
    LocalMux I__10509 (
            .O(N__46002),
            .I(N__45987));
    InMux I__10508 (
            .O(N__46001),
            .I(N__45984));
    InMux I__10507 (
            .O(N__46000),
            .I(N__45979));
    InMux I__10506 (
            .O(N__45999),
            .I(N__45979));
    InMux I__10505 (
            .O(N__45998),
            .I(N__45976));
    Span4Mux_h I__10504 (
            .O(N__45995),
            .I(N__45973));
    LocalMux I__10503 (
            .O(N__45992),
            .I(N__45970));
    Span4Mux_v I__10502 (
            .O(N__45987),
            .I(N__45961));
    LocalMux I__10501 (
            .O(N__45984),
            .I(N__45961));
    LocalMux I__10500 (
            .O(N__45979),
            .I(N__45961));
    LocalMux I__10499 (
            .O(N__45976),
            .I(N__45961));
    Odrv4 I__10498 (
            .O(N__45973),
            .I(n11896));
    Odrv12 I__10497 (
            .O(N__45970),
            .I(n11896));
    Odrv4 I__10496 (
            .O(N__45961),
            .I(n11896));
    InMux I__10495 (
            .O(N__45954),
            .I(N__45949));
    InMux I__10494 (
            .O(N__45953),
            .I(N__45944));
    InMux I__10493 (
            .O(N__45952),
            .I(N__45944));
    LocalMux I__10492 (
            .O(N__45949),
            .I(N__45939));
    LocalMux I__10491 (
            .O(N__45944),
            .I(N__45939));
    Span12Mux_v I__10490 (
            .O(N__45939),
            .I(N__45936));
    Odrv12 I__10489 (
            .O(N__45936),
            .I(n10697));
    InMux I__10488 (
            .O(N__45933),
            .I(N__45930));
    LocalMux I__10487 (
            .O(N__45930),
            .I(n18993));
    InMux I__10486 (
            .O(N__45927),
            .I(N__45924));
    LocalMux I__10485 (
            .O(N__45924),
            .I(N__45921));
    Span4Mux_h I__10484 (
            .O(N__45921),
            .I(N__45917));
    CascadeMux I__10483 (
            .O(N__45920),
            .I(N__45911));
    Span4Mux_h I__10482 (
            .O(N__45917),
            .I(N__45907));
    InMux I__10481 (
            .O(N__45916),
            .I(N__45904));
    InMux I__10480 (
            .O(N__45915),
            .I(N__45899));
    InMux I__10479 (
            .O(N__45914),
            .I(N__45899));
    InMux I__10478 (
            .O(N__45911),
            .I(N__45894));
    InMux I__10477 (
            .O(N__45910),
            .I(N__45894));
    Odrv4 I__10476 (
            .O(N__45907),
            .I(n20843));
    LocalMux I__10475 (
            .O(N__45904),
            .I(n20843));
    LocalMux I__10474 (
            .O(N__45899),
            .I(n20843));
    LocalMux I__10473 (
            .O(N__45894),
            .I(n20843));
    CascadeMux I__10472 (
            .O(N__45885),
            .I(n12_adj_1635_cascade_));
    InMux I__10471 (
            .O(N__45882),
            .I(N__45873));
    InMux I__10470 (
            .O(N__45881),
            .I(N__45870));
    InMux I__10469 (
            .O(N__45880),
            .I(N__45865));
    InMux I__10468 (
            .O(N__45879),
            .I(N__45865));
    CascadeMux I__10467 (
            .O(N__45878),
            .I(N__45862));
    InMux I__10466 (
            .O(N__45877),
            .I(N__45856));
    InMux I__10465 (
            .O(N__45876),
            .I(N__45856));
    LocalMux I__10464 (
            .O(N__45873),
            .I(N__45853));
    LocalMux I__10463 (
            .O(N__45870),
            .I(N__45850));
    LocalMux I__10462 (
            .O(N__45865),
            .I(N__45847));
    InMux I__10461 (
            .O(N__45862),
            .I(N__45843));
    InMux I__10460 (
            .O(N__45861),
            .I(N__45840));
    LocalMux I__10459 (
            .O(N__45856),
            .I(N__45837));
    Span4Mux_v I__10458 (
            .O(N__45853),
            .I(N__45834));
    Span4Mux_h I__10457 (
            .O(N__45850),
            .I(N__45829));
    Span4Mux_h I__10456 (
            .O(N__45847),
            .I(N__45829));
    InMux I__10455 (
            .O(N__45846),
            .I(N__45826));
    LocalMux I__10454 (
            .O(N__45843),
            .I(N__45819));
    LocalMux I__10453 (
            .O(N__45840),
            .I(N__45819));
    Span4Mux_h I__10452 (
            .O(N__45837),
            .I(N__45819));
    Odrv4 I__10451 (
            .O(N__45834),
            .I(n20917));
    Odrv4 I__10450 (
            .O(N__45829),
            .I(n20917));
    LocalMux I__10449 (
            .O(N__45826),
            .I(n20917));
    Odrv4 I__10448 (
            .O(N__45819),
            .I(n20917));
    CEMux I__10447 (
            .O(N__45810),
            .I(N__45807));
    LocalMux I__10446 (
            .O(N__45807),
            .I(N__45803));
    InMux I__10445 (
            .O(N__45806),
            .I(N__45800));
    Odrv4 I__10444 (
            .O(N__45803),
            .I(n12178));
    LocalMux I__10443 (
            .O(N__45800),
            .I(n12178));
    InMux I__10442 (
            .O(N__45795),
            .I(N__45788));
    CascadeMux I__10441 (
            .O(N__45794),
            .I(N__45784));
    InMux I__10440 (
            .O(N__45793),
            .I(N__45781));
    InMux I__10439 (
            .O(N__45792),
            .I(N__45778));
    CascadeMux I__10438 (
            .O(N__45791),
            .I(N__45775));
    LocalMux I__10437 (
            .O(N__45788),
            .I(N__45772));
    InMux I__10436 (
            .O(N__45787),
            .I(N__45769));
    InMux I__10435 (
            .O(N__45784),
            .I(N__45765));
    LocalMux I__10434 (
            .O(N__45781),
            .I(N__45760));
    LocalMux I__10433 (
            .O(N__45778),
            .I(N__45760));
    InMux I__10432 (
            .O(N__45775),
            .I(N__45757));
    Span4Mux_v I__10431 (
            .O(N__45772),
            .I(N__45754));
    LocalMux I__10430 (
            .O(N__45769),
            .I(N__45751));
    InMux I__10429 (
            .O(N__45768),
            .I(N__45748));
    LocalMux I__10428 (
            .O(N__45765),
            .I(N__45745));
    Span4Mux_v I__10427 (
            .O(N__45760),
            .I(N__45740));
    LocalMux I__10426 (
            .O(N__45757),
            .I(N__45740));
    Span4Mux_h I__10425 (
            .O(N__45754),
            .I(N__45737));
    Span4Mux_v I__10424 (
            .O(N__45751),
            .I(N__45732));
    LocalMux I__10423 (
            .O(N__45748),
            .I(N__45732));
    Span4Mux_v I__10422 (
            .O(N__45745),
            .I(N__45729));
    Span4Mux_h I__10421 (
            .O(N__45740),
            .I(N__45726));
    Sp12to4 I__10420 (
            .O(N__45737),
            .I(N__45721));
    Span4Mux_h I__10419 (
            .O(N__45732),
            .I(N__45716));
    Span4Mux_h I__10418 (
            .O(N__45729),
            .I(N__45716));
    Span4Mux_h I__10417 (
            .O(N__45726),
            .I(N__45713));
    InMux I__10416 (
            .O(N__45725),
            .I(N__45710));
    InMux I__10415 (
            .O(N__45724),
            .I(N__45707));
    Odrv12 I__10414 (
            .O(N__45721),
            .I(comm_rx_buf_1));
    Odrv4 I__10413 (
            .O(N__45716),
            .I(comm_rx_buf_1));
    Odrv4 I__10412 (
            .O(N__45713),
            .I(comm_rx_buf_1));
    LocalMux I__10411 (
            .O(N__45710),
            .I(comm_rx_buf_1));
    LocalMux I__10410 (
            .O(N__45707),
            .I(comm_rx_buf_1));
    InMux I__10409 (
            .O(N__45696),
            .I(N__45693));
    LocalMux I__10408 (
            .O(N__45693),
            .I(N__45690));
    Span4Mux_h I__10407 (
            .O(N__45690),
            .I(N__45687));
    Odrv4 I__10406 (
            .O(N__45687),
            .I(buf_data_vac_17));
    CascadeMux I__10405 (
            .O(N__45684),
            .I(N__45681));
    InMux I__10404 (
            .O(N__45681),
            .I(N__45678));
    LocalMux I__10403 (
            .O(N__45678),
            .I(N__45675));
    Span4Mux_h I__10402 (
            .O(N__45675),
            .I(N__45672));
    Span4Mux_h I__10401 (
            .O(N__45672),
            .I(N__45669));
    Odrv4 I__10400 (
            .O(N__45669),
            .I(comm_buf_3_1));
    InMux I__10399 (
            .O(N__45666),
            .I(N__45663));
    LocalMux I__10398 (
            .O(N__45663),
            .I(N__45660));
    Odrv12 I__10397 (
            .O(N__45660),
            .I(n20878));
    CascadeMux I__10396 (
            .O(N__45657),
            .I(n21352_cascade_));
    CascadeMux I__10395 (
            .O(N__45654),
            .I(n12_cascade_));
    CEMux I__10394 (
            .O(N__45651),
            .I(N__45648));
    LocalMux I__10393 (
            .O(N__45648),
            .I(n12136));
    CascadeMux I__10392 (
            .O(N__45645),
            .I(n12136_cascade_));
    SRMux I__10391 (
            .O(N__45642),
            .I(N__45639));
    LocalMux I__10390 (
            .O(N__45639),
            .I(n14771));
    InMux I__10389 (
            .O(N__45636),
            .I(N__45633));
    LocalMux I__10388 (
            .O(N__45633),
            .I(N__45628));
    InMux I__10387 (
            .O(N__45632),
            .I(N__45623));
    InMux I__10386 (
            .O(N__45631),
            .I(N__45623));
    Span4Mux_v I__10385 (
            .O(N__45628),
            .I(N__45620));
    LocalMux I__10384 (
            .O(N__45623),
            .I(N__45617));
    Sp12to4 I__10383 (
            .O(N__45620),
            .I(N__45614));
    Span4Mux_v I__10382 (
            .O(N__45617),
            .I(N__45611));
    Odrv12 I__10381 (
            .O(N__45614),
            .I(n19783));
    Odrv4 I__10380 (
            .O(N__45611),
            .I(n19783));
    CascadeMux I__10379 (
            .O(N__45606),
            .I(n18991_cascade_));
    CascadeMux I__10378 (
            .O(N__45603),
            .I(n4_adj_1545_cascade_));
    InMux I__10377 (
            .O(N__45600),
            .I(N__45597));
    LocalMux I__10376 (
            .O(N__45597),
            .I(N__45594));
    Span4Mux_h I__10375 (
            .O(N__45594),
            .I(N__45590));
    InMux I__10374 (
            .O(N__45593),
            .I(N__45587));
    Span4Mux_h I__10373 (
            .O(N__45590),
            .I(N__45584));
    LocalMux I__10372 (
            .O(N__45587),
            .I(comm_buf_6_6));
    Odrv4 I__10371 (
            .O(N__45584),
            .I(comm_buf_6_6));
    InMux I__10370 (
            .O(N__45579),
            .I(N__45576));
    LocalMux I__10369 (
            .O(N__45576),
            .I(n4_adj_1590));
    CascadeMux I__10368 (
            .O(N__45573),
            .I(n21539_cascade_));
    InMux I__10367 (
            .O(N__45570),
            .I(N__45567));
    LocalMux I__10366 (
            .O(N__45567),
            .I(n22339));
    InMux I__10365 (
            .O(N__45564),
            .I(N__45561));
    LocalMux I__10364 (
            .O(N__45561),
            .I(N__45558));
    Span4Mux_h I__10363 (
            .O(N__45558),
            .I(N__45555));
    Odrv4 I__10362 (
            .O(N__45555),
            .I(buf_data_vac_16));
    InMux I__10361 (
            .O(N__45552),
            .I(N__45549));
    LocalMux I__10360 (
            .O(N__45549),
            .I(comm_buf_3_0));
    InMux I__10359 (
            .O(N__45546),
            .I(N__45543));
    LocalMux I__10358 (
            .O(N__45543),
            .I(N__45540));
    Span4Mux_v I__10357 (
            .O(N__45540),
            .I(N__45537));
    Span4Mux_h I__10356 (
            .O(N__45537),
            .I(N__45534));
    Odrv4 I__10355 (
            .O(N__45534),
            .I(buf_data_vac_20));
    InMux I__10354 (
            .O(N__45531),
            .I(N__45528));
    LocalMux I__10353 (
            .O(N__45528),
            .I(N__45525));
    Span4Mux_v I__10352 (
            .O(N__45525),
            .I(N__45522));
    Odrv4 I__10351 (
            .O(N__45522),
            .I(comm_buf_3_4));
    InMux I__10350 (
            .O(N__45519),
            .I(N__45516));
    LocalMux I__10349 (
            .O(N__45516),
            .I(N__45513));
    Span4Mux_v I__10348 (
            .O(N__45513),
            .I(N__45510));
    Span4Mux_v I__10347 (
            .O(N__45510),
            .I(N__45507));
    Odrv4 I__10346 (
            .O(N__45507),
            .I(buf_data_vac_23));
    CascadeMux I__10345 (
            .O(N__45504),
            .I(N__45501));
    InMux I__10344 (
            .O(N__45501),
            .I(N__45498));
    LocalMux I__10343 (
            .O(N__45498),
            .I(N__45495));
    Span12Mux_h I__10342 (
            .O(N__45495),
            .I(N__45492));
    Odrv12 I__10341 (
            .O(N__45492),
            .I(comm_buf_3_7));
    InMux I__10340 (
            .O(N__45489),
            .I(N__45486));
    LocalMux I__10339 (
            .O(N__45486),
            .I(N__45483));
    Span4Mux_h I__10338 (
            .O(N__45483),
            .I(N__45480));
    Span4Mux_v I__10337 (
            .O(N__45480),
            .I(N__45477));
    Odrv4 I__10336 (
            .O(N__45477),
            .I(buf_data_vac_22));
    InMux I__10335 (
            .O(N__45474),
            .I(N__45471));
    LocalMux I__10334 (
            .O(N__45471),
            .I(N__45468));
    Odrv4 I__10333 (
            .O(N__45468),
            .I(comm_buf_3_6));
    InMux I__10332 (
            .O(N__45465),
            .I(N__45462));
    LocalMux I__10331 (
            .O(N__45462),
            .I(N__45459));
    Span4Mux_h I__10330 (
            .O(N__45459),
            .I(N__45456));
    Span4Mux_v I__10329 (
            .O(N__45456),
            .I(N__45453));
    Odrv4 I__10328 (
            .O(N__45453),
            .I(buf_data_vac_21));
    InMux I__10327 (
            .O(N__45450),
            .I(N__45447));
    LocalMux I__10326 (
            .O(N__45447),
            .I(comm_buf_3_5));
    InMux I__10325 (
            .O(N__45444),
            .I(N__45441));
    LocalMux I__10324 (
            .O(N__45441),
            .I(N__45438));
    Odrv4 I__10323 (
            .O(N__45438),
            .I(buf_data_vac_19));
    CascadeMux I__10322 (
            .O(N__45435),
            .I(N__45432));
    InMux I__10321 (
            .O(N__45432),
            .I(N__45429));
    LocalMux I__10320 (
            .O(N__45429),
            .I(N__45426));
    Span4Mux_h I__10319 (
            .O(N__45426),
            .I(N__45423));
    Odrv4 I__10318 (
            .O(N__45423),
            .I(comm_buf_3_3));
    InMux I__10317 (
            .O(N__45420),
            .I(N__45417));
    LocalMux I__10316 (
            .O(N__45417),
            .I(N__45414));
    Span4Mux_h I__10315 (
            .O(N__45414),
            .I(N__45411));
    Odrv4 I__10314 (
            .O(N__45411),
            .I(buf_data_vac_18));
    CascadeMux I__10313 (
            .O(N__45408),
            .I(N__45405));
    InMux I__10312 (
            .O(N__45405),
            .I(N__45402));
    LocalMux I__10311 (
            .O(N__45402),
            .I(N__45399));
    Odrv12 I__10310 (
            .O(N__45399),
            .I(comm_buf_3_2));
    CascadeMux I__10309 (
            .O(N__45396),
            .I(\ADC_VDC.genclk.n21446_cascade_ ));
    InMux I__10308 (
            .O(N__45393),
            .I(N__45390));
    LocalMux I__10307 (
            .O(N__45390),
            .I(\ADC_VDC.genclk.n26 ));
    InMux I__10306 (
            .O(N__45387),
            .I(N__45384));
    LocalMux I__10305 (
            .O(N__45384),
            .I(\ADC_VDC.genclk.n27 ));
    InMux I__10304 (
            .O(N__45381),
            .I(N__45378));
    LocalMux I__10303 (
            .O(N__45378),
            .I(\ADC_VDC.genclk.n28_adj_1397 ));
    SRMux I__10302 (
            .O(N__45375),
            .I(N__45372));
    LocalMux I__10301 (
            .O(N__45372),
            .I(N__45369));
    Span4Mux_h I__10300 (
            .O(N__45369),
            .I(N__45366));
    Odrv4 I__10299 (
            .O(N__45366),
            .I(\comm_spi.data_tx_7__N_767 ));
    CascadeMux I__10298 (
            .O(N__45363),
            .I(N__45359));
    CascadeMux I__10297 (
            .O(N__45362),
            .I(N__45354));
    InMux I__10296 (
            .O(N__45359),
            .I(N__45350));
    CascadeMux I__10295 (
            .O(N__45358),
            .I(N__45347));
    InMux I__10294 (
            .O(N__45357),
            .I(N__45344));
    InMux I__10293 (
            .O(N__45354),
            .I(N__45341));
    InMux I__10292 (
            .O(N__45353),
            .I(N__45335));
    LocalMux I__10291 (
            .O(N__45350),
            .I(N__45332));
    InMux I__10290 (
            .O(N__45347),
            .I(N__45329));
    LocalMux I__10289 (
            .O(N__45344),
            .I(N__45324));
    LocalMux I__10288 (
            .O(N__45341),
            .I(N__45324));
    InMux I__10287 (
            .O(N__45340),
            .I(N__45321));
    CascadeMux I__10286 (
            .O(N__45339),
            .I(N__45318));
    InMux I__10285 (
            .O(N__45338),
            .I(N__45315));
    LocalMux I__10284 (
            .O(N__45335),
            .I(N__45308));
    Span4Mux_h I__10283 (
            .O(N__45332),
            .I(N__45308));
    LocalMux I__10282 (
            .O(N__45329),
            .I(N__45308));
    Span4Mux_v I__10281 (
            .O(N__45324),
            .I(N__45303));
    LocalMux I__10280 (
            .O(N__45321),
            .I(N__45303));
    InMux I__10279 (
            .O(N__45318),
            .I(N__45300));
    LocalMux I__10278 (
            .O(N__45315),
            .I(N__45297));
    Span4Mux_v I__10277 (
            .O(N__45308),
            .I(N__45294));
    Span4Mux_h I__10276 (
            .O(N__45303),
            .I(N__45291));
    LocalMux I__10275 (
            .O(N__45300),
            .I(N__45288));
    Span4Mux_h I__10274 (
            .O(N__45297),
            .I(N__45285));
    Span4Mux_h I__10273 (
            .O(N__45294),
            .I(N__45280));
    Span4Mux_h I__10272 (
            .O(N__45291),
            .I(N__45280));
    Odrv12 I__10271 (
            .O(N__45288),
            .I(comm_buf_0_6));
    Odrv4 I__10270 (
            .O(N__45285),
            .I(comm_buf_0_6));
    Odrv4 I__10269 (
            .O(N__45280),
            .I(comm_buf_0_6));
    CascadeMux I__10268 (
            .O(N__45273),
            .I(n1_adj_1588_cascade_));
    InMux I__10267 (
            .O(N__45270),
            .I(N__45267));
    LocalMux I__10266 (
            .O(N__45267),
            .I(N__45264));
    Span4Mux_h I__10265 (
            .O(N__45264),
            .I(N__45261));
    Span4Mux_v I__10264 (
            .O(N__45261),
            .I(N__45256));
    InMux I__10263 (
            .O(N__45260),
            .I(N__45253));
    InMux I__10262 (
            .O(N__45259),
            .I(N__45250));
    Odrv4 I__10261 (
            .O(N__45256),
            .I(comm_tx_buf_6));
    LocalMux I__10260 (
            .O(N__45253),
            .I(comm_tx_buf_6));
    LocalMux I__10259 (
            .O(N__45250),
            .I(comm_tx_buf_6));
    CEMux I__10258 (
            .O(N__45243),
            .I(N__45240));
    LocalMux I__10257 (
            .O(N__45240),
            .I(N__45237));
    Span4Mux_v I__10256 (
            .O(N__45237),
            .I(N__45230));
    CEMux I__10255 (
            .O(N__45236),
            .I(N__45227));
    CEMux I__10254 (
            .O(N__45235),
            .I(N__45223));
    CEMux I__10253 (
            .O(N__45234),
            .I(N__45220));
    CEMux I__10252 (
            .O(N__45233),
            .I(N__45217));
    Span4Mux_v I__10251 (
            .O(N__45230),
            .I(N__45212));
    LocalMux I__10250 (
            .O(N__45227),
            .I(N__45212));
    CEMux I__10249 (
            .O(N__45226),
            .I(N__45209));
    LocalMux I__10248 (
            .O(N__45223),
            .I(N__45206));
    LocalMux I__10247 (
            .O(N__45220),
            .I(N__45203));
    LocalMux I__10246 (
            .O(N__45217),
            .I(N__45200));
    Span4Mux_v I__10245 (
            .O(N__45212),
            .I(N__45197));
    LocalMux I__10244 (
            .O(N__45209),
            .I(N__45194));
    Span4Mux_v I__10243 (
            .O(N__45206),
            .I(N__45187));
    Span4Mux_v I__10242 (
            .O(N__45203),
            .I(N__45187));
    Span4Mux_v I__10241 (
            .O(N__45200),
            .I(N__45187));
    Span4Mux_h I__10240 (
            .O(N__45197),
            .I(N__45184));
    Odrv4 I__10239 (
            .O(N__45194),
            .I(n12336));
    Odrv4 I__10238 (
            .O(N__45187),
            .I(n12336));
    Odrv4 I__10237 (
            .O(N__45184),
            .I(n12336));
    SRMux I__10236 (
            .O(N__45177),
            .I(N__45174));
    LocalMux I__10235 (
            .O(N__45174),
            .I(N__45168));
    SRMux I__10234 (
            .O(N__45173),
            .I(N__45165));
    SRMux I__10233 (
            .O(N__45172),
            .I(N__45161));
    SRMux I__10232 (
            .O(N__45171),
            .I(N__45158));
    Span4Mux_h I__10231 (
            .O(N__45168),
            .I(N__45152));
    LocalMux I__10230 (
            .O(N__45165),
            .I(N__45152));
    SRMux I__10229 (
            .O(N__45164),
            .I(N__45149));
    LocalMux I__10228 (
            .O(N__45161),
            .I(N__45146));
    LocalMux I__10227 (
            .O(N__45158),
            .I(N__45143));
    SRMux I__10226 (
            .O(N__45157),
            .I(N__45140));
    Span4Mux_v I__10225 (
            .O(N__45152),
            .I(N__45135));
    LocalMux I__10224 (
            .O(N__45149),
            .I(N__45135));
    Span4Mux_h I__10223 (
            .O(N__45146),
            .I(N__45132));
    Span4Mux_h I__10222 (
            .O(N__45143),
            .I(N__45129));
    LocalMux I__10221 (
            .O(N__45140),
            .I(N__45126));
    Span4Mux_h I__10220 (
            .O(N__45135),
            .I(N__45123));
    Odrv4 I__10219 (
            .O(N__45132),
            .I(n14799));
    Odrv4 I__10218 (
            .O(N__45129),
            .I(n14799));
    Odrv4 I__10217 (
            .O(N__45126),
            .I(n14799));
    Odrv4 I__10216 (
            .O(N__45123),
            .I(n14799));
    InMux I__10215 (
            .O(N__45114),
            .I(N__45111));
    LocalMux I__10214 (
            .O(N__45111),
            .I(N__45108));
    Odrv12 I__10213 (
            .O(N__45108),
            .I(comm_buf_2_6));
    InMux I__10212 (
            .O(N__45105),
            .I(N__45102));
    LocalMux I__10211 (
            .O(N__45102),
            .I(n2_adj_1589));
    InMux I__10210 (
            .O(N__45099),
            .I(N__45096));
    LocalMux I__10209 (
            .O(N__45096),
            .I(n8_adj_1571));
    InMux I__10208 (
            .O(N__45093),
            .I(N__45089));
    InMux I__10207 (
            .O(N__45092),
            .I(N__45086));
    LocalMux I__10206 (
            .O(N__45089),
            .I(N__45081));
    LocalMux I__10205 (
            .O(N__45086),
            .I(N__45081));
    Span4Mux_h I__10204 (
            .O(N__45081),
            .I(N__45078));
    Odrv4 I__10203 (
            .O(N__45078),
            .I(n7_adj_1570));
    CascadeMux I__10202 (
            .O(N__45075),
            .I(N__45072));
    CascadeBuf I__10201 (
            .O(N__45072),
            .I(N__45069));
    CascadeMux I__10200 (
            .O(N__45069),
            .I(N__45066));
    CascadeBuf I__10199 (
            .O(N__45066),
            .I(N__45063));
    CascadeMux I__10198 (
            .O(N__45063),
            .I(N__45060));
    CascadeBuf I__10197 (
            .O(N__45060),
            .I(N__45057));
    CascadeMux I__10196 (
            .O(N__45057),
            .I(N__45054));
    CascadeBuf I__10195 (
            .O(N__45054),
            .I(N__45051));
    CascadeMux I__10194 (
            .O(N__45051),
            .I(N__45048));
    CascadeBuf I__10193 (
            .O(N__45048),
            .I(N__45045));
    CascadeMux I__10192 (
            .O(N__45045),
            .I(N__45042));
    CascadeBuf I__10191 (
            .O(N__45042),
            .I(N__45039));
    CascadeMux I__10190 (
            .O(N__45039),
            .I(N__45036));
    CascadeBuf I__10189 (
            .O(N__45036),
            .I(N__45032));
    CascadeMux I__10188 (
            .O(N__45035),
            .I(N__45029));
    CascadeMux I__10187 (
            .O(N__45032),
            .I(N__45026));
    CascadeBuf I__10186 (
            .O(N__45029),
            .I(N__45023));
    CascadeBuf I__10185 (
            .O(N__45026),
            .I(N__45020));
    CascadeMux I__10184 (
            .O(N__45023),
            .I(N__45017));
    CascadeMux I__10183 (
            .O(N__45020),
            .I(N__45014));
    InMux I__10182 (
            .O(N__45017),
            .I(N__45011));
    CascadeBuf I__10181 (
            .O(N__45014),
            .I(N__45008));
    LocalMux I__10180 (
            .O(N__45011),
            .I(N__45005));
    CascadeMux I__10179 (
            .O(N__45008),
            .I(N__45002));
    Sp12to4 I__10178 (
            .O(N__45005),
            .I(N__44999));
    InMux I__10177 (
            .O(N__45002),
            .I(N__44996));
    Span12Mux_v I__10176 (
            .O(N__44999),
            .I(N__44993));
    LocalMux I__10175 (
            .O(N__44996),
            .I(N__44990));
    Span12Mux_h I__10174 (
            .O(N__44993),
            .I(N__44987));
    Span4Mux_h I__10173 (
            .O(N__44990),
            .I(N__44984));
    Odrv12 I__10172 (
            .O(N__44987),
            .I(data_index_9_N_216_2));
    Odrv4 I__10171 (
            .O(N__44984),
            .I(data_index_9_N_216_2));
    CascadeMux I__10170 (
            .O(N__44979),
            .I(N__44972));
    InMux I__10169 (
            .O(N__44978),
            .I(N__44967));
    InMux I__10168 (
            .O(N__44977),
            .I(N__44964));
    InMux I__10167 (
            .O(N__44976),
            .I(N__44961));
    InMux I__10166 (
            .O(N__44975),
            .I(N__44958));
    InMux I__10165 (
            .O(N__44972),
            .I(N__44954));
    InMux I__10164 (
            .O(N__44971),
            .I(N__44951));
    InMux I__10163 (
            .O(N__44970),
            .I(N__44948));
    LocalMux I__10162 (
            .O(N__44967),
            .I(N__44942));
    LocalMux I__10161 (
            .O(N__44964),
            .I(N__44942));
    LocalMux I__10160 (
            .O(N__44961),
            .I(N__44939));
    LocalMux I__10159 (
            .O(N__44958),
            .I(N__44936));
    InMux I__10158 (
            .O(N__44957),
            .I(N__44928));
    LocalMux I__10157 (
            .O(N__44954),
            .I(N__44923));
    LocalMux I__10156 (
            .O(N__44951),
            .I(N__44923));
    LocalMux I__10155 (
            .O(N__44948),
            .I(N__44920));
    InMux I__10154 (
            .O(N__44947),
            .I(N__44917));
    Span4Mux_v I__10153 (
            .O(N__44942),
            .I(N__44910));
    Span4Mux_h I__10152 (
            .O(N__44939),
            .I(N__44910));
    Span4Mux_v I__10151 (
            .O(N__44936),
            .I(N__44910));
    InMux I__10150 (
            .O(N__44935),
            .I(N__44902));
    InMux I__10149 (
            .O(N__44934),
            .I(N__44902));
    InMux I__10148 (
            .O(N__44933),
            .I(N__44895));
    InMux I__10147 (
            .O(N__44932),
            .I(N__44895));
    InMux I__10146 (
            .O(N__44931),
            .I(N__44895));
    LocalMux I__10145 (
            .O(N__44928),
            .I(N__44890));
    Span4Mux_v I__10144 (
            .O(N__44923),
            .I(N__44890));
    Span12Mux_v I__10143 (
            .O(N__44920),
            .I(N__44887));
    LocalMux I__10142 (
            .O(N__44917),
            .I(N__44882));
    Span4Mux_h I__10141 (
            .O(N__44910),
            .I(N__44882));
    InMux I__10140 (
            .O(N__44909),
            .I(N__44875));
    InMux I__10139 (
            .O(N__44908),
            .I(N__44875));
    InMux I__10138 (
            .O(N__44907),
            .I(N__44875));
    LocalMux I__10137 (
            .O(N__44902),
            .I(n11819));
    LocalMux I__10136 (
            .O(N__44895),
            .I(n11819));
    Odrv4 I__10135 (
            .O(N__44890),
            .I(n11819));
    Odrv12 I__10134 (
            .O(N__44887),
            .I(n11819));
    Odrv4 I__10133 (
            .O(N__44882),
            .I(n11819));
    LocalMux I__10132 (
            .O(N__44875),
            .I(n11819));
    InMux I__10131 (
            .O(N__44862),
            .I(N__44857));
    InMux I__10130 (
            .O(N__44861),
            .I(N__44853));
    InMux I__10129 (
            .O(N__44860),
            .I(N__44850));
    LocalMux I__10128 (
            .O(N__44857),
            .I(N__44846));
    InMux I__10127 (
            .O(N__44856),
            .I(N__44843));
    LocalMux I__10126 (
            .O(N__44853),
            .I(N__44838));
    LocalMux I__10125 (
            .O(N__44850),
            .I(N__44838));
    InMux I__10124 (
            .O(N__44849),
            .I(N__44835));
    Span4Mux_v I__10123 (
            .O(N__44846),
            .I(N__44830));
    LocalMux I__10122 (
            .O(N__44843),
            .I(N__44830));
    Span4Mux_h I__10121 (
            .O(N__44838),
            .I(N__44827));
    LocalMux I__10120 (
            .O(N__44835),
            .I(N__44824));
    Span4Mux_h I__10119 (
            .O(N__44830),
            .I(N__44821));
    Span4Mux_h I__10118 (
            .O(N__44827),
            .I(N__44816));
    Span12Mux_h I__10117 (
            .O(N__44824),
            .I(N__44813));
    Span4Mux_h I__10116 (
            .O(N__44821),
            .I(N__44810));
    InMux I__10115 (
            .O(N__44820),
            .I(N__44807));
    InMux I__10114 (
            .O(N__44819),
            .I(N__44804));
    Odrv4 I__10113 (
            .O(N__44816),
            .I(n12381));
    Odrv12 I__10112 (
            .O(N__44813),
            .I(n12381));
    Odrv4 I__10111 (
            .O(N__44810),
            .I(n12381));
    LocalMux I__10110 (
            .O(N__44807),
            .I(n12381));
    LocalMux I__10109 (
            .O(N__44804),
            .I(n12381));
    CascadeMux I__10108 (
            .O(N__44793),
            .I(N__44789));
    CascadeMux I__10107 (
            .O(N__44792),
            .I(N__44783));
    InMux I__10106 (
            .O(N__44789),
            .I(N__44780));
    CascadeMux I__10105 (
            .O(N__44788),
            .I(N__44776));
    InMux I__10104 (
            .O(N__44787),
            .I(N__44773));
    CascadeMux I__10103 (
            .O(N__44786),
            .I(N__44770));
    InMux I__10102 (
            .O(N__44783),
            .I(N__44766));
    LocalMux I__10101 (
            .O(N__44780),
            .I(N__44763));
    InMux I__10100 (
            .O(N__44779),
            .I(N__44760));
    InMux I__10099 (
            .O(N__44776),
            .I(N__44756));
    LocalMux I__10098 (
            .O(N__44773),
            .I(N__44753));
    InMux I__10097 (
            .O(N__44770),
            .I(N__44750));
    CascadeMux I__10096 (
            .O(N__44769),
            .I(N__44746));
    LocalMux I__10095 (
            .O(N__44766),
            .I(N__44743));
    Span4Mux_v I__10094 (
            .O(N__44763),
            .I(N__44740));
    LocalMux I__10093 (
            .O(N__44760),
            .I(N__44737));
    InMux I__10092 (
            .O(N__44759),
            .I(N__44734));
    LocalMux I__10091 (
            .O(N__44756),
            .I(N__44729));
    Span4Mux_v I__10090 (
            .O(N__44753),
            .I(N__44729));
    LocalMux I__10089 (
            .O(N__44750),
            .I(N__44726));
    InMux I__10088 (
            .O(N__44749),
            .I(N__44723));
    InMux I__10087 (
            .O(N__44746),
            .I(N__44720));
    Span4Mux_v I__10086 (
            .O(N__44743),
            .I(N__44713));
    Span4Mux_h I__10085 (
            .O(N__44740),
            .I(N__44713));
    Span4Mux_v I__10084 (
            .O(N__44737),
            .I(N__44713));
    LocalMux I__10083 (
            .O(N__44734),
            .I(N__44710));
    Span4Mux_h I__10082 (
            .O(N__44729),
            .I(N__44703));
    Span4Mux_h I__10081 (
            .O(N__44726),
            .I(N__44703));
    LocalMux I__10080 (
            .O(N__44723),
            .I(N__44703));
    LocalMux I__10079 (
            .O(N__44720),
            .I(N__44700));
    Span4Mux_h I__10078 (
            .O(N__44713),
            .I(N__44695));
    Span4Mux_v I__10077 (
            .O(N__44710),
            .I(N__44695));
    Span4Mux_v I__10076 (
            .O(N__44703),
            .I(N__44692));
    Odrv12 I__10075 (
            .O(N__44700),
            .I(comm_buf_0_2));
    Odrv4 I__10074 (
            .O(N__44695),
            .I(comm_buf_0_2));
    Odrv4 I__10073 (
            .O(N__44692),
            .I(comm_buf_0_2));
    IoInMux I__10072 (
            .O(N__44685),
            .I(N__44682));
    LocalMux I__10071 (
            .O(N__44682),
            .I(N__44679));
    Span4Mux_s3_v I__10070 (
            .O(N__44679),
            .I(N__44675));
    InMux I__10069 (
            .O(N__44678),
            .I(N__44672));
    Sp12to4 I__10068 (
            .O(N__44675),
            .I(N__44669));
    LocalMux I__10067 (
            .O(N__44672),
            .I(N__44665));
    Span12Mux_h I__10066 (
            .O(N__44669),
            .I(N__44662));
    InMux I__10065 (
            .O(N__44668),
            .I(N__44659));
    Span4Mux_v I__10064 (
            .O(N__44665),
            .I(N__44656));
    Odrv12 I__10063 (
            .O(N__44662),
            .I(IAC_FLT0));
    LocalMux I__10062 (
            .O(N__44659),
            .I(IAC_FLT0));
    Odrv4 I__10061 (
            .O(N__44656),
            .I(IAC_FLT0));
    InMux I__10060 (
            .O(N__44649),
            .I(N__44646));
    LocalMux I__10059 (
            .O(N__44646),
            .I(N__44643));
    Span4Mux_v I__10058 (
            .O(N__44643),
            .I(N__44640));
    Span4Mux_v I__10057 (
            .O(N__44640),
            .I(N__44637));
    Span4Mux_v I__10056 (
            .O(N__44637),
            .I(N__44634));
    Span4Mux_v I__10055 (
            .O(N__44634),
            .I(N__44629));
    InMux I__10054 (
            .O(N__44633),
            .I(N__44626));
    InMux I__10053 (
            .O(N__44632),
            .I(N__44623));
    Odrv4 I__10052 (
            .O(N__44629),
            .I(wdtick_flag));
    LocalMux I__10051 (
            .O(N__44626),
            .I(wdtick_flag));
    LocalMux I__10050 (
            .O(N__44623),
            .I(wdtick_flag));
    CascadeMux I__10049 (
            .O(N__44616),
            .I(N__44613));
    InMux I__10048 (
            .O(N__44613),
            .I(N__44608));
    InMux I__10047 (
            .O(N__44612),
            .I(N__44605));
    InMux I__10046 (
            .O(N__44611),
            .I(N__44602));
    LocalMux I__10045 (
            .O(N__44608),
            .I(N__44599));
    LocalMux I__10044 (
            .O(N__44605),
            .I(buf_control_0));
    LocalMux I__10043 (
            .O(N__44602),
            .I(buf_control_0));
    Odrv4 I__10042 (
            .O(N__44599),
            .I(buf_control_0));
    IoInMux I__10041 (
            .O(N__44592),
            .I(N__44589));
    LocalMux I__10040 (
            .O(N__44589),
            .I(N__44586));
    Span4Mux_s3_v I__10039 (
            .O(N__44586),
            .I(N__44583));
    Span4Mux_h I__10038 (
            .O(N__44583),
            .I(N__44580));
    Odrv4 I__10037 (
            .O(N__44580),
            .I(CONT_SD));
    SRMux I__10036 (
            .O(N__44577),
            .I(N__44574));
    LocalMux I__10035 (
            .O(N__44574),
            .I(N__44571));
    Span4Mux_h I__10034 (
            .O(N__44571),
            .I(N__44568));
    Span4Mux_h I__10033 (
            .O(N__44568),
            .I(N__44565));
    Odrv4 I__10032 (
            .O(N__44565),
            .I(\comm_spi.imosi_N_753 ));
    InMux I__10031 (
            .O(N__44562),
            .I(N__44558));
    InMux I__10030 (
            .O(N__44561),
            .I(N__44555));
    LocalMux I__10029 (
            .O(N__44558),
            .I(N__44550));
    LocalMux I__10028 (
            .O(N__44555),
            .I(N__44550));
    Span4Mux_h I__10027 (
            .O(N__44550),
            .I(N__44547));
    Sp12to4 I__10026 (
            .O(N__44547),
            .I(N__44543));
    InMux I__10025 (
            .O(N__44546),
            .I(N__44540));
    Odrv12 I__10024 (
            .O(N__44543),
            .I(\comm_spi.n22872 ));
    LocalMux I__10023 (
            .O(N__44540),
            .I(\comm_spi.n22872 ));
    InMux I__10022 (
            .O(N__44535),
            .I(N__44532));
    LocalMux I__10021 (
            .O(N__44532),
            .I(N__44529));
    Span4Mux_v I__10020 (
            .O(N__44529),
            .I(N__44525));
    InMux I__10019 (
            .O(N__44528),
            .I(N__44522));
    Odrv4 I__10018 (
            .O(N__44525),
            .I(\comm_spi.n14630 ));
    LocalMux I__10017 (
            .O(N__44522),
            .I(\comm_spi.n14630 ));
    InMux I__10016 (
            .O(N__44517),
            .I(N__44513));
    InMux I__10015 (
            .O(N__44516),
            .I(N__44510));
    LocalMux I__10014 (
            .O(N__44513),
            .I(N__44505));
    LocalMux I__10013 (
            .O(N__44510),
            .I(N__44505));
    Span4Mux_v I__10012 (
            .O(N__44505),
            .I(N__44502));
    Odrv4 I__10011 (
            .O(N__44502),
            .I(\comm_spi.n14631 ));
    SRMux I__10010 (
            .O(N__44499),
            .I(N__44496));
    LocalMux I__10009 (
            .O(N__44496),
            .I(N__44493));
    Span4Mux_v I__10008 (
            .O(N__44493),
            .I(N__44490));
    Odrv4 I__10007 (
            .O(N__44490),
            .I(\comm_spi.data_tx_7__N_768 ));
    InMux I__10006 (
            .O(N__44487),
            .I(N__44482));
    InMux I__10005 (
            .O(N__44486),
            .I(N__44479));
    InMux I__10004 (
            .O(N__44485),
            .I(N__44476));
    LocalMux I__10003 (
            .O(N__44482),
            .I(\comm_spi.n22869 ));
    LocalMux I__10002 (
            .O(N__44479),
            .I(\comm_spi.n22869 ));
    LocalMux I__10001 (
            .O(N__44476),
            .I(\comm_spi.n22869 ));
    InMux I__10000 (
            .O(N__44469),
            .I(N__44465));
    InMux I__9999 (
            .O(N__44468),
            .I(N__44462));
    LocalMux I__9998 (
            .O(N__44465),
            .I(\comm_spi.n14634 ));
    LocalMux I__9997 (
            .O(N__44462),
            .I(\comm_spi.n14634 ));
    InMux I__9996 (
            .O(N__44457),
            .I(N__44453));
    InMux I__9995 (
            .O(N__44456),
            .I(N__44450));
    LocalMux I__9994 (
            .O(N__44453),
            .I(\comm_spi.n14635 ));
    LocalMux I__9993 (
            .O(N__44450),
            .I(\comm_spi.n14635 ));
    InMux I__9992 (
            .O(N__44445),
            .I(N__44442));
    LocalMux I__9991 (
            .O(N__44442),
            .I(N__44438));
    InMux I__9990 (
            .O(N__44441),
            .I(N__44435));
    Sp12to4 I__9989 (
            .O(N__44438),
            .I(N__44430));
    LocalMux I__9988 (
            .O(N__44435),
            .I(N__44430));
    Odrv12 I__9987 (
            .O(N__44430),
            .I(\comm_spi.n14638 ));
    InMux I__9986 (
            .O(N__44427),
            .I(N__44423));
    InMux I__9985 (
            .O(N__44426),
            .I(N__44420));
    LocalMux I__9984 (
            .O(N__44423),
            .I(N__44415));
    LocalMux I__9983 (
            .O(N__44420),
            .I(N__44415));
    Span4Mux_v I__9982 (
            .O(N__44415),
            .I(N__44412));
    Odrv4 I__9981 (
            .O(N__44412),
            .I(n14_adj_1578));
    CascadeMux I__9980 (
            .O(N__44409),
            .I(N__44406));
    InMux I__9979 (
            .O(N__44406),
            .I(N__44403));
    LocalMux I__9978 (
            .O(N__44403),
            .I(N__44400));
    Span4Mux_v I__9977 (
            .O(N__44400),
            .I(N__44397));
    Odrv4 I__9976 (
            .O(N__44397),
            .I(n9_adj_1415));
    CascadeMux I__9975 (
            .O(N__44394),
            .I(N__44391));
    InMux I__9974 (
            .O(N__44391),
            .I(N__44388));
    LocalMux I__9973 (
            .O(N__44388),
            .I(N__44385));
    Span4Mux_h I__9972 (
            .O(N__44385),
            .I(N__44382));
    Span4Mux_v I__9971 (
            .O(N__44382),
            .I(N__44379));
    Odrv4 I__9970 (
            .O(N__44379),
            .I(buf_data_iac_16));
    InMux I__9969 (
            .O(N__44376),
            .I(N__44373));
    LocalMux I__9968 (
            .O(N__44373),
            .I(n21165));
    CascadeMux I__9967 (
            .O(N__44370),
            .I(n21167_cascade_));
    InMux I__9966 (
            .O(N__44367),
            .I(N__44364));
    LocalMux I__9965 (
            .O(N__44364),
            .I(n22222));
    CascadeMux I__9964 (
            .O(N__44361),
            .I(N__44358));
    InMux I__9963 (
            .O(N__44358),
            .I(N__44355));
    LocalMux I__9962 (
            .O(N__44355),
            .I(n21070));
    InMux I__9961 (
            .O(N__44352),
            .I(N__44349));
    LocalMux I__9960 (
            .O(N__44349),
            .I(n21084));
    InMux I__9959 (
            .O(N__44346),
            .I(N__44343));
    LocalMux I__9958 (
            .O(N__44343),
            .I(n21085));
    InMux I__9957 (
            .O(N__44340),
            .I(N__44337));
    LocalMux I__9956 (
            .O(N__44337),
            .I(N__44334));
    Odrv4 I__9955 (
            .O(N__44334),
            .I(n22309));
    CascadeMux I__9954 (
            .O(N__44331),
            .I(N__44318));
    InMux I__9953 (
            .O(N__44330),
            .I(N__44311));
    InMux I__9952 (
            .O(N__44329),
            .I(N__44311));
    InMux I__9951 (
            .O(N__44328),
            .I(N__44308));
    InMux I__9950 (
            .O(N__44327),
            .I(N__44303));
    InMux I__9949 (
            .O(N__44326),
            .I(N__44303));
    InMux I__9948 (
            .O(N__44325),
            .I(N__44300));
    InMux I__9947 (
            .O(N__44324),
            .I(N__44288));
    InMux I__9946 (
            .O(N__44323),
            .I(N__44288));
    InMux I__9945 (
            .O(N__44322),
            .I(N__44288));
    InMux I__9944 (
            .O(N__44321),
            .I(N__44288));
    InMux I__9943 (
            .O(N__44318),
            .I(N__44285));
    InMux I__9942 (
            .O(N__44317),
            .I(N__44282));
    InMux I__9941 (
            .O(N__44316),
            .I(N__44279));
    LocalMux I__9940 (
            .O(N__44311),
            .I(N__44276));
    LocalMux I__9939 (
            .O(N__44308),
            .I(N__44271));
    LocalMux I__9938 (
            .O(N__44303),
            .I(N__44271));
    LocalMux I__9937 (
            .O(N__44300),
            .I(N__44268));
    InMux I__9936 (
            .O(N__44299),
            .I(N__44261));
    InMux I__9935 (
            .O(N__44298),
            .I(N__44261));
    InMux I__9934 (
            .O(N__44297),
            .I(N__44261));
    LocalMux I__9933 (
            .O(N__44288),
            .I(N__44258));
    LocalMux I__9932 (
            .O(N__44285),
            .I(N__44253));
    LocalMux I__9931 (
            .O(N__44282),
            .I(N__44253));
    LocalMux I__9930 (
            .O(N__44279),
            .I(N__44248));
    Span4Mux_v I__9929 (
            .O(N__44276),
            .I(N__44248));
    Span4Mux_v I__9928 (
            .O(N__44271),
            .I(N__44245));
    Span4Mux_v I__9927 (
            .O(N__44268),
            .I(N__44242));
    LocalMux I__9926 (
            .O(N__44261),
            .I(n12399));
    Odrv4 I__9925 (
            .O(N__44258),
            .I(n12399));
    Odrv12 I__9924 (
            .O(N__44253),
            .I(n12399));
    Odrv4 I__9923 (
            .O(N__44248),
            .I(n12399));
    Odrv4 I__9922 (
            .O(N__44245),
            .I(n12399));
    Odrv4 I__9921 (
            .O(N__44242),
            .I(n12399));
    CascadeMux I__9920 (
            .O(N__44229),
            .I(N__44223));
    CascadeMux I__9919 (
            .O(N__44228),
            .I(N__44219));
    CascadeMux I__9918 (
            .O(N__44227),
            .I(N__44216));
    CascadeMux I__9917 (
            .O(N__44226),
            .I(N__44213));
    InMux I__9916 (
            .O(N__44223),
            .I(N__44210));
    InMux I__9915 (
            .O(N__44222),
            .I(N__44207));
    InMux I__9914 (
            .O(N__44219),
            .I(N__44204));
    InMux I__9913 (
            .O(N__44216),
            .I(N__44201));
    InMux I__9912 (
            .O(N__44213),
            .I(N__44198));
    LocalMux I__9911 (
            .O(N__44210),
            .I(N__44194));
    LocalMux I__9910 (
            .O(N__44207),
            .I(N__44191));
    LocalMux I__9909 (
            .O(N__44204),
            .I(N__44188));
    LocalMux I__9908 (
            .O(N__44201),
            .I(N__44184));
    LocalMux I__9907 (
            .O(N__44198),
            .I(N__44181));
    CascadeMux I__9906 (
            .O(N__44197),
            .I(N__44178));
    Span4Mux_h I__9905 (
            .O(N__44194),
            .I(N__44174));
    Span4Mux_v I__9904 (
            .O(N__44191),
            .I(N__44171));
    Span4Mux_h I__9903 (
            .O(N__44188),
            .I(N__44168));
    InMux I__9902 (
            .O(N__44187),
            .I(N__44165));
    Span4Mux_h I__9901 (
            .O(N__44184),
            .I(N__44160));
    Span4Mux_v I__9900 (
            .O(N__44181),
            .I(N__44160));
    InMux I__9899 (
            .O(N__44178),
            .I(N__44157));
    InMux I__9898 (
            .O(N__44177),
            .I(N__44154));
    Span4Mux_h I__9897 (
            .O(N__44174),
            .I(N__44151));
    Span4Mux_h I__9896 (
            .O(N__44171),
            .I(N__44148));
    Span4Mux_h I__9895 (
            .O(N__44168),
            .I(N__44143));
    LocalMux I__9894 (
            .O(N__44165),
            .I(N__44143));
    Span4Mux_h I__9893 (
            .O(N__44160),
            .I(N__44140));
    LocalMux I__9892 (
            .O(N__44157),
            .I(N__44133));
    LocalMux I__9891 (
            .O(N__44154),
            .I(N__44133));
    Span4Mux_h I__9890 (
            .O(N__44151),
            .I(N__44133));
    Span4Mux_v I__9889 (
            .O(N__44148),
            .I(N__44128));
    Span4Mux_v I__9888 (
            .O(N__44143),
            .I(N__44128));
    Odrv4 I__9887 (
            .O(N__44140),
            .I(comm_buf_0_3));
    Odrv4 I__9886 (
            .O(N__44133),
            .I(comm_buf_0_3));
    Odrv4 I__9885 (
            .O(N__44128),
            .I(comm_buf_0_3));
    IoInMux I__9884 (
            .O(N__44121),
            .I(N__44118));
    LocalMux I__9883 (
            .O(N__44118),
            .I(N__44115));
    Span4Mux_s3_v I__9882 (
            .O(N__44115),
            .I(N__44112));
    Span4Mux_v I__9881 (
            .O(N__44112),
            .I(N__44109));
    Sp12to4 I__9880 (
            .O(N__44109),
            .I(N__44105));
    InMux I__9879 (
            .O(N__44108),
            .I(N__44101));
    Span12Mux_h I__9878 (
            .O(N__44105),
            .I(N__44098));
    InMux I__9877 (
            .O(N__44104),
            .I(N__44095));
    LocalMux I__9876 (
            .O(N__44101),
            .I(N__44092));
    Odrv12 I__9875 (
            .O(N__44098),
            .I(IAC_FLT1));
    LocalMux I__9874 (
            .O(N__44095),
            .I(IAC_FLT1));
    Odrv4 I__9873 (
            .O(N__44092),
            .I(IAC_FLT1));
    InMux I__9872 (
            .O(N__44085),
            .I(N__44082));
    LocalMux I__9871 (
            .O(N__44082),
            .I(N__44079));
    Span12Mux_h I__9870 (
            .O(N__44079),
            .I(N__44076));
    Odrv12 I__9869 (
            .O(N__44076),
            .I(n20914));
    CascadeMux I__9868 (
            .O(N__44073),
            .I(N__44070));
    InMux I__9867 (
            .O(N__44070),
            .I(N__44066));
    CascadeMux I__9866 (
            .O(N__44069),
            .I(N__44063));
    LocalMux I__9865 (
            .O(N__44066),
            .I(N__44060));
    InMux I__9864 (
            .O(N__44063),
            .I(N__44056));
    Span4Mux_v I__9863 (
            .O(N__44060),
            .I(N__44053));
    CascadeMux I__9862 (
            .O(N__44059),
            .I(N__44050));
    LocalMux I__9861 (
            .O(N__44056),
            .I(N__44047));
    Span4Mux_h I__9860 (
            .O(N__44053),
            .I(N__44044));
    InMux I__9859 (
            .O(N__44050),
            .I(N__44041));
    Span4Mux_h I__9858 (
            .O(N__44047),
            .I(N__44038));
    Span4Mux_h I__9857 (
            .O(N__44044),
            .I(N__44033));
    LocalMux I__9856 (
            .O(N__44041),
            .I(N__44033));
    Span4Mux_v I__9855 (
            .O(N__44038),
            .I(N__44029));
    Span4Mux_h I__9854 (
            .O(N__44033),
            .I(N__44026));
    CascadeMux I__9853 (
            .O(N__44032),
            .I(N__44023));
    Span4Mux_h I__9852 (
            .O(N__44029),
            .I(N__44020));
    Span4Mux_v I__9851 (
            .O(N__44026),
            .I(N__44017));
    InMux I__9850 (
            .O(N__44023),
            .I(N__44014));
    Span4Mux_h I__9849 (
            .O(N__44020),
            .I(N__44011));
    Span4Mux_v I__9848 (
            .O(N__44017),
            .I(N__44008));
    LocalMux I__9847 (
            .O(N__44014),
            .I(trig_dds1));
    Odrv4 I__9846 (
            .O(N__44011),
            .I(trig_dds1));
    Odrv4 I__9845 (
            .O(N__44008),
            .I(trig_dds1));
    InMux I__9844 (
            .O(N__44001),
            .I(N__43997));
    InMux I__9843 (
            .O(N__44000),
            .I(N__43994));
    LocalMux I__9842 (
            .O(N__43997),
            .I(N__43990));
    LocalMux I__9841 (
            .O(N__43994),
            .I(N__43987));
    InMux I__9840 (
            .O(N__43993),
            .I(N__43984));
    Span4Mux_h I__9839 (
            .O(N__43990),
            .I(N__43981));
    Odrv4 I__9838 (
            .O(N__43987),
            .I(buf_dds0_11));
    LocalMux I__9837 (
            .O(N__43984),
            .I(buf_dds0_11));
    Odrv4 I__9836 (
            .O(N__43981),
            .I(buf_dds0_11));
    CascadeMux I__9835 (
            .O(N__43974),
            .I(n22297_cascade_));
    InMux I__9834 (
            .O(N__43971),
            .I(N__43967));
    InMux I__9833 (
            .O(N__43970),
            .I(N__43963));
    LocalMux I__9832 (
            .O(N__43967),
            .I(N__43960));
    InMux I__9831 (
            .O(N__43966),
            .I(N__43957));
    LocalMux I__9830 (
            .O(N__43963),
            .I(N__43954));
    Span12Mux_h I__9829 (
            .O(N__43960),
            .I(N__43951));
    LocalMux I__9828 (
            .O(N__43957),
            .I(N__43946));
    Span4Mux_h I__9827 (
            .O(N__43954),
            .I(N__43946));
    Odrv12 I__9826 (
            .O(N__43951),
            .I(buf_dds1_11));
    Odrv4 I__9825 (
            .O(N__43946),
            .I(buf_dds1_11));
    InMux I__9824 (
            .O(N__43941),
            .I(N__43938));
    LocalMux I__9823 (
            .O(N__43938),
            .I(N__43935));
    Odrv12 I__9822 (
            .O(N__43935),
            .I(n21076));
    CascadeMux I__9821 (
            .O(N__43932),
            .I(N__43929));
    InMux I__9820 (
            .O(N__43929),
            .I(N__43926));
    LocalMux I__9819 (
            .O(N__43926),
            .I(n22300));
    CascadeMux I__9818 (
            .O(N__43923),
            .I(n22312_cascade_));
    CascadeMux I__9817 (
            .O(N__43920),
            .I(N__43917));
    InMux I__9816 (
            .O(N__43917),
            .I(N__43914));
    LocalMux I__9815 (
            .O(N__43914),
            .I(N__43911));
    Span4Mux_h I__9814 (
            .O(N__43911),
            .I(N__43907));
    InMux I__9813 (
            .O(N__43910),
            .I(N__43901));
    Span4Mux_h I__9812 (
            .O(N__43907),
            .I(N__43898));
    InMux I__9811 (
            .O(N__43906),
            .I(N__43895));
    InMux I__9810 (
            .O(N__43905),
            .I(N__43890));
    InMux I__9809 (
            .O(N__43904),
            .I(N__43890));
    LocalMux I__9808 (
            .O(N__43901),
            .I(eis_start));
    Odrv4 I__9807 (
            .O(N__43898),
            .I(eis_start));
    LocalMux I__9806 (
            .O(N__43895),
            .I(eis_start));
    LocalMux I__9805 (
            .O(N__43890),
            .I(eis_start));
    InMux I__9804 (
            .O(N__43881),
            .I(N__43878));
    LocalMux I__9803 (
            .O(N__43878),
            .I(N__43873));
    CascadeMux I__9802 (
            .O(N__43877),
            .I(N__43870));
    InMux I__9801 (
            .O(N__43876),
            .I(N__43867));
    Span4Mux_h I__9800 (
            .O(N__43873),
            .I(N__43864));
    InMux I__9799 (
            .O(N__43870),
            .I(N__43861));
    LocalMux I__9798 (
            .O(N__43867),
            .I(req_data_cnt_8));
    Odrv4 I__9797 (
            .O(N__43864),
            .I(req_data_cnt_8));
    LocalMux I__9796 (
            .O(N__43861),
            .I(req_data_cnt_8));
    InMux I__9795 (
            .O(N__43854),
            .I(N__43851));
    LocalMux I__9794 (
            .O(N__43851),
            .I(N__43848));
    Span4Mux_h I__9793 (
            .O(N__43848),
            .I(N__43845));
    Span4Mux_h I__9792 (
            .O(N__43845),
            .I(N__43842));
    Odrv4 I__9791 (
            .O(N__43842),
            .I(n22294));
    CascadeMux I__9790 (
            .O(N__43839),
            .I(n21071_cascade_));
    CascadeMux I__9789 (
            .O(N__43836),
            .I(N__43832));
    CascadeMux I__9788 (
            .O(N__43835),
            .I(N__43826));
    InMux I__9787 (
            .O(N__43832),
            .I(N__43819));
    InMux I__9786 (
            .O(N__43831),
            .I(N__43819));
    InMux I__9785 (
            .O(N__43830),
            .I(N__43816));
    CascadeMux I__9784 (
            .O(N__43829),
            .I(N__43812));
    InMux I__9783 (
            .O(N__43826),
            .I(N__43809));
    InMux I__9782 (
            .O(N__43825),
            .I(N__43805));
    InMux I__9781 (
            .O(N__43824),
            .I(N__43802));
    LocalMux I__9780 (
            .O(N__43819),
            .I(N__43799));
    LocalMux I__9779 (
            .O(N__43816),
            .I(N__43796));
    InMux I__9778 (
            .O(N__43815),
            .I(N__43793));
    InMux I__9777 (
            .O(N__43812),
            .I(N__43790));
    LocalMux I__9776 (
            .O(N__43809),
            .I(N__43787));
    CascadeMux I__9775 (
            .O(N__43808),
            .I(N__43784));
    LocalMux I__9774 (
            .O(N__43805),
            .I(N__43780));
    LocalMux I__9773 (
            .O(N__43802),
            .I(N__43775));
    Span4Mux_v I__9772 (
            .O(N__43799),
            .I(N__43775));
    Span4Mux_v I__9771 (
            .O(N__43796),
            .I(N__43770));
    LocalMux I__9770 (
            .O(N__43793),
            .I(N__43770));
    LocalMux I__9769 (
            .O(N__43790),
            .I(N__43767));
    Span4Mux_h I__9768 (
            .O(N__43787),
            .I(N__43764));
    InMux I__9767 (
            .O(N__43784),
            .I(N__43761));
    InMux I__9766 (
            .O(N__43783),
            .I(N__43758));
    Span4Mux_v I__9765 (
            .O(N__43780),
            .I(N__43755));
    Span4Mux_h I__9764 (
            .O(N__43775),
            .I(N__43750));
    Span4Mux_h I__9763 (
            .O(N__43770),
            .I(N__43750));
    Span4Mux_h I__9762 (
            .O(N__43767),
            .I(N__43745));
    Span4Mux_v I__9761 (
            .O(N__43764),
            .I(N__43745));
    LocalMux I__9760 (
            .O(N__43761),
            .I(N__43740));
    LocalMux I__9759 (
            .O(N__43758),
            .I(N__43740));
    Span4Mux_v I__9758 (
            .O(N__43755),
            .I(N__43735));
    Span4Mux_h I__9757 (
            .O(N__43750),
            .I(N__43735));
    Span4Mux_h I__9756 (
            .O(N__43745),
            .I(N__43730));
    Span4Mux_v I__9755 (
            .O(N__43740),
            .I(N__43730));
    Odrv4 I__9754 (
            .O(N__43735),
            .I(comm_buf_0_0));
    Odrv4 I__9753 (
            .O(N__43730),
            .I(comm_buf_0_0));
    SRMux I__9752 (
            .O(N__43725),
            .I(N__43720));
    SRMux I__9751 (
            .O(N__43724),
            .I(N__43717));
    SRMux I__9750 (
            .O(N__43723),
            .I(N__43714));
    LocalMux I__9749 (
            .O(N__43720),
            .I(N__43711));
    LocalMux I__9748 (
            .O(N__43717),
            .I(N__43707));
    LocalMux I__9747 (
            .O(N__43714),
            .I(N__43704));
    Span4Mux_h I__9746 (
            .O(N__43711),
            .I(N__43701));
    SRMux I__9745 (
            .O(N__43710),
            .I(N__43695));
    Span4Mux_v I__9744 (
            .O(N__43707),
            .I(N__43690));
    Span4Mux_v I__9743 (
            .O(N__43704),
            .I(N__43690));
    Span4Mux_h I__9742 (
            .O(N__43701),
            .I(N__43687));
    SRMux I__9741 (
            .O(N__43700),
            .I(N__43684));
    SRMux I__9740 (
            .O(N__43699),
            .I(N__43681));
    SRMux I__9739 (
            .O(N__43698),
            .I(N__43678));
    LocalMux I__9738 (
            .O(N__43695),
            .I(N__43675));
    Sp12to4 I__9737 (
            .O(N__43690),
            .I(N__43672));
    Span4Mux_v I__9736 (
            .O(N__43687),
            .I(N__43669));
    LocalMux I__9735 (
            .O(N__43684),
            .I(n14750));
    LocalMux I__9734 (
            .O(N__43681),
            .I(n14750));
    LocalMux I__9733 (
            .O(N__43678),
            .I(n14750));
    Odrv12 I__9732 (
            .O(N__43675),
            .I(n14750));
    Odrv12 I__9731 (
            .O(N__43672),
            .I(n14750));
    Odrv4 I__9730 (
            .O(N__43669),
            .I(n14750));
    InMux I__9729 (
            .O(N__43656),
            .I(N__43653));
    LocalMux I__9728 (
            .O(N__43653),
            .I(n22219));
    InMux I__9727 (
            .O(N__43650),
            .I(N__43646));
    InMux I__9726 (
            .O(N__43649),
            .I(N__43643));
    LocalMux I__9725 (
            .O(N__43646),
            .I(N__43640));
    LocalMux I__9724 (
            .O(N__43643),
            .I(N__43636));
    Span12Mux_h I__9723 (
            .O(N__43640),
            .I(N__43633));
    InMux I__9722 (
            .O(N__43639),
            .I(N__43630));
    Odrv4 I__9721 (
            .O(N__43636),
            .I(acadc_skipCount_8));
    Odrv12 I__9720 (
            .O(N__43633),
            .I(acadc_skipCount_8));
    LocalMux I__9719 (
            .O(N__43630),
            .I(acadc_skipCount_8));
    InMux I__9718 (
            .O(N__43623),
            .I(N__43620));
    LocalMux I__9717 (
            .O(N__43620),
            .I(N__43617));
    Span4Mux_v I__9716 (
            .O(N__43617),
            .I(N__43614));
    Span4Mux_h I__9715 (
            .O(N__43614),
            .I(N__43611));
    Span4Mux_h I__9714 (
            .O(N__43611),
            .I(N__43608));
    Odrv4 I__9713 (
            .O(N__43608),
            .I(n22324));
    CascadeMux I__9712 (
            .O(N__43605),
            .I(N__43602));
    InMux I__9711 (
            .O(N__43602),
            .I(N__43597));
    CascadeMux I__9710 (
            .O(N__43601),
            .I(N__43594));
    CascadeMux I__9709 (
            .O(N__43600),
            .I(N__43590));
    LocalMux I__9708 (
            .O(N__43597),
            .I(N__43586));
    InMux I__9707 (
            .O(N__43594),
            .I(N__43583));
    InMux I__9706 (
            .O(N__43593),
            .I(N__43580));
    InMux I__9705 (
            .O(N__43590),
            .I(N__43577));
    InMux I__9704 (
            .O(N__43589),
            .I(N__43574));
    Span4Mux_v I__9703 (
            .O(N__43586),
            .I(N__43569));
    LocalMux I__9702 (
            .O(N__43583),
            .I(N__43569));
    LocalMux I__9701 (
            .O(N__43580),
            .I(N__43564));
    LocalMux I__9700 (
            .O(N__43577),
            .I(N__43561));
    LocalMux I__9699 (
            .O(N__43574),
            .I(N__43556));
    Span4Mux_h I__9698 (
            .O(N__43569),
            .I(N__43556));
    InMux I__9697 (
            .O(N__43568),
            .I(N__43553));
    InMux I__9696 (
            .O(N__43567),
            .I(N__43550));
    Span4Mux_v I__9695 (
            .O(N__43564),
            .I(N__43547));
    Span12Mux_v I__9694 (
            .O(N__43561),
            .I(N__43544));
    Sp12to4 I__9693 (
            .O(N__43556),
            .I(N__43539));
    LocalMux I__9692 (
            .O(N__43553),
            .I(N__43539));
    LocalMux I__9691 (
            .O(N__43550),
            .I(N__43536));
    Sp12to4 I__9690 (
            .O(N__43547),
            .I(N__43531));
    Span12Mux_h I__9689 (
            .O(N__43544),
            .I(N__43531));
    Span12Mux_v I__9688 (
            .O(N__43539),
            .I(N__43528));
    Odrv4 I__9687 (
            .O(N__43536),
            .I(comm_buf_0_5));
    Odrv12 I__9686 (
            .O(N__43531),
            .I(comm_buf_0_5));
    Odrv12 I__9685 (
            .O(N__43528),
            .I(comm_buf_0_5));
    CascadeMux I__9684 (
            .O(N__43521),
            .I(N__43518));
    InMux I__9683 (
            .O(N__43518),
            .I(N__43514));
    InMux I__9682 (
            .O(N__43517),
            .I(N__43511));
    LocalMux I__9681 (
            .O(N__43514),
            .I(N__43508));
    LocalMux I__9680 (
            .O(N__43511),
            .I(N__43505));
    Span4Mux_v I__9679 (
            .O(N__43508),
            .I(N__43499));
    Span4Mux_v I__9678 (
            .O(N__43505),
            .I(N__43499));
    CascadeMux I__9677 (
            .O(N__43504),
            .I(N__43496));
    Sp12to4 I__9676 (
            .O(N__43499),
            .I(N__43493));
    InMux I__9675 (
            .O(N__43496),
            .I(N__43490));
    Span12Mux_h I__9674 (
            .O(N__43493),
            .I(N__43487));
    LocalMux I__9673 (
            .O(N__43490),
            .I(buf_adcdata_iac_8));
    Odrv12 I__9672 (
            .O(N__43487),
            .I(buf_adcdata_iac_8));
    InMux I__9671 (
            .O(N__43482),
            .I(N__43479));
    LocalMux I__9670 (
            .O(N__43479),
            .I(N__43476));
    Span4Mux_v I__9669 (
            .O(N__43476),
            .I(N__43473));
    Span4Mux_h I__9668 (
            .O(N__43473),
            .I(N__43470));
    Odrv4 I__9667 (
            .O(N__43470),
            .I(n16_adj_1487));
    InMux I__9666 (
            .O(N__43467),
            .I(N__43464));
    LocalMux I__9665 (
            .O(N__43464),
            .I(N__43461));
    Span4Mux_h I__9664 (
            .O(N__43461),
            .I(N__43458));
    Span4Mux_h I__9663 (
            .O(N__43458),
            .I(N__43455));
    Span4Mux_h I__9662 (
            .O(N__43455),
            .I(N__43452));
    Odrv4 I__9661 (
            .O(N__43452),
            .I(n19_adj_1486));
    CascadeMux I__9660 (
            .O(N__43449),
            .I(N__43446));
    InMux I__9659 (
            .O(N__43446),
            .I(N__43443));
    LocalMux I__9658 (
            .O(N__43443),
            .I(N__43440));
    Span12Mux_v I__9657 (
            .O(N__43440),
            .I(N__43436));
    CascadeMux I__9656 (
            .O(N__43439),
            .I(N__43433));
    Span12Mux_h I__9655 (
            .O(N__43436),
            .I(N__43430));
    InMux I__9654 (
            .O(N__43433),
            .I(N__43427));
    Odrv12 I__9653 (
            .O(N__43430),
            .I(buf_readRTD_0));
    LocalMux I__9652 (
            .O(N__43427),
            .I(buf_readRTD_0));
    InMux I__9651 (
            .O(N__43422),
            .I(N__43419));
    LocalMux I__9650 (
            .O(N__43419),
            .I(n22213));
    InMux I__9649 (
            .O(N__43416),
            .I(N__43413));
    LocalMux I__9648 (
            .O(N__43413),
            .I(N__43409));
    CascadeMux I__9647 (
            .O(N__43412),
            .I(N__43406));
    Span4Mux_v I__9646 (
            .O(N__43409),
            .I(N__43403));
    InMux I__9645 (
            .O(N__43406),
            .I(N__43400));
    Span4Mux_h I__9644 (
            .O(N__43403),
            .I(N__43397));
    LocalMux I__9643 (
            .O(N__43400),
            .I(data_idxvec_0));
    Odrv4 I__9642 (
            .O(N__43397),
            .I(data_idxvec_0));
    InMux I__9641 (
            .O(N__43392),
            .I(N__43388));
    InMux I__9640 (
            .O(N__43391),
            .I(N__43384));
    LocalMux I__9639 (
            .O(N__43388),
            .I(N__43381));
    InMux I__9638 (
            .O(N__43387),
            .I(N__43378));
    LocalMux I__9637 (
            .O(N__43384),
            .I(N__43373));
    Span4Mux_h I__9636 (
            .O(N__43381),
            .I(N__43373));
    LocalMux I__9635 (
            .O(N__43378),
            .I(data_cntvec_0));
    Odrv4 I__9634 (
            .O(N__43373),
            .I(data_cntvec_0));
    CascadeMux I__9633 (
            .O(N__43368),
            .I(n26_cascade_));
    InMux I__9632 (
            .O(N__43365),
            .I(N__43362));
    LocalMux I__9631 (
            .O(N__43362),
            .I(N__43358));
    InMux I__9630 (
            .O(N__43361),
            .I(N__43354));
    Span4Mux_v I__9629 (
            .O(N__43358),
            .I(N__43351));
    InMux I__9628 (
            .O(N__43357),
            .I(N__43348));
    LocalMux I__9627 (
            .O(N__43354),
            .I(acadc_skipCount_0));
    Odrv4 I__9626 (
            .O(N__43351),
            .I(acadc_skipCount_0));
    LocalMux I__9625 (
            .O(N__43348),
            .I(acadc_skipCount_0));
    CascadeMux I__9624 (
            .O(N__43341),
            .I(n22201_cascade_));
    InMux I__9623 (
            .O(N__43338),
            .I(N__43335));
    LocalMux I__9622 (
            .O(N__43335),
            .I(N__43330));
    CascadeMux I__9621 (
            .O(N__43334),
            .I(N__43327));
    CascadeMux I__9620 (
            .O(N__43333),
            .I(N__43324));
    Span4Mux_v I__9619 (
            .O(N__43330),
            .I(N__43321));
    InMux I__9618 (
            .O(N__43327),
            .I(N__43316));
    InMux I__9617 (
            .O(N__43324),
            .I(N__43316));
    Odrv4 I__9616 (
            .O(N__43321),
            .I(req_data_cnt_0));
    LocalMux I__9615 (
            .O(N__43316),
            .I(req_data_cnt_0));
    InMux I__9614 (
            .O(N__43311),
            .I(N__43308));
    LocalMux I__9613 (
            .O(N__43308),
            .I(n22216));
    CascadeMux I__9612 (
            .O(N__43305),
            .I(n22204_cascade_));
    CascadeMux I__9611 (
            .O(N__43302),
            .I(n30_adj_1485_cascade_));
    CascadeMux I__9610 (
            .O(N__43299),
            .I(N__43296));
    InMux I__9609 (
            .O(N__43296),
            .I(N__43293));
    LocalMux I__9608 (
            .O(N__43293),
            .I(N__43287));
    InMux I__9607 (
            .O(N__43292),
            .I(N__43284));
    InMux I__9606 (
            .O(N__43291),
            .I(N__43279));
    InMux I__9605 (
            .O(N__43290),
            .I(N__43276));
    Span4Mux_v I__9604 (
            .O(N__43287),
            .I(N__43271));
    LocalMux I__9603 (
            .O(N__43284),
            .I(N__43271));
    InMux I__9602 (
            .O(N__43283),
            .I(N__43268));
    InMux I__9601 (
            .O(N__43282),
            .I(N__43265));
    LocalMux I__9600 (
            .O(N__43279),
            .I(N__43262));
    LocalMux I__9599 (
            .O(N__43276),
            .I(N__43259));
    Span4Mux_v I__9598 (
            .O(N__43271),
            .I(N__43254));
    LocalMux I__9597 (
            .O(N__43268),
            .I(N__43254));
    LocalMux I__9596 (
            .O(N__43265),
            .I(N__43251));
    Span4Mux_h I__9595 (
            .O(N__43262),
            .I(N__43248));
    Span4Mux_v I__9594 (
            .O(N__43259),
            .I(N__43243));
    Span4Mux_v I__9593 (
            .O(N__43254),
            .I(N__43243));
    Span4Mux_v I__9592 (
            .O(N__43251),
            .I(N__43240));
    Span4Mux_v I__9591 (
            .O(N__43248),
            .I(N__43235));
    Span4Mux_h I__9590 (
            .O(N__43243),
            .I(N__43235));
    Odrv4 I__9589 (
            .O(N__43240),
            .I(comm_buf_1_0));
    Odrv4 I__9588 (
            .O(N__43235),
            .I(comm_buf_1_0));
    InMux I__9587 (
            .O(N__43230),
            .I(N__43226));
    CascadeMux I__9586 (
            .O(N__43229),
            .I(N__43223));
    LocalMux I__9585 (
            .O(N__43226),
            .I(N__43220));
    InMux I__9584 (
            .O(N__43223),
            .I(N__43217));
    Span12Mux_v I__9583 (
            .O(N__43220),
            .I(N__43213));
    LocalMux I__9582 (
            .O(N__43217),
            .I(N__43210));
    InMux I__9581 (
            .O(N__43216),
            .I(N__43207));
    Span12Mux_h I__9580 (
            .O(N__43213),
            .I(N__43204));
    Span12Mux_v I__9579 (
            .O(N__43210),
            .I(N__43201));
    LocalMux I__9578 (
            .O(N__43207),
            .I(buf_adcdata_iac_19));
    Odrv12 I__9577 (
            .O(N__43204),
            .I(buf_adcdata_iac_19));
    Odrv12 I__9576 (
            .O(N__43201),
            .I(buf_adcdata_iac_19));
    InMux I__9575 (
            .O(N__43194),
            .I(N__43191));
    LocalMux I__9574 (
            .O(N__43191),
            .I(comm_buf_4_1));
    InMux I__9573 (
            .O(N__43188),
            .I(N__43185));
    LocalMux I__9572 (
            .O(N__43185),
            .I(N__43181));
    InMux I__9571 (
            .O(N__43184),
            .I(N__43178));
    Span4Mux_h I__9570 (
            .O(N__43181),
            .I(N__43175));
    LocalMux I__9569 (
            .O(N__43178),
            .I(\SIG_DDS.bit_cnt_3 ));
    Odrv4 I__9568 (
            .O(N__43175),
            .I(\SIG_DDS.bit_cnt_3 ));
    InMux I__9567 (
            .O(N__43170),
            .I(N__43161));
    InMux I__9566 (
            .O(N__43169),
            .I(N__43161));
    InMux I__9565 (
            .O(N__43168),
            .I(N__43161));
    LocalMux I__9564 (
            .O(N__43161),
            .I(N__43158));
    Span4Mux_v I__9563 (
            .O(N__43158),
            .I(N__43154));
    InMux I__9562 (
            .O(N__43157),
            .I(N__43151));
    Span4Mux_h I__9561 (
            .O(N__43154),
            .I(N__43147));
    LocalMux I__9560 (
            .O(N__43151),
            .I(N__43144));
    InMux I__9559 (
            .O(N__43150),
            .I(N__43141));
    Odrv4 I__9558 (
            .O(N__43147),
            .I(bit_cnt_0));
    Odrv4 I__9557 (
            .O(N__43144),
            .I(bit_cnt_0));
    LocalMux I__9556 (
            .O(N__43141),
            .I(bit_cnt_0));
    InMux I__9555 (
            .O(N__43134),
            .I(N__43131));
    LocalMux I__9554 (
            .O(N__43131),
            .I(N__43128));
    Span4Mux_v I__9553 (
            .O(N__43128),
            .I(N__43123));
    CascadeMux I__9552 (
            .O(N__43127),
            .I(N__43120));
    CascadeMux I__9551 (
            .O(N__43126),
            .I(N__43117));
    Sp12to4 I__9550 (
            .O(N__43123),
            .I(N__43113));
    InMux I__9549 (
            .O(N__43120),
            .I(N__43106));
    InMux I__9548 (
            .O(N__43117),
            .I(N__43106));
    InMux I__9547 (
            .O(N__43116),
            .I(N__43106));
    Span12Mux_v I__9546 (
            .O(N__43113),
            .I(N__43103));
    LocalMux I__9545 (
            .O(N__43106),
            .I(\SIG_DDS.bit_cnt_1 ));
    Odrv12 I__9544 (
            .O(N__43103),
            .I(\SIG_DDS.bit_cnt_1 ));
    CascadeMux I__9543 (
            .O(N__43098),
            .I(N__43095));
    InMux I__9542 (
            .O(N__43095),
            .I(N__43092));
    LocalMux I__9541 (
            .O(N__43092),
            .I(N__43087));
    InMux I__9540 (
            .O(N__43091),
            .I(N__43082));
    InMux I__9539 (
            .O(N__43090),
            .I(N__43082));
    Span12Mux_h I__9538 (
            .O(N__43087),
            .I(N__43079));
    LocalMux I__9537 (
            .O(N__43082),
            .I(\SIG_DDS.bit_cnt_2 ));
    Odrv12 I__9536 (
            .O(N__43079),
            .I(\SIG_DDS.bit_cnt_2 ));
    CEMux I__9535 (
            .O(N__43074),
            .I(N__43071));
    LocalMux I__9534 (
            .O(N__43071),
            .I(N__43056));
    InMux I__9533 (
            .O(N__43070),
            .I(N__43053));
    InMux I__9532 (
            .O(N__43069),
            .I(N__43027));
    InMux I__9531 (
            .O(N__43068),
            .I(N__43027));
    InMux I__9530 (
            .O(N__43067),
            .I(N__43027));
    InMux I__9529 (
            .O(N__43066),
            .I(N__43027));
    InMux I__9528 (
            .O(N__43065),
            .I(N__43027));
    InMux I__9527 (
            .O(N__43064),
            .I(N__43027));
    InMux I__9526 (
            .O(N__43063),
            .I(N__43027));
    InMux I__9525 (
            .O(N__43062),
            .I(N__43027));
    InMux I__9524 (
            .O(N__43061),
            .I(N__43024));
    SRMux I__9523 (
            .O(N__43060),
            .I(N__43021));
    CascadeMux I__9522 (
            .O(N__43059),
            .I(N__43017));
    Span4Mux_v I__9521 (
            .O(N__43056),
            .I(N__43014));
    LocalMux I__9520 (
            .O(N__43053),
            .I(N__43011));
    InMux I__9519 (
            .O(N__43052),
            .I(N__43006));
    InMux I__9518 (
            .O(N__43051),
            .I(N__43006));
    InMux I__9517 (
            .O(N__43050),
            .I(N__42993));
    InMux I__9516 (
            .O(N__43049),
            .I(N__42993));
    InMux I__9515 (
            .O(N__43048),
            .I(N__42993));
    InMux I__9514 (
            .O(N__43047),
            .I(N__42993));
    InMux I__9513 (
            .O(N__43046),
            .I(N__42993));
    InMux I__9512 (
            .O(N__43045),
            .I(N__42993));
    InMux I__9511 (
            .O(N__43044),
            .I(N__42990));
    LocalMux I__9510 (
            .O(N__43027),
            .I(N__42987));
    LocalMux I__9509 (
            .O(N__43024),
            .I(N__42984));
    LocalMux I__9508 (
            .O(N__43021),
            .I(N__42980));
    InMux I__9507 (
            .O(N__43020),
            .I(N__42977));
    InMux I__9506 (
            .O(N__43017),
            .I(N__42973));
    Span4Mux_h I__9505 (
            .O(N__43014),
            .I(N__42968));
    Span4Mux_h I__9504 (
            .O(N__43011),
            .I(N__42968));
    LocalMux I__9503 (
            .O(N__43006),
            .I(N__42965));
    LocalMux I__9502 (
            .O(N__42993),
            .I(N__42962));
    LocalMux I__9501 (
            .O(N__42990),
            .I(N__42959));
    Span4Mux_v I__9500 (
            .O(N__42987),
            .I(N__42953));
    Span4Mux_h I__9499 (
            .O(N__42984),
            .I(N__42950));
    InMux I__9498 (
            .O(N__42983),
            .I(N__42947));
    Span4Mux_h I__9497 (
            .O(N__42980),
            .I(N__42944));
    LocalMux I__9496 (
            .O(N__42977),
            .I(N__42941));
    InMux I__9495 (
            .O(N__42976),
            .I(N__42938));
    LocalMux I__9494 (
            .O(N__42973),
            .I(N__42933));
    Span4Mux_v I__9493 (
            .O(N__42968),
            .I(N__42933));
    Span4Mux_v I__9492 (
            .O(N__42965),
            .I(N__42930));
    Span4Mux_v I__9491 (
            .O(N__42962),
            .I(N__42925));
    Span4Mux_v I__9490 (
            .O(N__42959),
            .I(N__42925));
    InMux I__9489 (
            .O(N__42958),
            .I(N__42918));
    InMux I__9488 (
            .O(N__42957),
            .I(N__42918));
    InMux I__9487 (
            .O(N__42956),
            .I(N__42918));
    Span4Mux_v I__9486 (
            .O(N__42953),
            .I(N__42915));
    Sp12to4 I__9485 (
            .O(N__42950),
            .I(N__42912));
    LocalMux I__9484 (
            .O(N__42947),
            .I(N__42905));
    Span4Mux_h I__9483 (
            .O(N__42944),
            .I(N__42905));
    Span4Mux_v I__9482 (
            .O(N__42941),
            .I(N__42905));
    LocalMux I__9481 (
            .O(N__42938),
            .I(N__42900));
    Span4Mux_v I__9480 (
            .O(N__42933),
            .I(N__42900));
    Odrv4 I__9479 (
            .O(N__42930),
            .I(dds_state_1));
    Odrv4 I__9478 (
            .O(N__42925),
            .I(dds_state_1));
    LocalMux I__9477 (
            .O(N__42918),
            .I(dds_state_1));
    Odrv4 I__9476 (
            .O(N__42915),
            .I(dds_state_1));
    Odrv12 I__9475 (
            .O(N__42912),
            .I(dds_state_1));
    Odrv4 I__9474 (
            .O(N__42905),
            .I(dds_state_1));
    Odrv4 I__9473 (
            .O(N__42900),
            .I(dds_state_1));
    SRMux I__9472 (
            .O(N__42885),
            .I(N__42882));
    LocalMux I__9471 (
            .O(N__42882),
            .I(N__42878));
    InMux I__9470 (
            .O(N__42881),
            .I(N__42875));
    Span4Mux_v I__9469 (
            .O(N__42878),
            .I(N__42872));
    LocalMux I__9468 (
            .O(N__42875),
            .I(N__42869));
    Span4Mux_h I__9467 (
            .O(N__42872),
            .I(N__42866));
    Span4Mux_v I__9466 (
            .O(N__42869),
            .I(N__42863));
    Odrv4 I__9465 (
            .O(N__42866),
            .I(n14884));
    Odrv4 I__9464 (
            .O(N__42863),
            .I(n14884));
    CEMux I__9463 (
            .O(N__42858),
            .I(N__42855));
    LocalMux I__9462 (
            .O(N__42855),
            .I(n12220));
    CascadeMux I__9461 (
            .O(N__42852),
            .I(n12220_cascade_));
    SRMux I__9460 (
            .O(N__42849),
            .I(N__42846));
    LocalMux I__9459 (
            .O(N__42846),
            .I(n14785));
    SRMux I__9458 (
            .O(N__42843),
            .I(N__42840));
    LocalMux I__9457 (
            .O(N__42840),
            .I(N__42837));
    Span4Mux_h I__9456 (
            .O(N__42837),
            .I(N__42834));
    Odrv4 I__9455 (
            .O(N__42834),
            .I(n14778));
    InMux I__9454 (
            .O(N__42831),
            .I(N__42828));
    LocalMux I__9453 (
            .O(N__42828),
            .I(N__42825));
    Span4Mux_v I__9452 (
            .O(N__42825),
            .I(N__42822));
    Span4Mux_h I__9451 (
            .O(N__42822),
            .I(N__42819));
    Odrv4 I__9450 (
            .O(N__42819),
            .I(n30_adj_1531));
    CascadeMux I__9449 (
            .O(N__42816),
            .I(N__42811));
    CascadeMux I__9448 (
            .O(N__42815),
            .I(N__42807));
    CascadeMux I__9447 (
            .O(N__42814),
            .I(N__42804));
    InMux I__9446 (
            .O(N__42811),
            .I(N__42799));
    InMux I__9445 (
            .O(N__42810),
            .I(N__42794));
    InMux I__9444 (
            .O(N__42807),
            .I(N__42794));
    InMux I__9443 (
            .O(N__42804),
            .I(N__42791));
    InMux I__9442 (
            .O(N__42803),
            .I(N__42788));
    InMux I__9441 (
            .O(N__42802),
            .I(N__42785));
    LocalMux I__9440 (
            .O(N__42799),
            .I(N__42782));
    LocalMux I__9439 (
            .O(N__42794),
            .I(N__42777));
    LocalMux I__9438 (
            .O(N__42791),
            .I(N__42777));
    LocalMux I__9437 (
            .O(N__42788),
            .I(N__42774));
    LocalMux I__9436 (
            .O(N__42785),
            .I(N__42771));
    Span4Mux_h I__9435 (
            .O(N__42782),
            .I(N__42767));
    Span4Mux_v I__9434 (
            .O(N__42777),
            .I(N__42762));
    Span4Mux_v I__9433 (
            .O(N__42774),
            .I(N__42762));
    Span4Mux_h I__9432 (
            .O(N__42771),
            .I(N__42759));
    InMux I__9431 (
            .O(N__42770),
            .I(N__42756));
    Span4Mux_h I__9430 (
            .O(N__42767),
            .I(N__42753));
    Span4Mux_h I__9429 (
            .O(N__42762),
            .I(N__42746));
    Span4Mux_v I__9428 (
            .O(N__42759),
            .I(N__42746));
    LocalMux I__9427 (
            .O(N__42756),
            .I(N__42746));
    Span4Mux_v I__9426 (
            .O(N__42753),
            .I(N__42743));
    Span4Mux_h I__9425 (
            .O(N__42746),
            .I(N__42740));
    Odrv4 I__9424 (
            .O(N__42743),
            .I(comm_buf_0_7));
    Odrv4 I__9423 (
            .O(N__42740),
            .I(comm_buf_0_7));
    InMux I__9422 (
            .O(N__42735),
            .I(N__42729));
    InMux I__9421 (
            .O(N__42734),
            .I(N__42729));
    LocalMux I__9420 (
            .O(N__42729),
            .I(N__42725));
    InMux I__9419 (
            .O(N__42728),
            .I(N__42722));
    Odrv12 I__9418 (
            .O(N__42725),
            .I(comm_tx_buf_5));
    LocalMux I__9417 (
            .O(N__42722),
            .I(comm_tx_buf_5));
    InMux I__9416 (
            .O(N__42717),
            .I(N__42714));
    LocalMux I__9415 (
            .O(N__42714),
            .I(N__42711));
    Span4Mux_h I__9414 (
            .O(N__42711),
            .I(N__42708));
    Span4Mux_v I__9413 (
            .O(N__42708),
            .I(N__42705));
    Span4Mux_v I__9412 (
            .O(N__42705),
            .I(N__42702));
    Odrv4 I__9411 (
            .O(N__42702),
            .I(buf_data_vac_8));
    InMux I__9410 (
            .O(N__42699),
            .I(N__42696));
    LocalMux I__9409 (
            .O(N__42696),
            .I(N__42693));
    Odrv4 I__9408 (
            .O(N__42693),
            .I(comm_buf_4_0));
    InMux I__9407 (
            .O(N__42690),
            .I(N__42687));
    LocalMux I__9406 (
            .O(N__42687),
            .I(N__42684));
    Span4Mux_h I__9405 (
            .O(N__42684),
            .I(N__42681));
    Span4Mux_h I__9404 (
            .O(N__42681),
            .I(N__42678));
    Odrv4 I__9403 (
            .O(N__42678),
            .I(buf_data_vac_15));
    InMux I__9402 (
            .O(N__42675),
            .I(N__42672));
    LocalMux I__9401 (
            .O(N__42672),
            .I(N__42669));
    Span4Mux_v I__9400 (
            .O(N__42669),
            .I(N__42666));
    Span4Mux_h I__9399 (
            .O(N__42666),
            .I(N__42663));
    Odrv4 I__9398 (
            .O(N__42663),
            .I(comm_buf_4_7));
    InMux I__9397 (
            .O(N__42660),
            .I(N__42657));
    LocalMux I__9396 (
            .O(N__42657),
            .I(N__42654));
    Span4Mux_v I__9395 (
            .O(N__42654),
            .I(N__42651));
    Span4Mux_v I__9394 (
            .O(N__42651),
            .I(N__42648));
    Odrv4 I__9393 (
            .O(N__42648),
            .I(buf_data_vac_14));
    InMux I__9392 (
            .O(N__42645),
            .I(N__42642));
    LocalMux I__9391 (
            .O(N__42642),
            .I(N__42639));
    Odrv4 I__9390 (
            .O(N__42639),
            .I(comm_buf_4_6));
    InMux I__9389 (
            .O(N__42636),
            .I(N__42633));
    LocalMux I__9388 (
            .O(N__42633),
            .I(N__42630));
    Span4Mux_h I__9387 (
            .O(N__42630),
            .I(N__42627));
    Span4Mux_v I__9386 (
            .O(N__42627),
            .I(N__42624));
    Odrv4 I__9385 (
            .O(N__42624),
            .I(buf_data_vac_13));
    InMux I__9384 (
            .O(N__42621),
            .I(N__42618));
    LocalMux I__9383 (
            .O(N__42618),
            .I(comm_buf_4_5));
    InMux I__9382 (
            .O(N__42615),
            .I(N__42612));
    LocalMux I__9381 (
            .O(N__42612),
            .I(N__42609));
    Span12Mux_h I__9380 (
            .O(N__42609),
            .I(N__42606));
    Odrv12 I__9379 (
            .O(N__42606),
            .I(buf_data_vac_12));
    InMux I__9378 (
            .O(N__42603),
            .I(N__42600));
    LocalMux I__9377 (
            .O(N__42600),
            .I(N__42597));
    Span4Mux_h I__9376 (
            .O(N__42597),
            .I(N__42594));
    Odrv4 I__9375 (
            .O(N__42594),
            .I(comm_buf_4_4));
    InMux I__9374 (
            .O(N__42591),
            .I(N__42588));
    LocalMux I__9373 (
            .O(N__42588),
            .I(N__42585));
    Span4Mux_h I__9372 (
            .O(N__42585),
            .I(N__42582));
    Span4Mux_v I__9371 (
            .O(N__42582),
            .I(N__42579));
    Odrv4 I__9370 (
            .O(N__42579),
            .I(buf_data_vac_11));
    InMux I__9369 (
            .O(N__42576),
            .I(N__42573));
    LocalMux I__9368 (
            .O(N__42573),
            .I(N__42570));
    Span4Mux_h I__9367 (
            .O(N__42570),
            .I(N__42567));
    Odrv4 I__9366 (
            .O(N__42567),
            .I(comm_buf_4_3));
    InMux I__9365 (
            .O(N__42564),
            .I(N__42561));
    LocalMux I__9364 (
            .O(N__42561),
            .I(N__42558));
    Span4Mux_h I__9363 (
            .O(N__42558),
            .I(N__42555));
    Span4Mux_v I__9362 (
            .O(N__42555),
            .I(N__42552));
    Span4Mux_v I__9361 (
            .O(N__42552),
            .I(N__42549));
    Odrv4 I__9360 (
            .O(N__42549),
            .I(buf_data_vac_10));
    InMux I__9359 (
            .O(N__42546),
            .I(N__42543));
    LocalMux I__9358 (
            .O(N__42543),
            .I(comm_buf_4_2));
    InMux I__9357 (
            .O(N__42540),
            .I(N__42537));
    LocalMux I__9356 (
            .O(N__42537),
            .I(N__42534));
    Span4Mux_v I__9355 (
            .O(N__42534),
            .I(N__42531));
    Span4Mux_h I__9354 (
            .O(N__42531),
            .I(N__42528));
    Span4Mux_v I__9353 (
            .O(N__42528),
            .I(N__42525));
    Odrv4 I__9352 (
            .O(N__42525),
            .I(buf_data_vac_9));
    InMux I__9351 (
            .O(N__42522),
            .I(N__42519));
    LocalMux I__9350 (
            .O(N__42519),
            .I(N__42516));
    Odrv4 I__9349 (
            .O(N__42516),
            .I(n1));
    InMux I__9348 (
            .O(N__42513),
            .I(N__42510));
    LocalMux I__9347 (
            .O(N__42510),
            .I(N__42507));
    Span4Mux_h I__9346 (
            .O(N__42507),
            .I(N__42504));
    Odrv4 I__9345 (
            .O(N__42504),
            .I(comm_buf_2_0));
    InMux I__9344 (
            .O(N__42501),
            .I(N__42498));
    LocalMux I__9343 (
            .O(N__42498),
            .I(n2));
    InMux I__9342 (
            .O(N__42495),
            .I(N__42491));
    InMux I__9341 (
            .O(N__42494),
            .I(N__42488));
    LocalMux I__9340 (
            .O(N__42491),
            .I(N__42485));
    LocalMux I__9339 (
            .O(N__42488),
            .I(N__42482));
    Span4Mux_h I__9338 (
            .O(N__42485),
            .I(N__42478));
    Span4Mux_v I__9337 (
            .O(N__42482),
            .I(N__42475));
    InMux I__9336 (
            .O(N__42481),
            .I(N__42472));
    Odrv4 I__9335 (
            .O(N__42478),
            .I(comm_tx_buf_0));
    Odrv4 I__9334 (
            .O(N__42475),
            .I(comm_tx_buf_0));
    LocalMux I__9333 (
            .O(N__42472),
            .I(comm_tx_buf_0));
    SRMux I__9332 (
            .O(N__42465),
            .I(N__42462));
    LocalMux I__9331 (
            .O(N__42462),
            .I(N__42459));
    Span4Mux_h I__9330 (
            .O(N__42459),
            .I(N__42456));
    Span4Mux_v I__9329 (
            .O(N__42456),
            .I(N__42453));
    Odrv4 I__9328 (
            .O(N__42453),
            .I(\comm_spi.data_tx_7__N_773 ));
    CascadeMux I__9327 (
            .O(N__42450),
            .I(n17479_cascade_));
    InMux I__9326 (
            .O(N__42447),
            .I(N__42443));
    InMux I__9325 (
            .O(N__42446),
            .I(N__42440));
    LocalMux I__9324 (
            .O(N__42443),
            .I(N__42437));
    LocalMux I__9323 (
            .O(N__42440),
            .I(N__42432));
    Span4Mux_v I__9322 (
            .O(N__42437),
            .I(N__42432));
    Odrv4 I__9321 (
            .O(N__42432),
            .I(comm_buf_6_5));
    InMux I__9320 (
            .O(N__42429),
            .I(N__42426));
    LocalMux I__9319 (
            .O(N__42426),
            .I(N__42423));
    Span4Mux_h I__9318 (
            .O(N__42423),
            .I(N__42420));
    Odrv4 I__9317 (
            .O(N__42420),
            .I(comm_buf_2_5));
    InMux I__9316 (
            .O(N__42417),
            .I(N__42414));
    LocalMux I__9315 (
            .O(N__42414),
            .I(N__42411));
    Odrv4 I__9314 (
            .O(N__42411),
            .I(n17480));
    InMux I__9313 (
            .O(N__42408),
            .I(N__42405));
    LocalMux I__9312 (
            .O(N__42405),
            .I(comm_buf_5_5));
    InMux I__9311 (
            .O(N__42402),
            .I(N__42399));
    LocalMux I__9310 (
            .O(N__42399),
            .I(n21212));
    CascadeMux I__9309 (
            .O(N__42396),
            .I(n17482_cascade_));
    InMux I__9308 (
            .O(N__42393),
            .I(N__42390));
    LocalMux I__9307 (
            .O(N__42390),
            .I(n22189));
    InMux I__9306 (
            .O(N__42387),
            .I(N__42383));
    InMux I__9305 (
            .O(N__42386),
            .I(N__42380));
    LocalMux I__9304 (
            .O(N__42383),
            .I(N__42375));
    LocalMux I__9303 (
            .O(N__42380),
            .I(N__42375));
    Odrv12 I__9302 (
            .O(N__42375),
            .I(\comm_spi.n14639 ));
    SRMux I__9301 (
            .O(N__42372),
            .I(N__42369));
    LocalMux I__9300 (
            .O(N__42369),
            .I(N__42366));
    Span4Mux_h I__9299 (
            .O(N__42366),
            .I(N__42363));
    Odrv4 I__9298 (
            .O(N__42363),
            .I(\comm_spi.data_tx_7__N_777 ));
    SRMux I__9297 (
            .O(N__42360),
            .I(N__42357));
    LocalMux I__9296 (
            .O(N__42357),
            .I(N__42354));
    Span4Mux_v I__9295 (
            .O(N__42354),
            .I(N__42351));
    Odrv4 I__9294 (
            .O(N__42351),
            .I(\comm_spi.data_tx_7__N_780 ));
    InMux I__9293 (
            .O(N__42348),
            .I(N__42345));
    LocalMux I__9292 (
            .O(N__42345),
            .I(N__42342));
    Odrv4 I__9291 (
            .O(N__42342),
            .I(comm_buf_5_6));
    CascadeMux I__9290 (
            .O(N__42339),
            .I(n22183_cascade_));
    InMux I__9289 (
            .O(N__42336),
            .I(N__42333));
    LocalMux I__9288 (
            .O(N__42333),
            .I(N__42330));
    Span4Mux_h I__9287 (
            .O(N__42330),
            .I(N__42327));
    Odrv4 I__9286 (
            .O(N__42327),
            .I(comm_buf_5_0));
    InMux I__9285 (
            .O(N__42324),
            .I(N__42321));
    LocalMux I__9284 (
            .O(N__42321),
            .I(n4));
    InMux I__9283 (
            .O(N__42318),
            .I(N__42314));
    CascadeMux I__9282 (
            .O(N__42317),
            .I(N__42311));
    LocalMux I__9281 (
            .O(N__42314),
            .I(N__42308));
    InMux I__9280 (
            .O(N__42311),
            .I(N__42305));
    Span4Mux_v I__9279 (
            .O(N__42308),
            .I(N__42302));
    LocalMux I__9278 (
            .O(N__42305),
            .I(comm_buf_6_0));
    Odrv4 I__9277 (
            .O(N__42302),
            .I(comm_buf_6_0));
    CascadeMux I__9276 (
            .O(N__42297),
            .I(N__42294));
    InMux I__9275 (
            .O(N__42294),
            .I(N__42291));
    LocalMux I__9274 (
            .O(N__42291),
            .I(n21211));
    InMux I__9273 (
            .O(N__42288),
            .I(N__42279));
    CascadeMux I__9272 (
            .O(N__42287),
            .I(N__42276));
    InMux I__9271 (
            .O(N__42286),
            .I(N__42263));
    CascadeMux I__9270 (
            .O(N__42285),
            .I(N__42259));
    CascadeMux I__9269 (
            .O(N__42284),
            .I(N__42256));
    CascadeMux I__9268 (
            .O(N__42283),
            .I(N__42253));
    CascadeMux I__9267 (
            .O(N__42282),
            .I(N__42250));
    LocalMux I__9266 (
            .O(N__42279),
            .I(N__42245));
    InMux I__9265 (
            .O(N__42276),
            .I(N__42242));
    InMux I__9264 (
            .O(N__42275),
            .I(N__42225));
    InMux I__9263 (
            .O(N__42274),
            .I(N__42225));
    InMux I__9262 (
            .O(N__42273),
            .I(N__42225));
    InMux I__9261 (
            .O(N__42272),
            .I(N__42225));
    InMux I__9260 (
            .O(N__42271),
            .I(N__42225));
    InMux I__9259 (
            .O(N__42270),
            .I(N__42225));
    InMux I__9258 (
            .O(N__42269),
            .I(N__42225));
    InMux I__9257 (
            .O(N__42268),
            .I(N__42225));
    InMux I__9256 (
            .O(N__42267),
            .I(N__42222));
    InMux I__9255 (
            .O(N__42266),
            .I(N__42219));
    LocalMux I__9254 (
            .O(N__42263),
            .I(N__42216));
    InMux I__9253 (
            .O(N__42262),
            .I(N__42201));
    InMux I__9252 (
            .O(N__42259),
            .I(N__42201));
    InMux I__9251 (
            .O(N__42256),
            .I(N__42201));
    InMux I__9250 (
            .O(N__42253),
            .I(N__42201));
    InMux I__9249 (
            .O(N__42250),
            .I(N__42201));
    InMux I__9248 (
            .O(N__42249),
            .I(N__42201));
    InMux I__9247 (
            .O(N__42248),
            .I(N__42201));
    Span4Mux_h I__9246 (
            .O(N__42245),
            .I(N__42198));
    LocalMux I__9245 (
            .O(N__42242),
            .I(N__42191));
    LocalMux I__9244 (
            .O(N__42225),
            .I(N__42191));
    LocalMux I__9243 (
            .O(N__42222),
            .I(N__42185));
    LocalMux I__9242 (
            .O(N__42219),
            .I(N__42182));
    Span4Mux_v I__9241 (
            .O(N__42216),
            .I(N__42179));
    LocalMux I__9240 (
            .O(N__42201),
            .I(N__42174));
    Span4Mux_v I__9239 (
            .O(N__42198),
            .I(N__42174));
    InMux I__9238 (
            .O(N__42197),
            .I(N__42171));
    InMux I__9237 (
            .O(N__42196),
            .I(N__42168));
    Span4Mux_h I__9236 (
            .O(N__42191),
            .I(N__42165));
    InMux I__9235 (
            .O(N__42190),
            .I(N__42158));
    InMux I__9234 (
            .O(N__42189),
            .I(N__42158));
    InMux I__9233 (
            .O(N__42188),
            .I(N__42158));
    Span4Mux_h I__9232 (
            .O(N__42185),
            .I(N__42153));
    Span4Mux_v I__9231 (
            .O(N__42182),
            .I(N__42153));
    Span4Mux_v I__9230 (
            .O(N__42179),
            .I(N__42150));
    Span4Mux_v I__9229 (
            .O(N__42174),
            .I(N__42147));
    LocalMux I__9228 (
            .O(N__42171),
            .I(dds_state_2));
    LocalMux I__9227 (
            .O(N__42168),
            .I(dds_state_2));
    Odrv4 I__9226 (
            .O(N__42165),
            .I(dds_state_2));
    LocalMux I__9225 (
            .O(N__42158),
            .I(dds_state_2));
    Odrv4 I__9224 (
            .O(N__42153),
            .I(dds_state_2));
    Odrv4 I__9223 (
            .O(N__42150),
            .I(dds_state_2));
    Odrv4 I__9222 (
            .O(N__42147),
            .I(dds_state_2));
    CascadeMux I__9221 (
            .O(N__42132),
            .I(N__42128));
    InMux I__9220 (
            .O(N__42131),
            .I(N__42125));
    InMux I__9219 (
            .O(N__42128),
            .I(N__42121));
    LocalMux I__9218 (
            .O(N__42125),
            .I(N__42117));
    InMux I__9217 (
            .O(N__42124),
            .I(N__42114));
    LocalMux I__9216 (
            .O(N__42121),
            .I(N__42111));
    CascadeMux I__9215 (
            .O(N__42120),
            .I(N__42108));
    Span4Mux_v I__9214 (
            .O(N__42117),
            .I(N__42105));
    LocalMux I__9213 (
            .O(N__42114),
            .I(N__42100));
    Span4Mux_h I__9212 (
            .O(N__42111),
            .I(N__42100));
    InMux I__9211 (
            .O(N__42108),
            .I(N__42097));
    Odrv4 I__9210 (
            .O(N__42105),
            .I(trig_dds0));
    Odrv4 I__9209 (
            .O(N__42100),
            .I(trig_dds0));
    LocalMux I__9208 (
            .O(N__42097),
            .I(trig_dds0));
    CEMux I__9207 (
            .O(N__42090),
            .I(N__42086));
    CEMux I__9206 (
            .O(N__42089),
            .I(N__42083));
    LocalMux I__9205 (
            .O(N__42086),
            .I(N__42080));
    LocalMux I__9204 (
            .O(N__42083),
            .I(N__42077));
    Span4Mux_h I__9203 (
            .O(N__42080),
            .I(N__42074));
    Span4Mux_h I__9202 (
            .O(N__42077),
            .I(N__42071));
    Span4Mux_h I__9201 (
            .O(N__42074),
            .I(N__42068));
    Odrv4 I__9200 (
            .O(N__42071),
            .I(\SIG_DDS.n12722 ));
    Odrv4 I__9199 (
            .O(N__42068),
            .I(\SIG_DDS.n12722 ));
    InMux I__9198 (
            .O(N__42063),
            .I(N__42059));
    InMux I__9197 (
            .O(N__42062),
            .I(N__42055));
    LocalMux I__9196 (
            .O(N__42059),
            .I(N__42052));
    InMux I__9195 (
            .O(N__42058),
            .I(N__42049));
    LocalMux I__9194 (
            .O(N__42055),
            .I(data_index_8));
    Odrv4 I__9193 (
            .O(N__42052),
            .I(data_index_8));
    LocalMux I__9192 (
            .O(N__42049),
            .I(data_index_8));
    InMux I__9191 (
            .O(N__42042),
            .I(N__42039));
    LocalMux I__9190 (
            .O(N__42039),
            .I(N__42036));
    Span4Mux_h I__9189 (
            .O(N__42036),
            .I(N__42032));
    InMux I__9188 (
            .O(N__42035),
            .I(N__42029));
    Odrv4 I__9187 (
            .O(N__42032),
            .I(n8_adj_1561));
    LocalMux I__9186 (
            .O(N__42029),
            .I(n8_adj_1561));
    InMux I__9185 (
            .O(N__42024),
            .I(N__42020));
    InMux I__9184 (
            .O(N__42023),
            .I(N__42017));
    LocalMux I__9183 (
            .O(N__42020),
            .I(n8_adj_1563));
    LocalMux I__9182 (
            .O(N__42017),
            .I(n8_adj_1563));
    CascadeMux I__9181 (
            .O(N__42012),
            .I(N__42009));
    InMux I__9180 (
            .O(N__42009),
            .I(N__42006));
    LocalMux I__9179 (
            .O(N__42006),
            .I(N__42003));
    Span4Mux_h I__9178 (
            .O(N__42003),
            .I(N__41999));
    InMux I__9177 (
            .O(N__42002),
            .I(N__41996));
    Odrv4 I__9176 (
            .O(N__41999),
            .I(n7_adj_1562));
    LocalMux I__9175 (
            .O(N__41996),
            .I(n7_adj_1562));
    InMux I__9174 (
            .O(N__41991),
            .I(N__41987));
    InMux I__9173 (
            .O(N__41990),
            .I(N__41984));
    LocalMux I__9172 (
            .O(N__41987),
            .I(N__41979));
    LocalMux I__9171 (
            .O(N__41984),
            .I(N__41979));
    Span4Mux_h I__9170 (
            .O(N__41979),
            .I(N__41975));
    InMux I__9169 (
            .O(N__41978),
            .I(N__41972));
    Span4Mux_h I__9168 (
            .O(N__41975),
            .I(N__41969));
    LocalMux I__9167 (
            .O(N__41972),
            .I(data_index_7));
    Odrv4 I__9166 (
            .O(N__41969),
            .I(data_index_7));
    IoInMux I__9165 (
            .O(N__41964),
            .I(N__41961));
    LocalMux I__9164 (
            .O(N__41961),
            .I(N__41958));
    IoSpan4Mux I__9163 (
            .O(N__41958),
            .I(N__41955));
    Span4Mux_s3_v I__9162 (
            .O(N__41955),
            .I(N__41950));
    InMux I__9161 (
            .O(N__41954),
            .I(N__41947));
    InMux I__9160 (
            .O(N__41953),
            .I(N__41944));
    Span4Mux_v I__9159 (
            .O(N__41950),
            .I(N__41939));
    LocalMux I__9158 (
            .O(N__41947),
            .I(N__41939));
    LocalMux I__9157 (
            .O(N__41944),
            .I(SELIRNG1));
    Odrv4 I__9156 (
            .O(N__41939),
            .I(SELIRNG1));
    InMux I__9155 (
            .O(N__41934),
            .I(N__41931));
    LocalMux I__9154 (
            .O(N__41931),
            .I(N__41928));
    Span4Mux_h I__9153 (
            .O(N__41928),
            .I(N__41923));
    CascadeMux I__9152 (
            .O(N__41927),
            .I(N__41920));
    InMux I__9151 (
            .O(N__41926),
            .I(N__41917));
    Span4Mux_h I__9150 (
            .O(N__41923),
            .I(N__41914));
    InMux I__9149 (
            .O(N__41920),
            .I(N__41911));
    LocalMux I__9148 (
            .O(N__41917),
            .I(acadc_skipCount_11));
    Odrv4 I__9147 (
            .O(N__41914),
            .I(acadc_skipCount_11));
    LocalMux I__9146 (
            .O(N__41911),
            .I(acadc_skipCount_11));
    CascadeMux I__9145 (
            .O(N__41904),
            .I(N__41901));
    InMux I__9144 (
            .O(N__41901),
            .I(N__41898));
    LocalMux I__9143 (
            .O(N__41898),
            .I(N__41895));
    Odrv4 I__9142 (
            .O(N__41895),
            .I(n23_adj_1543));
    InMux I__9141 (
            .O(N__41892),
            .I(N__41888));
    InMux I__9140 (
            .O(N__41891),
            .I(N__41883));
    LocalMux I__9139 (
            .O(N__41888),
            .I(N__41880));
    InMux I__9138 (
            .O(N__41887),
            .I(N__41875));
    InMux I__9137 (
            .O(N__41886),
            .I(N__41875));
    LocalMux I__9136 (
            .O(N__41883),
            .I(N__41871));
    Span4Mux_h I__9135 (
            .O(N__41880),
            .I(N__41866));
    LocalMux I__9134 (
            .O(N__41875),
            .I(N__41866));
    InMux I__9133 (
            .O(N__41874),
            .I(N__41863));
    Span12Mux_h I__9132 (
            .O(N__41871),
            .I(N__41858));
    Span4Mux_h I__9131 (
            .O(N__41866),
            .I(N__41853));
    LocalMux I__9130 (
            .O(N__41863),
            .I(N__41853));
    InMux I__9129 (
            .O(N__41862),
            .I(N__41850));
    InMux I__9128 (
            .O(N__41861),
            .I(N__41847));
    Odrv12 I__9127 (
            .O(N__41858),
            .I(n11915));
    Odrv4 I__9126 (
            .O(N__41853),
            .I(n11915));
    LocalMux I__9125 (
            .O(N__41850),
            .I(n11915));
    LocalMux I__9124 (
            .O(N__41847),
            .I(n11915));
    InMux I__9123 (
            .O(N__41838),
            .I(N__41835));
    LocalMux I__9122 (
            .O(N__41835),
            .I(N__41832));
    Odrv12 I__9121 (
            .O(N__41832),
            .I(buf_data_iac_22));
    InMux I__9120 (
            .O(N__41829),
            .I(N__41826));
    LocalMux I__9119 (
            .O(N__41826),
            .I(N__41823));
    Span12Mux_h I__9118 (
            .O(N__41823),
            .I(N__41820));
    Odrv12 I__9117 (
            .O(N__41820),
            .I(n21273));
    InMux I__9116 (
            .O(N__41817),
            .I(N__41814));
    LocalMux I__9115 (
            .O(N__41814),
            .I(N__41811));
    Span4Mux_h I__9114 (
            .O(N__41811),
            .I(N__41808));
    Odrv4 I__9113 (
            .O(N__41808),
            .I(buf_data_iac_20));
    InMux I__9112 (
            .O(N__41805),
            .I(N__41802));
    LocalMux I__9111 (
            .O(N__41802),
            .I(N__41799));
    Span4Mux_v I__9110 (
            .O(N__41799),
            .I(N__41796));
    Span4Mux_v I__9109 (
            .O(N__41796),
            .I(N__41793));
    Odrv4 I__9108 (
            .O(N__41793),
            .I(n21569));
    InMux I__9107 (
            .O(N__41790),
            .I(N__41786));
    InMux I__9106 (
            .O(N__41789),
            .I(N__41783));
    LocalMux I__9105 (
            .O(N__41786),
            .I(\comm_spi.n14592 ));
    LocalMux I__9104 (
            .O(N__41783),
            .I(\comm_spi.n14592 ));
    InMux I__9103 (
            .O(N__41778),
            .I(N__41774));
    InMux I__9102 (
            .O(N__41777),
            .I(N__41771));
    LocalMux I__9101 (
            .O(N__41774),
            .I(N__41768));
    LocalMux I__9100 (
            .O(N__41771),
            .I(N__41765));
    Span4Mux_h I__9099 (
            .O(N__41768),
            .I(N__41757));
    Span4Mux_v I__9098 (
            .O(N__41765),
            .I(N__41757));
    InMux I__9097 (
            .O(N__41764),
            .I(N__41754));
    InMux I__9096 (
            .O(N__41763),
            .I(N__41749));
    InMux I__9095 (
            .O(N__41762),
            .I(N__41749));
    Odrv4 I__9094 (
            .O(N__41757),
            .I(n20907));
    LocalMux I__9093 (
            .O(N__41754),
            .I(n20907));
    LocalMux I__9092 (
            .O(N__41749),
            .I(n20907));
    InMux I__9091 (
            .O(N__41742),
            .I(N__41736));
    InMux I__9090 (
            .O(N__41741),
            .I(N__41731));
    InMux I__9089 (
            .O(N__41740),
            .I(N__41731));
    CascadeMux I__9088 (
            .O(N__41739),
            .I(N__41726));
    LocalMux I__9087 (
            .O(N__41736),
            .I(N__41718));
    LocalMux I__9086 (
            .O(N__41731),
            .I(N__41718));
    InMux I__9085 (
            .O(N__41730),
            .I(N__41713));
    InMux I__9084 (
            .O(N__41729),
            .I(N__41713));
    InMux I__9083 (
            .O(N__41726),
            .I(N__41708));
    InMux I__9082 (
            .O(N__41725),
            .I(N__41708));
    CascadeMux I__9081 (
            .O(N__41724),
            .I(N__41705));
    InMux I__9080 (
            .O(N__41723),
            .I(N__41695));
    Span4Mux_v I__9079 (
            .O(N__41718),
            .I(N__41688));
    LocalMux I__9078 (
            .O(N__41713),
            .I(N__41688));
    LocalMux I__9077 (
            .O(N__41708),
            .I(N__41688));
    InMux I__9076 (
            .O(N__41705),
            .I(N__41679));
    InMux I__9075 (
            .O(N__41704),
            .I(N__41679));
    InMux I__9074 (
            .O(N__41703),
            .I(N__41679));
    InMux I__9073 (
            .O(N__41702),
            .I(N__41679));
    InMux I__9072 (
            .O(N__41701),
            .I(N__41672));
    InMux I__9071 (
            .O(N__41700),
            .I(N__41672));
    InMux I__9070 (
            .O(N__41699),
            .I(N__41672));
    InMux I__9069 (
            .O(N__41698),
            .I(N__41669));
    LocalMux I__9068 (
            .O(N__41695),
            .I(N__41666));
    Span4Mux_h I__9067 (
            .O(N__41688),
            .I(N__41663));
    LocalMux I__9066 (
            .O(N__41679),
            .I(N__41660));
    LocalMux I__9065 (
            .O(N__41672),
            .I(N__41655));
    LocalMux I__9064 (
            .O(N__41669),
            .I(N__41655));
    Span4Mux_v I__9063 (
            .O(N__41666),
            .I(N__41652));
    Span4Mux_h I__9062 (
            .O(N__41663),
            .I(N__41649));
    Span4Mux_h I__9061 (
            .O(N__41660),
            .I(N__41646));
    Span4Mux_h I__9060 (
            .O(N__41655),
            .I(N__41643));
    Odrv4 I__9059 (
            .O(N__41652),
            .I(n12429));
    Odrv4 I__9058 (
            .O(N__41649),
            .I(n12429));
    Odrv4 I__9057 (
            .O(N__41646),
            .I(n12429));
    Odrv4 I__9056 (
            .O(N__41643),
            .I(n12429));
    CascadeMux I__9055 (
            .O(N__41634),
            .I(n9306_cascade_));
    InMux I__9054 (
            .O(N__41631),
            .I(N__41627));
    InMux I__9053 (
            .O(N__41630),
            .I(N__41624));
    LocalMux I__9052 (
            .O(N__41627),
            .I(N__41621));
    LocalMux I__9051 (
            .O(N__41624),
            .I(N__41618));
    Span4Mux_v I__9050 (
            .O(N__41621),
            .I(N__41612));
    Span4Mux_h I__9049 (
            .O(N__41618),
            .I(N__41612));
    InMux I__9048 (
            .O(N__41617),
            .I(N__41609));
    Span4Mux_h I__9047 (
            .O(N__41612),
            .I(N__41606));
    LocalMux I__9046 (
            .O(N__41609),
            .I(buf_dds0_13));
    Odrv4 I__9045 (
            .O(N__41606),
            .I(buf_dds0_13));
    InMux I__9044 (
            .O(N__41601),
            .I(N__41598));
    LocalMux I__9043 (
            .O(N__41598),
            .I(N__41594));
    InMux I__9042 (
            .O(N__41597),
            .I(N__41591));
    Span4Mux_h I__9041 (
            .O(N__41594),
            .I(N__41588));
    LocalMux I__9040 (
            .O(N__41591),
            .I(acadc_skipcnt_7));
    Odrv4 I__9039 (
            .O(N__41588),
            .I(acadc_skipcnt_7));
    InMux I__9038 (
            .O(N__41583),
            .I(N__41580));
    LocalMux I__9037 (
            .O(N__41580),
            .I(N__41576));
    InMux I__9036 (
            .O(N__41579),
            .I(N__41573));
    Span4Mux_v I__9035 (
            .O(N__41576),
            .I(N__41570));
    LocalMux I__9034 (
            .O(N__41573),
            .I(acadc_skipcnt_2));
    Odrv4 I__9033 (
            .O(N__41570),
            .I(acadc_skipcnt_2));
    InMux I__9032 (
            .O(N__41565),
            .I(N__41562));
    LocalMux I__9031 (
            .O(N__41562),
            .I(N__41559));
    Span4Mux_h I__9030 (
            .O(N__41559),
            .I(N__41556));
    Odrv4 I__9029 (
            .O(N__41556),
            .I(n22));
    InMux I__9028 (
            .O(N__41553),
            .I(N__41549));
    InMux I__9027 (
            .O(N__41552),
            .I(N__41546));
    LocalMux I__9026 (
            .O(N__41549),
            .I(n9));
    LocalMux I__9025 (
            .O(N__41546),
            .I(n9));
    CascadeMux I__9024 (
            .O(N__41541),
            .I(N__41537));
    CascadeMux I__9023 (
            .O(N__41540),
            .I(N__41534));
    InMux I__9022 (
            .O(N__41537),
            .I(N__41529));
    InMux I__9021 (
            .O(N__41534),
            .I(N__41526));
    InMux I__9020 (
            .O(N__41533),
            .I(N__41523));
    CascadeMux I__9019 (
            .O(N__41532),
            .I(N__41520));
    LocalMux I__9018 (
            .O(N__41529),
            .I(N__41517));
    LocalMux I__9017 (
            .O(N__41526),
            .I(N__41514));
    LocalMux I__9016 (
            .O(N__41523),
            .I(N__41511));
    InMux I__9015 (
            .O(N__41520),
            .I(N__41508));
    Span4Mux_v I__9014 (
            .O(N__41517),
            .I(N__41503));
    Span4Mux_v I__9013 (
            .O(N__41514),
            .I(N__41503));
    Odrv12 I__9012 (
            .O(N__41511),
            .I(n20912));
    LocalMux I__9011 (
            .O(N__41508),
            .I(n20912));
    Odrv4 I__9010 (
            .O(N__41503),
            .I(n20912));
    CascadeMux I__9009 (
            .O(N__41496),
            .I(N__41488));
    CascadeMux I__9008 (
            .O(N__41495),
            .I(N__41485));
    InMux I__9007 (
            .O(N__41494),
            .I(N__41481));
    CascadeMux I__9006 (
            .O(N__41493),
            .I(N__41478));
    CascadeMux I__9005 (
            .O(N__41492),
            .I(N__41475));
    CascadeMux I__9004 (
            .O(N__41491),
            .I(N__41472));
    InMux I__9003 (
            .O(N__41488),
            .I(N__41469));
    InMux I__9002 (
            .O(N__41485),
            .I(N__41466));
    InMux I__9001 (
            .O(N__41484),
            .I(N__41462));
    LocalMux I__9000 (
            .O(N__41481),
            .I(N__41459));
    InMux I__8999 (
            .O(N__41478),
            .I(N__41456));
    InMux I__8998 (
            .O(N__41475),
            .I(N__41453));
    InMux I__8997 (
            .O(N__41472),
            .I(N__41450));
    LocalMux I__8996 (
            .O(N__41469),
            .I(N__41447));
    LocalMux I__8995 (
            .O(N__41466),
            .I(N__41444));
    InMux I__8994 (
            .O(N__41465),
            .I(N__41441));
    LocalMux I__8993 (
            .O(N__41462),
            .I(N__41438));
    Span4Mux_v I__8992 (
            .O(N__41459),
            .I(N__41433));
    LocalMux I__8991 (
            .O(N__41456),
            .I(N__41433));
    LocalMux I__8990 (
            .O(N__41453),
            .I(N__41428));
    LocalMux I__8989 (
            .O(N__41450),
            .I(N__41428));
    Span12Mux_h I__8988 (
            .O(N__41447),
            .I(N__41425));
    Span4Mux_v I__8987 (
            .O(N__41444),
            .I(N__41422));
    LocalMux I__8986 (
            .O(N__41441),
            .I(N__41417));
    Sp12to4 I__8985 (
            .O(N__41438),
            .I(N__41417));
    Span4Mux_h I__8984 (
            .O(N__41433),
            .I(N__41412));
    Span4Mux_v I__8983 (
            .O(N__41428),
            .I(N__41412));
    Odrv12 I__8982 (
            .O(N__41425),
            .I(comm_buf_0_4));
    Odrv4 I__8981 (
            .O(N__41422),
            .I(comm_buf_0_4));
    Odrv12 I__8980 (
            .O(N__41417),
            .I(comm_buf_0_4));
    Odrv4 I__8979 (
            .O(N__41412),
            .I(comm_buf_0_4));
    CascadeMux I__8978 (
            .O(N__41403),
            .I(n12381_cascade_));
    IoInMux I__8977 (
            .O(N__41400),
            .I(N__41397));
    LocalMux I__8976 (
            .O(N__41397),
            .I(N__41394));
    Span4Mux_s3_h I__8975 (
            .O(N__41394),
            .I(N__41391));
    Span4Mux_h I__8974 (
            .O(N__41391),
            .I(N__41388));
    Sp12to4 I__8973 (
            .O(N__41388),
            .I(N__41384));
    InMux I__8972 (
            .O(N__41387),
            .I(N__41381));
    Span12Mux_s11_v I__8971 (
            .O(N__41384),
            .I(N__41378));
    LocalMux I__8970 (
            .O(N__41381),
            .I(N__41374));
    Span12Mux_h I__8969 (
            .O(N__41378),
            .I(N__41371));
    InMux I__8968 (
            .O(N__41377),
            .I(N__41368));
    Span4Mux_v I__8967 (
            .O(N__41374),
            .I(N__41365));
    Odrv12 I__8966 (
            .O(N__41371),
            .I(VAC_OSR0));
    LocalMux I__8965 (
            .O(N__41368),
            .I(VAC_OSR0));
    Odrv4 I__8964 (
            .O(N__41365),
            .I(VAC_OSR0));
    InMux I__8963 (
            .O(N__41358),
            .I(N__41354));
    InMux I__8962 (
            .O(N__41357),
            .I(N__41351));
    LocalMux I__8961 (
            .O(N__41354),
            .I(N__41345));
    LocalMux I__8960 (
            .O(N__41351),
            .I(N__41345));
    InMux I__8959 (
            .O(N__41350),
            .I(N__41342));
    Odrv4 I__8958 (
            .O(N__41345),
            .I(acadc_skipCount_6));
    LocalMux I__8957 (
            .O(N__41342),
            .I(acadc_skipCount_6));
    InMux I__8956 (
            .O(N__41337),
            .I(N__41331));
    CascadeMux I__8955 (
            .O(N__41336),
            .I(N__41328));
    InMux I__8954 (
            .O(N__41335),
            .I(N__41324));
    InMux I__8953 (
            .O(N__41334),
            .I(N__41320));
    LocalMux I__8952 (
            .O(N__41331),
            .I(N__41317));
    InMux I__8951 (
            .O(N__41328),
            .I(N__41312));
    InMux I__8950 (
            .O(N__41327),
            .I(N__41312));
    LocalMux I__8949 (
            .O(N__41324),
            .I(N__41308));
    InMux I__8948 (
            .O(N__41323),
            .I(N__41305));
    LocalMux I__8947 (
            .O(N__41320),
            .I(N__41302));
    Span4Mux_v I__8946 (
            .O(N__41317),
            .I(N__41296));
    LocalMux I__8945 (
            .O(N__41312),
            .I(N__41296));
    InMux I__8944 (
            .O(N__41311),
            .I(N__41293));
    Span4Mux_h I__8943 (
            .O(N__41308),
            .I(N__41288));
    LocalMux I__8942 (
            .O(N__41305),
            .I(N__41288));
    Span4Mux_v I__8941 (
            .O(N__41302),
            .I(N__41285));
    InMux I__8940 (
            .O(N__41301),
            .I(N__41281));
    Span4Mux_v I__8939 (
            .O(N__41296),
            .I(N__41276));
    LocalMux I__8938 (
            .O(N__41293),
            .I(N__41276));
    Span4Mux_v I__8937 (
            .O(N__41288),
            .I(N__41273));
    Sp12to4 I__8936 (
            .O(N__41285),
            .I(N__41270));
    InMux I__8935 (
            .O(N__41284),
            .I(N__41267));
    LocalMux I__8934 (
            .O(N__41281),
            .I(N__41264));
    Span4Mux_h I__8933 (
            .O(N__41276),
            .I(N__41261));
    Span4Mux_h I__8932 (
            .O(N__41273),
            .I(N__41258));
    Span12Mux_h I__8931 (
            .O(N__41270),
            .I(N__41255));
    LocalMux I__8930 (
            .O(N__41267),
            .I(dds_state_0));
    Odrv12 I__8929 (
            .O(N__41264),
            .I(dds_state_0));
    Odrv4 I__8928 (
            .O(N__41261),
            .I(dds_state_0));
    Odrv4 I__8927 (
            .O(N__41258),
            .I(dds_state_0));
    Odrv12 I__8926 (
            .O(N__41255),
            .I(dds_state_0));
    CascadeMux I__8925 (
            .O(N__41244),
            .I(N__41241));
    InMux I__8924 (
            .O(N__41241),
            .I(N__41237));
    InMux I__8923 (
            .O(N__41240),
            .I(N__41234));
    LocalMux I__8922 (
            .O(N__41237),
            .I(data_idxvec_10));
    LocalMux I__8921 (
            .O(N__41234),
            .I(data_idxvec_10));
    InMux I__8920 (
            .O(N__41229),
            .I(N__41226));
    LocalMux I__8919 (
            .O(N__41226),
            .I(N__41222));
    InMux I__8918 (
            .O(N__41225),
            .I(N__41218));
    Span4Mux_h I__8917 (
            .O(N__41222),
            .I(N__41215));
    InMux I__8916 (
            .O(N__41221),
            .I(N__41212));
    LocalMux I__8915 (
            .O(N__41218),
            .I(data_cntvec_10));
    Odrv4 I__8914 (
            .O(N__41215),
            .I(data_cntvec_10));
    LocalMux I__8913 (
            .O(N__41212),
            .I(data_cntvec_10));
    InMux I__8912 (
            .O(N__41205),
            .I(N__41202));
    LocalMux I__8911 (
            .O(N__41202),
            .I(N__41199));
    Odrv4 I__8910 (
            .O(N__41199),
            .I(n21150));
    CascadeMux I__8909 (
            .O(N__41196),
            .I(N__41192));
    CascadeMux I__8908 (
            .O(N__41195),
            .I(N__41189));
    InMux I__8907 (
            .O(N__41192),
            .I(N__41186));
    InMux I__8906 (
            .O(N__41189),
            .I(N__41183));
    LocalMux I__8905 (
            .O(N__41186),
            .I(N__41180));
    LocalMux I__8904 (
            .O(N__41183),
            .I(data_idxvec_9));
    Odrv4 I__8903 (
            .O(N__41180),
            .I(data_idxvec_9));
    InMux I__8902 (
            .O(N__41175),
            .I(N__41172));
    LocalMux I__8901 (
            .O(N__41172),
            .I(N__41168));
    InMux I__8900 (
            .O(N__41171),
            .I(N__41164));
    Span4Mux_v I__8899 (
            .O(N__41168),
            .I(N__41161));
    InMux I__8898 (
            .O(N__41167),
            .I(N__41158));
    LocalMux I__8897 (
            .O(N__41164),
            .I(data_cntvec_9));
    Odrv4 I__8896 (
            .O(N__41161),
            .I(data_cntvec_9));
    LocalMux I__8895 (
            .O(N__41158),
            .I(data_cntvec_9));
    InMux I__8894 (
            .O(N__41151),
            .I(N__41148));
    LocalMux I__8893 (
            .O(N__41148),
            .I(N__41145));
    Odrv12 I__8892 (
            .O(N__41145),
            .I(n21060));
    InMux I__8891 (
            .O(N__41142),
            .I(N__41139));
    LocalMux I__8890 (
            .O(N__41139),
            .I(N__41136));
    Span4Mux_h I__8889 (
            .O(N__41136),
            .I(N__41132));
    InMux I__8888 (
            .O(N__41135),
            .I(N__41129));
    Odrv4 I__8887 (
            .O(N__41132),
            .I(n8_adj_1569));
    LocalMux I__8886 (
            .O(N__41129),
            .I(n8_adj_1569));
    InMux I__8885 (
            .O(N__41124),
            .I(N__41120));
    CascadeMux I__8884 (
            .O(N__41123),
            .I(N__41117));
    LocalMux I__8883 (
            .O(N__41120),
            .I(N__41114));
    InMux I__8882 (
            .O(N__41117),
            .I(N__41111));
    Span4Mux_v I__8881 (
            .O(N__41114),
            .I(N__41108));
    LocalMux I__8880 (
            .O(N__41111),
            .I(N__41105));
    Odrv4 I__8879 (
            .O(N__41108),
            .I(n7_adj_1568));
    Odrv4 I__8878 (
            .O(N__41105),
            .I(n7_adj_1568));
    InMux I__8877 (
            .O(N__41100),
            .I(N__41095));
    InMux I__8876 (
            .O(N__41099),
            .I(N__41092));
    InMux I__8875 (
            .O(N__41098),
            .I(N__41089));
    LocalMux I__8874 (
            .O(N__41095),
            .I(N__41084));
    LocalMux I__8873 (
            .O(N__41092),
            .I(N__41084));
    LocalMux I__8872 (
            .O(N__41089),
            .I(N__41081));
    Span4Mux_v I__8871 (
            .O(N__41084),
            .I(N__41078));
    Span4Mux_h I__8870 (
            .O(N__41081),
            .I(N__41075));
    Odrv4 I__8869 (
            .O(N__41078),
            .I(data_index_3));
    Odrv4 I__8868 (
            .O(N__41075),
            .I(data_index_3));
    InMux I__8867 (
            .O(N__41070),
            .I(N__41066));
    CascadeMux I__8866 (
            .O(N__41069),
            .I(N__41063));
    LocalMux I__8865 (
            .O(N__41066),
            .I(N__41060));
    InMux I__8864 (
            .O(N__41063),
            .I(N__41057));
    Span4Mux_h I__8863 (
            .O(N__41060),
            .I(N__41054));
    LocalMux I__8862 (
            .O(N__41057),
            .I(data_idxvec_8));
    Odrv4 I__8861 (
            .O(N__41054),
            .I(data_idxvec_8));
    InMux I__8860 (
            .O(N__41049),
            .I(N__41046));
    LocalMux I__8859 (
            .O(N__41046),
            .I(N__41042));
    InMux I__8858 (
            .O(N__41045),
            .I(N__41038));
    Span4Mux_h I__8857 (
            .O(N__41042),
            .I(N__41035));
    InMux I__8856 (
            .O(N__41041),
            .I(N__41032));
    LocalMux I__8855 (
            .O(N__41038),
            .I(data_cntvec_8));
    Odrv4 I__8854 (
            .O(N__41035),
            .I(data_cntvec_8));
    LocalMux I__8853 (
            .O(N__41032),
            .I(data_cntvec_8));
    InMux I__8852 (
            .O(N__41025),
            .I(N__41022));
    LocalMux I__8851 (
            .O(N__41022),
            .I(N__41017));
    InMux I__8850 (
            .O(N__41021),
            .I(N__41012));
    InMux I__8849 (
            .O(N__41020),
            .I(N__41012));
    Odrv4 I__8848 (
            .O(N__41017),
            .I(req_data_cnt_11));
    LocalMux I__8847 (
            .O(N__41012),
            .I(req_data_cnt_11));
    CascadeMux I__8846 (
            .O(N__41007),
            .I(n8_adj_1571_cascade_));
    InMux I__8845 (
            .O(N__41004),
            .I(N__41000));
    InMux I__8844 (
            .O(N__41003),
            .I(N__40997));
    LocalMux I__8843 (
            .O(N__41000),
            .I(N__40991));
    LocalMux I__8842 (
            .O(N__40997),
            .I(N__40991));
    InMux I__8841 (
            .O(N__40996),
            .I(N__40988));
    Span4Mux_h I__8840 (
            .O(N__40991),
            .I(N__40985));
    LocalMux I__8839 (
            .O(N__40988),
            .I(data_index_2));
    Odrv4 I__8838 (
            .O(N__40985),
            .I(data_index_2));
    InMux I__8837 (
            .O(N__40980),
            .I(N__40977));
    LocalMux I__8836 (
            .O(N__40977),
            .I(N__40973));
    InMux I__8835 (
            .O(N__40976),
            .I(N__40970));
    Span4Mux_v I__8834 (
            .O(N__40973),
            .I(N__40964));
    LocalMux I__8833 (
            .O(N__40970),
            .I(N__40964));
    InMux I__8832 (
            .O(N__40969),
            .I(N__40961));
    Span4Mux_h I__8831 (
            .O(N__40964),
            .I(N__40958));
    LocalMux I__8830 (
            .O(N__40961),
            .I(buf_dds0_10));
    Odrv4 I__8829 (
            .O(N__40958),
            .I(buf_dds0_10));
    CascadeMux I__8828 (
            .O(N__40953),
            .I(N__40950));
    InMux I__8827 (
            .O(N__40950),
            .I(N__40946));
    InMux I__8826 (
            .O(N__40949),
            .I(N__40943));
    LocalMux I__8825 (
            .O(N__40946),
            .I(data_idxvec_11));
    LocalMux I__8824 (
            .O(N__40943),
            .I(data_idxvec_11));
    InMux I__8823 (
            .O(N__40938),
            .I(N__40933));
    InMux I__8822 (
            .O(N__40937),
            .I(N__40930));
    InMux I__8821 (
            .O(N__40936),
            .I(N__40927));
    LocalMux I__8820 (
            .O(N__40933),
            .I(N__40924));
    LocalMux I__8819 (
            .O(N__40930),
            .I(data_cntvec_11));
    LocalMux I__8818 (
            .O(N__40927),
            .I(data_cntvec_11));
    Odrv4 I__8817 (
            .O(N__40924),
            .I(data_cntvec_11));
    InMux I__8816 (
            .O(N__40917),
            .I(N__40914));
    LocalMux I__8815 (
            .O(N__40914),
            .I(N__40911));
    Span4Mux_v I__8814 (
            .O(N__40911),
            .I(N__40908));
    Span4Mux_h I__8813 (
            .O(N__40908),
            .I(N__40905));
    Odrv4 I__8812 (
            .O(N__40905),
            .I(buf_data_iac_19));
    CascadeMux I__8811 (
            .O(N__40902),
            .I(n26_adj_1544_cascade_));
    InMux I__8810 (
            .O(N__40899),
            .I(N__40895));
    InMux I__8809 (
            .O(N__40898),
            .I(N__40892));
    LocalMux I__8808 (
            .O(N__40895),
            .I(N__40886));
    LocalMux I__8807 (
            .O(N__40892),
            .I(N__40881));
    SRMux I__8806 (
            .O(N__40891),
            .I(N__40878));
    InMux I__8805 (
            .O(N__40890),
            .I(N__40874));
    SRMux I__8804 (
            .O(N__40889),
            .I(N__40871));
    Span4Mux_h I__8803 (
            .O(N__40886),
            .I(N__40868));
    InMux I__8802 (
            .O(N__40885),
            .I(N__40865));
    InMux I__8801 (
            .O(N__40884),
            .I(N__40859));
    Span4Mux_h I__8800 (
            .O(N__40881),
            .I(N__40854));
    LocalMux I__8799 (
            .O(N__40878),
            .I(N__40854));
    InMux I__8798 (
            .O(N__40877),
            .I(N__40851));
    LocalMux I__8797 (
            .O(N__40874),
            .I(N__40848));
    LocalMux I__8796 (
            .O(N__40871),
            .I(N__40841));
    Span4Mux_h I__8795 (
            .O(N__40868),
            .I(N__40841));
    LocalMux I__8794 (
            .O(N__40865),
            .I(N__40841));
    InMux I__8793 (
            .O(N__40864),
            .I(N__40834));
    InMux I__8792 (
            .O(N__40863),
            .I(N__40834));
    InMux I__8791 (
            .O(N__40862),
            .I(N__40834));
    LocalMux I__8790 (
            .O(N__40859),
            .I(acadc_rst));
    Odrv4 I__8789 (
            .O(N__40854),
            .I(acadc_rst));
    LocalMux I__8788 (
            .O(N__40851),
            .I(acadc_rst));
    Odrv12 I__8787 (
            .O(N__40848),
            .I(acadc_rst));
    Odrv4 I__8786 (
            .O(N__40841),
            .I(acadc_rst));
    LocalMux I__8785 (
            .O(N__40834),
            .I(acadc_rst));
    InMux I__8784 (
            .O(N__40821),
            .I(N__40817));
    CascadeMux I__8783 (
            .O(N__40820),
            .I(N__40814));
    LocalMux I__8782 (
            .O(N__40817),
            .I(N__40810));
    InMux I__8781 (
            .O(N__40814),
            .I(N__40807));
    InMux I__8780 (
            .O(N__40813),
            .I(N__40804));
    Span4Mux_h I__8779 (
            .O(N__40810),
            .I(N__40801));
    LocalMux I__8778 (
            .O(N__40807),
            .I(N__40798));
    LocalMux I__8777 (
            .O(N__40804),
            .I(req_data_cnt_10));
    Odrv4 I__8776 (
            .O(N__40801),
            .I(req_data_cnt_10));
    Odrv4 I__8775 (
            .O(N__40798),
            .I(req_data_cnt_10));
    InMux I__8774 (
            .O(N__40791),
            .I(N__40788));
    LocalMux I__8773 (
            .O(N__40788),
            .I(n21088));
    InMux I__8772 (
            .O(N__40785),
            .I(N__40782));
    LocalMux I__8771 (
            .O(N__40782),
            .I(N__40778));
    InMux I__8770 (
            .O(N__40781),
            .I(N__40774));
    Span4Mux_v I__8769 (
            .O(N__40778),
            .I(N__40771));
    InMux I__8768 (
            .O(N__40777),
            .I(N__40768));
    LocalMux I__8767 (
            .O(N__40774),
            .I(req_data_cnt_6));
    Odrv4 I__8766 (
            .O(N__40771),
            .I(req_data_cnt_6));
    LocalMux I__8765 (
            .O(N__40768),
            .I(req_data_cnt_6));
    InMux I__8764 (
            .O(N__40761),
            .I(N__40758));
    LocalMux I__8763 (
            .O(N__40758),
            .I(N__40755));
    Span4Mux_v I__8762 (
            .O(N__40755),
            .I(N__40751));
    InMux I__8761 (
            .O(N__40754),
            .I(N__40747));
    Span4Mux_h I__8760 (
            .O(N__40751),
            .I(N__40744));
    InMux I__8759 (
            .O(N__40750),
            .I(N__40741));
    LocalMux I__8758 (
            .O(N__40747),
            .I(buf_dds1_6));
    Odrv4 I__8757 (
            .O(N__40744),
            .I(buf_dds1_6));
    LocalMux I__8756 (
            .O(N__40741),
            .I(buf_dds1_6));
    InMux I__8755 (
            .O(N__40734),
            .I(N__40731));
    LocalMux I__8754 (
            .O(N__40731),
            .I(N__40726));
    InMux I__8753 (
            .O(N__40730),
            .I(N__40721));
    InMux I__8752 (
            .O(N__40729),
            .I(N__40721));
    Odrv12 I__8751 (
            .O(N__40726),
            .I(buf_dds0_6));
    LocalMux I__8750 (
            .O(N__40721),
            .I(buf_dds0_6));
    InMux I__8749 (
            .O(N__40716),
            .I(N__40712));
    InMux I__8748 (
            .O(N__40715),
            .I(N__40709));
    LocalMux I__8747 (
            .O(N__40712),
            .I(N__40706));
    LocalMux I__8746 (
            .O(N__40709),
            .I(N__40703));
    Span4Mux_v I__8745 (
            .O(N__40706),
            .I(N__40700));
    Span4Mux_v I__8744 (
            .O(N__40703),
            .I(N__40697));
    Sp12to4 I__8743 (
            .O(N__40700),
            .I(N__40691));
    Sp12to4 I__8742 (
            .O(N__40697),
            .I(N__40691));
    InMux I__8741 (
            .O(N__40696),
            .I(N__40688));
    Span12Mux_h I__8740 (
            .O(N__40691),
            .I(N__40685));
    LocalMux I__8739 (
            .O(N__40688),
            .I(buf_adcdata_iac_18));
    Odrv12 I__8738 (
            .O(N__40685),
            .I(buf_adcdata_iac_18));
    InMux I__8737 (
            .O(N__40680),
            .I(N__40677));
    LocalMux I__8736 (
            .O(N__40677),
            .I(n21073));
    CascadeMux I__8735 (
            .O(N__40674),
            .I(N__40671));
    InMux I__8734 (
            .O(N__40671),
            .I(N__40663));
    InMux I__8733 (
            .O(N__40670),
            .I(N__40660));
    InMux I__8732 (
            .O(N__40669),
            .I(N__40657));
    InMux I__8731 (
            .O(N__40668),
            .I(N__40652));
    InMux I__8730 (
            .O(N__40667),
            .I(N__40649));
    InMux I__8729 (
            .O(N__40666),
            .I(N__40646));
    LocalMux I__8728 (
            .O(N__40663),
            .I(N__40643));
    LocalMux I__8727 (
            .O(N__40660),
            .I(N__40638));
    LocalMux I__8726 (
            .O(N__40657),
            .I(N__40638));
    CascadeMux I__8725 (
            .O(N__40656),
            .I(N__40632));
    InMux I__8724 (
            .O(N__40655),
            .I(N__40628));
    LocalMux I__8723 (
            .O(N__40652),
            .I(N__40625));
    LocalMux I__8722 (
            .O(N__40649),
            .I(N__40622));
    LocalMux I__8721 (
            .O(N__40646),
            .I(N__40619));
    Span4Mux_v I__8720 (
            .O(N__40643),
            .I(N__40614));
    Span4Mux_v I__8719 (
            .O(N__40638),
            .I(N__40614));
    InMux I__8718 (
            .O(N__40637),
            .I(N__40611));
    InMux I__8717 (
            .O(N__40636),
            .I(N__40608));
    InMux I__8716 (
            .O(N__40635),
            .I(N__40605));
    InMux I__8715 (
            .O(N__40632),
            .I(N__40600));
    InMux I__8714 (
            .O(N__40631),
            .I(N__40600));
    LocalMux I__8713 (
            .O(N__40628),
            .I(N__40597));
    Span4Mux_h I__8712 (
            .O(N__40625),
            .I(N__40594));
    Span4Mux_h I__8711 (
            .O(N__40622),
            .I(N__40591));
    Span4Mux_v I__8710 (
            .O(N__40619),
            .I(N__40586));
    Span4Mux_h I__8709 (
            .O(N__40614),
            .I(N__40586));
    LocalMux I__8708 (
            .O(N__40611),
            .I(n16891));
    LocalMux I__8707 (
            .O(N__40608),
            .I(n16891));
    LocalMux I__8706 (
            .O(N__40605),
            .I(n16891));
    LocalMux I__8705 (
            .O(N__40600),
            .I(n16891));
    Odrv12 I__8704 (
            .O(N__40597),
            .I(n16891));
    Odrv4 I__8703 (
            .O(N__40594),
            .I(n16891));
    Odrv4 I__8702 (
            .O(N__40591),
            .I(n16891));
    Odrv4 I__8701 (
            .O(N__40586),
            .I(n16891));
    InMux I__8700 (
            .O(N__40569),
            .I(N__40564));
    InMux I__8699 (
            .O(N__40568),
            .I(N__40561));
    InMux I__8698 (
            .O(N__40567),
            .I(N__40558));
    LocalMux I__8697 (
            .O(N__40564),
            .I(N__40551));
    LocalMux I__8696 (
            .O(N__40561),
            .I(N__40551));
    LocalMux I__8695 (
            .O(N__40558),
            .I(N__40551));
    Span4Mux_h I__8694 (
            .O(N__40551),
            .I(N__40548));
    Odrv4 I__8693 (
            .O(N__40548),
            .I(data_index_5));
    InMux I__8692 (
            .O(N__40545),
            .I(N__40542));
    LocalMux I__8691 (
            .O(N__40542),
            .I(n22306));
    InMux I__8690 (
            .O(N__40539),
            .I(N__40536));
    LocalMux I__8689 (
            .O(N__40536),
            .I(N__40533));
    Odrv12 I__8688 (
            .O(N__40533),
            .I(n22420));
    InMux I__8687 (
            .O(N__40530),
            .I(N__40527));
    LocalMux I__8686 (
            .O(N__40527),
            .I(n22246));
    CascadeMux I__8685 (
            .O(N__40524),
            .I(n21092_cascade_));
    CascadeMux I__8684 (
            .O(N__40521),
            .I(n30_adj_1542_cascade_));
    InMux I__8683 (
            .O(N__40518),
            .I(N__40515));
    LocalMux I__8682 (
            .O(N__40515),
            .I(N__40512));
    Odrv12 I__8681 (
            .O(N__40512),
            .I(n21087));
    CascadeMux I__8680 (
            .O(N__40509),
            .I(n22357_cascade_));
    CascadeMux I__8679 (
            .O(N__40506),
            .I(n22360_cascade_));
    CascadeMux I__8678 (
            .O(N__40503),
            .I(n21137_cascade_));
    CascadeMux I__8677 (
            .O(N__40500),
            .I(N__40497));
    InMux I__8676 (
            .O(N__40497),
            .I(N__40494));
    LocalMux I__8675 (
            .O(N__40494),
            .I(N__40491));
    Odrv12 I__8674 (
            .O(N__40491),
            .I(n21072));
    InMux I__8673 (
            .O(N__40488),
            .I(N__40485));
    LocalMux I__8672 (
            .O(N__40485),
            .I(N__40482));
    Odrv12 I__8671 (
            .O(N__40482),
            .I(n22327));
    InMux I__8670 (
            .O(N__40479),
            .I(N__40476));
    LocalMux I__8669 (
            .O(N__40476),
            .I(n22330));
    CascadeMux I__8668 (
            .O(N__40473),
            .I(n22288_cascade_));
    InMux I__8667 (
            .O(N__40470),
            .I(N__40467));
    LocalMux I__8666 (
            .O(N__40467),
            .I(n22276));
    CascadeMux I__8665 (
            .O(N__40464),
            .I(n30_adj_1539_cascade_));
    InMux I__8664 (
            .O(N__40461),
            .I(N__40458));
    LocalMux I__8663 (
            .O(N__40458),
            .I(N__40455));
    Span4Mux_v I__8662 (
            .O(N__40455),
            .I(N__40452));
    Span4Mux_v I__8661 (
            .O(N__40452),
            .I(N__40448));
    CascadeMux I__8660 (
            .O(N__40451),
            .I(N__40445));
    Span4Mux_h I__8659 (
            .O(N__40448),
            .I(N__40442));
    InMux I__8658 (
            .O(N__40445),
            .I(N__40439));
    Odrv4 I__8657 (
            .O(N__40442),
            .I(buf_adcdata_vdc_22));
    LocalMux I__8656 (
            .O(N__40439),
            .I(buf_adcdata_vdc_22));
    InMux I__8655 (
            .O(N__40434),
            .I(N__40430));
    InMux I__8654 (
            .O(N__40433),
            .I(N__40426));
    LocalMux I__8653 (
            .O(N__40430),
            .I(N__40423));
    CascadeMux I__8652 (
            .O(N__40429),
            .I(N__40420));
    LocalMux I__8651 (
            .O(N__40426),
            .I(N__40415));
    Span12Mux_v I__8650 (
            .O(N__40423),
            .I(N__40415));
    InMux I__8649 (
            .O(N__40420),
            .I(N__40412));
    Span12Mux_h I__8648 (
            .O(N__40415),
            .I(N__40409));
    LocalMux I__8647 (
            .O(N__40412),
            .I(buf_adcdata_vac_22));
    Odrv12 I__8646 (
            .O(N__40409),
            .I(buf_adcdata_vac_22));
    InMux I__8645 (
            .O(N__40404),
            .I(N__40401));
    LocalMux I__8644 (
            .O(N__40401),
            .I(N__40398));
    Odrv12 I__8643 (
            .O(N__40398),
            .I(n20_adj_1537));
    CascadeMux I__8642 (
            .O(N__40395),
            .I(n19_adj_1536_cascade_));
    InMux I__8641 (
            .O(N__40392),
            .I(N__40389));
    LocalMux I__8640 (
            .O(N__40389),
            .I(n22285));
    InMux I__8639 (
            .O(N__40386),
            .I(N__40382));
    CascadeMux I__8638 (
            .O(N__40385),
            .I(N__40379));
    LocalMux I__8637 (
            .O(N__40382),
            .I(N__40376));
    InMux I__8636 (
            .O(N__40379),
            .I(N__40373));
    Sp12to4 I__8635 (
            .O(N__40376),
            .I(N__40370));
    LocalMux I__8634 (
            .O(N__40373),
            .I(N__40366));
    Span12Mux_v I__8633 (
            .O(N__40370),
            .I(N__40363));
    InMux I__8632 (
            .O(N__40369),
            .I(N__40360));
    Span12Mux_h I__8631 (
            .O(N__40366),
            .I(N__40357));
    Span12Mux_h I__8630 (
            .O(N__40363),
            .I(N__40354));
    LocalMux I__8629 (
            .O(N__40360),
            .I(buf_adcdata_iac_20));
    Odrv12 I__8628 (
            .O(N__40357),
            .I(buf_adcdata_iac_20));
    Odrv12 I__8627 (
            .O(N__40354),
            .I(buf_adcdata_iac_20));
    InMux I__8626 (
            .O(N__40347),
            .I(N__40343));
    InMux I__8625 (
            .O(N__40346),
            .I(N__40340));
    LocalMux I__8624 (
            .O(N__40343),
            .I(N__40336));
    LocalMux I__8623 (
            .O(N__40340),
            .I(N__40333));
    InMux I__8622 (
            .O(N__40339),
            .I(N__40330));
    Span12Mux_h I__8621 (
            .O(N__40336),
            .I(N__40327));
    Odrv4 I__8620 (
            .O(N__40333),
            .I(buf_dds0_12));
    LocalMux I__8619 (
            .O(N__40330),
            .I(buf_dds0_12));
    Odrv12 I__8618 (
            .O(N__40327),
            .I(buf_dds0_12));
    CascadeMux I__8617 (
            .O(N__40320),
            .I(n22303_cascade_));
    InMux I__8616 (
            .O(N__40317),
            .I(N__40313));
    InMux I__8615 (
            .O(N__40316),
            .I(N__40310));
    LocalMux I__8614 (
            .O(N__40313),
            .I(N__40306));
    LocalMux I__8613 (
            .O(N__40310),
            .I(N__40303));
    InMux I__8612 (
            .O(N__40309),
            .I(N__40300));
    Span4Mux_h I__8611 (
            .O(N__40306),
            .I(N__40297));
    Span4Mux_v I__8610 (
            .O(N__40303),
            .I(N__40294));
    LocalMux I__8609 (
            .O(N__40300),
            .I(buf_dds1_12));
    Odrv4 I__8608 (
            .O(N__40297),
            .I(buf_dds1_12));
    Odrv4 I__8607 (
            .O(N__40294),
            .I(buf_dds1_12));
    InMux I__8606 (
            .O(N__40287),
            .I(N__40284));
    LocalMux I__8605 (
            .O(N__40284),
            .I(N__40281));
    Span12Mux_v I__8604 (
            .O(N__40281),
            .I(N__40278));
    Odrv12 I__8603 (
            .O(N__40278),
            .I(n21309));
    CascadeMux I__8602 (
            .O(N__40275),
            .I(N__40272));
    InMux I__8601 (
            .O(N__40272),
            .I(N__40269));
    LocalMux I__8600 (
            .O(N__40269),
            .I(N__40266));
    Span4Mux_h I__8599 (
            .O(N__40266),
            .I(N__40263));
    Odrv4 I__8598 (
            .O(N__40263),
            .I(n23_adj_1541));
    CascadeMux I__8597 (
            .O(N__40260),
            .I(N__40257));
    InMux I__8596 (
            .O(N__40257),
            .I(N__40254));
    LocalMux I__8595 (
            .O(N__40254),
            .I(n21568));
    InMux I__8594 (
            .O(N__40251),
            .I(N__40248));
    LocalMux I__8593 (
            .O(N__40248),
            .I(n22243));
    CascadeMux I__8592 (
            .O(N__40245),
            .I(n22237_cascade_));
    InMux I__8591 (
            .O(N__40242),
            .I(N__40238));
    InMux I__8590 (
            .O(N__40241),
            .I(N__40234));
    LocalMux I__8589 (
            .O(N__40238),
            .I(N__40231));
    InMux I__8588 (
            .O(N__40237),
            .I(N__40228));
    LocalMux I__8587 (
            .O(N__40234),
            .I(N__40225));
    Span4Mux_h I__8586 (
            .O(N__40231),
            .I(N__40222));
    LocalMux I__8585 (
            .O(N__40228),
            .I(buf_dds1_9));
    Odrv4 I__8584 (
            .O(N__40225),
            .I(buf_dds1_9));
    Odrv4 I__8583 (
            .O(N__40222),
            .I(buf_dds1_9));
    InMux I__8582 (
            .O(N__40215),
            .I(N__40212));
    LocalMux I__8581 (
            .O(N__40212),
            .I(N__40209));
    Odrv12 I__8580 (
            .O(N__40209),
            .I(buf_data_iac_17));
    InMux I__8579 (
            .O(N__40206),
            .I(N__40203));
    LocalMux I__8578 (
            .O(N__40203),
            .I(N__40200));
    Span4Mux_h I__8577 (
            .O(N__40200),
            .I(N__40197));
    Span4Mux_v I__8576 (
            .O(N__40197),
            .I(N__40194));
    Odrv4 I__8575 (
            .O(N__40194),
            .I(n22378));
    CascadeMux I__8574 (
            .O(N__40191),
            .I(n21062_cascade_));
    InMux I__8573 (
            .O(N__40188),
            .I(N__40185));
    LocalMux I__8572 (
            .O(N__40185),
            .I(n22240));
    InMux I__8571 (
            .O(N__40182),
            .I(N__40179));
    LocalMux I__8570 (
            .O(N__40179),
            .I(N__40176));
    Span4Mux_h I__8569 (
            .O(N__40176),
            .I(N__40173));
    Span4Mux_h I__8568 (
            .O(N__40173),
            .I(N__40170));
    Odrv4 I__8567 (
            .O(N__40170),
            .I(n22444));
    CascadeMux I__8566 (
            .O(N__40167),
            .I(n22447_cascade_));
    CascadeMux I__8565 (
            .O(N__40164),
            .I(n22450_cascade_));
    CascadeMux I__8564 (
            .O(N__40161),
            .I(N__40157));
    CascadeMux I__8563 (
            .O(N__40160),
            .I(N__40152));
    InMux I__8562 (
            .O(N__40157),
            .I(N__40149));
    CascadeMux I__8561 (
            .O(N__40156),
            .I(N__40146));
    CascadeMux I__8560 (
            .O(N__40155),
            .I(N__40142));
    InMux I__8559 (
            .O(N__40152),
            .I(N__40139));
    LocalMux I__8558 (
            .O(N__40149),
            .I(N__40136));
    InMux I__8557 (
            .O(N__40146),
            .I(N__40132));
    InMux I__8556 (
            .O(N__40145),
            .I(N__40129));
    InMux I__8555 (
            .O(N__40142),
            .I(N__40126));
    LocalMux I__8554 (
            .O(N__40139),
            .I(N__40123));
    Span4Mux_v I__8553 (
            .O(N__40136),
            .I(N__40116));
    InMux I__8552 (
            .O(N__40135),
            .I(N__40113));
    LocalMux I__8551 (
            .O(N__40132),
            .I(N__40110));
    LocalMux I__8550 (
            .O(N__40129),
            .I(N__40107));
    LocalMux I__8549 (
            .O(N__40126),
            .I(N__40104));
    Span4Mux_v I__8548 (
            .O(N__40123),
            .I(N__40101));
    InMux I__8547 (
            .O(N__40122),
            .I(N__40098));
    InMux I__8546 (
            .O(N__40121),
            .I(N__40095));
    InMux I__8545 (
            .O(N__40120),
            .I(N__40092));
    InMux I__8544 (
            .O(N__40119),
            .I(N__40089));
    Span4Mux_h I__8543 (
            .O(N__40116),
            .I(N__40084));
    LocalMux I__8542 (
            .O(N__40113),
            .I(N__40084));
    Span4Mux_v I__8541 (
            .O(N__40110),
            .I(N__40081));
    Span4Mux_h I__8540 (
            .O(N__40107),
            .I(N__40078));
    Span4Mux_h I__8539 (
            .O(N__40104),
            .I(N__40071));
    Span4Mux_h I__8538 (
            .O(N__40101),
            .I(N__40071));
    LocalMux I__8537 (
            .O(N__40098),
            .I(N__40071));
    LocalMux I__8536 (
            .O(N__40095),
            .I(N__40068));
    LocalMux I__8535 (
            .O(N__40092),
            .I(N__40065));
    LocalMux I__8534 (
            .O(N__40089),
            .I(N__40054));
    Span4Mux_h I__8533 (
            .O(N__40084),
            .I(N__40054));
    Span4Mux_h I__8532 (
            .O(N__40081),
            .I(N__40054));
    Span4Mux_v I__8531 (
            .O(N__40078),
            .I(N__40054));
    Span4Mux_v I__8530 (
            .O(N__40071),
            .I(N__40054));
    Span12Mux_h I__8529 (
            .O(N__40068),
            .I(N__40051));
    Span12Mux_v I__8528 (
            .O(N__40065),
            .I(N__40048));
    Span4Mux_v I__8527 (
            .O(N__40054),
            .I(N__40045));
    Odrv12 I__8526 (
            .O(N__40051),
            .I(comm_buf_0_1));
    Odrv12 I__8525 (
            .O(N__40048),
            .I(comm_buf_0_1));
    Odrv4 I__8524 (
            .O(N__40045),
            .I(comm_buf_0_1));
    CascadeMux I__8523 (
            .O(N__40038),
            .I(N__40035));
    InMux I__8522 (
            .O(N__40035),
            .I(N__40032));
    LocalMux I__8521 (
            .O(N__40032),
            .I(n30));
    CascadeMux I__8520 (
            .O(N__40029),
            .I(N__40026));
    InMux I__8519 (
            .O(N__40026),
            .I(N__40023));
    LocalMux I__8518 (
            .O(N__40023),
            .I(n21272));
    InMux I__8517 (
            .O(N__40020),
            .I(N__40017));
    LocalMux I__8516 (
            .O(N__40017),
            .I(N__40014));
    Span4Mux_h I__8515 (
            .O(N__40014),
            .I(N__40011));
    Odrv4 I__8514 (
            .O(N__40011),
            .I(n23_adj_1538));
    CascadeMux I__8513 (
            .O(N__40008),
            .I(n22273_cascade_));
    InMux I__8512 (
            .O(N__40005),
            .I(N__40002));
    LocalMux I__8511 (
            .O(N__40002),
            .I(N__39999));
    Span4Mux_h I__8510 (
            .O(N__39999),
            .I(N__39996));
    Odrv4 I__8509 (
            .O(N__39996),
            .I(n21286));
    InMux I__8508 (
            .O(N__39993),
            .I(N__39990));
    LocalMux I__8507 (
            .O(N__39990),
            .I(N__39987));
    Span4Mux_h I__8506 (
            .O(N__39987),
            .I(N__39984));
    Span4Mux_h I__8505 (
            .O(N__39984),
            .I(N__39981));
    Odrv4 I__8504 (
            .O(N__39981),
            .I(n17_adj_1535));
    CascadeMux I__8503 (
            .O(N__39978),
            .I(N__39975));
    InMux I__8502 (
            .O(N__39975),
            .I(N__39972));
    LocalMux I__8501 (
            .O(N__39972),
            .I(N__39969));
    Span4Mux_v I__8500 (
            .O(N__39969),
            .I(N__39966));
    Sp12to4 I__8499 (
            .O(N__39966),
            .I(N__39963));
    Odrv12 I__8498 (
            .O(N__39963),
            .I(n16_adj_1534));
    CascadeMux I__8497 (
            .O(N__39960),
            .I(N__39957));
    InMux I__8496 (
            .O(N__39957),
            .I(N__39954));
    LocalMux I__8495 (
            .O(N__39954),
            .I(N__39951));
    Span12Mux_v I__8494 (
            .O(N__39951),
            .I(N__39948));
    Span12Mux_h I__8493 (
            .O(N__39948),
            .I(N__39945));
    Odrv12 I__8492 (
            .O(N__39945),
            .I(buf_data_vac_7));
    InMux I__8491 (
            .O(N__39942),
            .I(N__39939));
    LocalMux I__8490 (
            .O(N__39939),
            .I(N__39936));
    Span4Mux_v I__8489 (
            .O(N__39936),
            .I(N__39933));
    Odrv4 I__8488 (
            .O(N__39933),
            .I(comm_buf_5_7));
    InMux I__8487 (
            .O(N__39930),
            .I(N__39927));
    LocalMux I__8486 (
            .O(N__39927),
            .I(N__39924));
    Span12Mux_v I__8485 (
            .O(N__39924),
            .I(N__39921));
    Span12Mux_h I__8484 (
            .O(N__39921),
            .I(N__39918));
    Odrv12 I__8483 (
            .O(N__39918),
            .I(buf_data_vac_6));
    InMux I__8482 (
            .O(N__39915),
            .I(N__39912));
    LocalMux I__8481 (
            .O(N__39912),
            .I(N__39909));
    Span12Mux_v I__8480 (
            .O(N__39909),
            .I(N__39906));
    Span12Mux_h I__8479 (
            .O(N__39906),
            .I(N__39903));
    Odrv12 I__8478 (
            .O(N__39903),
            .I(buf_data_vac_5));
    InMux I__8477 (
            .O(N__39900),
            .I(N__39897));
    LocalMux I__8476 (
            .O(N__39897),
            .I(N__39894));
    Span12Mux_v I__8475 (
            .O(N__39894),
            .I(N__39891));
    Span12Mux_h I__8474 (
            .O(N__39891),
            .I(N__39888));
    Odrv12 I__8473 (
            .O(N__39888),
            .I(buf_data_vac_4));
    InMux I__8472 (
            .O(N__39885),
            .I(N__39882));
    LocalMux I__8471 (
            .O(N__39882),
            .I(N__39879));
    Odrv4 I__8470 (
            .O(N__39879),
            .I(comm_buf_5_4));
    InMux I__8469 (
            .O(N__39876),
            .I(N__39873));
    LocalMux I__8468 (
            .O(N__39873),
            .I(N__39870));
    Span4Mux_v I__8467 (
            .O(N__39870),
            .I(N__39867));
    Span4Mux_h I__8466 (
            .O(N__39867),
            .I(N__39864));
    Odrv4 I__8465 (
            .O(N__39864),
            .I(buf_data_vac_3));
    InMux I__8464 (
            .O(N__39861),
            .I(N__39858));
    LocalMux I__8463 (
            .O(N__39858),
            .I(N__39855));
    Span4Mux_h I__8462 (
            .O(N__39855),
            .I(N__39852));
    Odrv4 I__8461 (
            .O(N__39852),
            .I(comm_buf_5_3));
    InMux I__8460 (
            .O(N__39849),
            .I(N__39846));
    LocalMux I__8459 (
            .O(N__39846),
            .I(N__39843));
    Span4Mux_v I__8458 (
            .O(N__39843),
            .I(N__39840));
    Span4Mux_h I__8457 (
            .O(N__39840),
            .I(N__39837));
    Odrv4 I__8456 (
            .O(N__39837),
            .I(buf_data_vac_2));
    InMux I__8455 (
            .O(N__39834),
            .I(N__39831));
    LocalMux I__8454 (
            .O(N__39831),
            .I(comm_buf_5_2));
    InMux I__8453 (
            .O(N__39828),
            .I(N__39825));
    LocalMux I__8452 (
            .O(N__39825),
            .I(N__39822));
    Span4Mux_h I__8451 (
            .O(N__39822),
            .I(N__39819));
    Span4Mux_h I__8450 (
            .O(N__39819),
            .I(N__39816));
    Odrv4 I__8449 (
            .O(N__39816),
            .I(buf_data_vac_1));
    InMux I__8448 (
            .O(N__39813),
            .I(N__39810));
    LocalMux I__8447 (
            .O(N__39810),
            .I(comm_buf_5_1));
    IoInMux I__8446 (
            .O(N__39807),
            .I(N__39804));
    LocalMux I__8445 (
            .O(N__39804),
            .I(N__39801));
    Span4Mux_s3_v I__8444 (
            .O(N__39801),
            .I(N__39797));
    InMux I__8443 (
            .O(N__39800),
            .I(N__39794));
    Span4Mux_h I__8442 (
            .O(N__39797),
            .I(N__39791));
    LocalMux I__8441 (
            .O(N__39794),
            .I(N__39788));
    Span4Mux_v I__8440 (
            .O(N__39791),
            .I(N__39784));
    Span4Mux_h I__8439 (
            .O(N__39788),
            .I(N__39781));
    InMux I__8438 (
            .O(N__39787),
            .I(N__39778));
    Span4Mux_v I__8437 (
            .O(N__39784),
            .I(N__39773));
    Span4Mux_h I__8436 (
            .O(N__39781),
            .I(N__39773));
    LocalMux I__8435 (
            .O(N__39778),
            .I(IAC_OSR1));
    Odrv4 I__8434 (
            .O(N__39773),
            .I(IAC_OSR1));
    InMux I__8433 (
            .O(N__39768),
            .I(N__39765));
    LocalMux I__8432 (
            .O(N__39765),
            .I(N__39762));
    Span4Mux_h I__8431 (
            .O(N__39762),
            .I(N__39758));
    InMux I__8430 (
            .O(N__39761),
            .I(N__39755));
    Span4Mux_h I__8429 (
            .O(N__39758),
            .I(N__39749));
    LocalMux I__8428 (
            .O(N__39755),
            .I(N__39749));
    InMux I__8427 (
            .O(N__39754),
            .I(N__39746));
    Span4Mux_h I__8426 (
            .O(N__39749),
            .I(N__39743));
    LocalMux I__8425 (
            .O(N__39746),
            .I(buf_adcdata_iac_17));
    Odrv4 I__8424 (
            .O(N__39743),
            .I(buf_adcdata_iac_17));
    InMux I__8423 (
            .O(N__39738),
            .I(N__39735));
    LocalMux I__8422 (
            .O(N__39735),
            .I(N__39732));
    Span4Mux_v I__8421 (
            .O(N__39732),
            .I(N__39729));
    Span4Mux_h I__8420 (
            .O(N__39729),
            .I(N__39724));
    InMux I__8419 (
            .O(N__39728),
            .I(N__39721));
    InMux I__8418 (
            .O(N__39727),
            .I(N__39718));
    Span4Mux_v I__8417 (
            .O(N__39724),
            .I(N__39715));
    LocalMux I__8416 (
            .O(N__39721),
            .I(buf_dds0_9));
    LocalMux I__8415 (
            .O(N__39718),
            .I(buf_dds0_9));
    Odrv4 I__8414 (
            .O(N__39715),
            .I(buf_dds0_9));
    InMux I__8413 (
            .O(N__39708),
            .I(N__39705));
    LocalMux I__8412 (
            .O(N__39705),
            .I(N__39702));
    Span4Mux_h I__8411 (
            .O(N__39702),
            .I(N__39699));
    Odrv4 I__8410 (
            .O(N__39699),
            .I(comm_buf_2_2));
    CascadeMux I__8409 (
            .O(N__39696),
            .I(n22393_cascade_));
    InMux I__8408 (
            .O(N__39693),
            .I(N__39690));
    LocalMux I__8407 (
            .O(N__39690),
            .I(N__39687));
    Span4Mux_v I__8406 (
            .O(N__39687),
            .I(N__39683));
    InMux I__8405 (
            .O(N__39686),
            .I(N__39680));
    Span4Mux_h I__8404 (
            .O(N__39683),
            .I(N__39677));
    LocalMux I__8403 (
            .O(N__39680),
            .I(comm_buf_6_2));
    Odrv4 I__8402 (
            .O(N__39677),
            .I(comm_buf_6_2));
    CascadeMux I__8401 (
            .O(N__39672),
            .I(n4_adj_1595_cascade_));
    InMux I__8400 (
            .O(N__39669),
            .I(N__39666));
    LocalMux I__8399 (
            .O(N__39666),
            .I(n22396));
    CascadeMux I__8398 (
            .O(N__39663),
            .I(n21196_cascade_));
    InMux I__8397 (
            .O(N__39660),
            .I(N__39651));
    InMux I__8396 (
            .O(N__39659),
            .I(N__39651));
    InMux I__8395 (
            .O(N__39658),
            .I(N__39651));
    LocalMux I__8394 (
            .O(N__39651),
            .I(N__39648));
    Span4Mux_v I__8393 (
            .O(N__39648),
            .I(N__39645));
    Odrv4 I__8392 (
            .O(N__39645),
            .I(comm_tx_buf_2));
    InMux I__8391 (
            .O(N__39642),
            .I(N__39639));
    LocalMux I__8390 (
            .O(N__39639),
            .I(N__39635));
    InMux I__8389 (
            .O(N__39638),
            .I(N__39632));
    Span4Mux_h I__8388 (
            .O(N__39635),
            .I(N__39629));
    LocalMux I__8387 (
            .O(N__39632),
            .I(comm_buf_6_1));
    Odrv4 I__8386 (
            .O(N__39629),
            .I(comm_buf_6_1));
    CascadeMux I__8385 (
            .O(N__39624),
            .I(n4_adj_1596_cascade_));
    InMux I__8384 (
            .O(N__39621),
            .I(N__39618));
    LocalMux I__8383 (
            .O(N__39618),
            .I(N__39615));
    Span4Mux_h I__8382 (
            .O(N__39615),
            .I(N__39612));
    Odrv4 I__8381 (
            .O(N__39612),
            .I(n22252));
    CascadeMux I__8380 (
            .O(N__39609),
            .I(n21052_cascade_));
    InMux I__8379 (
            .O(N__39606),
            .I(N__39597));
    InMux I__8378 (
            .O(N__39605),
            .I(N__39597));
    InMux I__8377 (
            .O(N__39604),
            .I(N__39597));
    LocalMux I__8376 (
            .O(N__39597),
            .I(N__39594));
    Span4Mux_v I__8375 (
            .O(N__39594),
            .I(N__39591));
    Odrv4 I__8374 (
            .O(N__39591),
            .I(comm_tx_buf_1));
    InMux I__8373 (
            .O(N__39588),
            .I(N__39585));
    LocalMux I__8372 (
            .O(N__39585),
            .I(N__39582));
    Span4Mux_h I__8371 (
            .O(N__39582),
            .I(N__39579));
    Span4Mux_h I__8370 (
            .O(N__39579),
            .I(N__39576));
    Odrv4 I__8369 (
            .O(N__39576),
            .I(buf_data_vac_0));
    SRMux I__8368 (
            .O(N__39573),
            .I(N__39570));
    LocalMux I__8367 (
            .O(N__39570),
            .I(N__39566));
    SRMux I__8366 (
            .O(N__39569),
            .I(N__39563));
    Span4Mux_v I__8365 (
            .O(N__39566),
            .I(N__39560));
    LocalMux I__8364 (
            .O(N__39563),
            .I(N__39557));
    Span4Mux_h I__8363 (
            .O(N__39560),
            .I(N__39554));
    Span4Mux_v I__8362 (
            .O(N__39557),
            .I(N__39551));
    Odrv4 I__8361 (
            .O(N__39554),
            .I(n20378));
    Odrv4 I__8360 (
            .O(N__39551),
            .I(n20378));
    InMux I__8359 (
            .O(N__39546),
            .I(N__39543));
    LocalMux I__8358 (
            .O(N__39543),
            .I(N__39540));
    Odrv12 I__8357 (
            .O(N__39540),
            .I(comm_buf_2_4));
    InMux I__8356 (
            .O(N__39537),
            .I(N__39534));
    LocalMux I__8355 (
            .O(N__39534),
            .I(N__39531));
    Span4Mux_h I__8354 (
            .O(N__39531),
            .I(N__39527));
    InMux I__8353 (
            .O(N__39530),
            .I(N__39524));
    Span4Mux_h I__8352 (
            .O(N__39527),
            .I(N__39521));
    LocalMux I__8351 (
            .O(N__39524),
            .I(comm_buf_6_4));
    Odrv4 I__8350 (
            .O(N__39521),
            .I(comm_buf_6_4));
    CascadeMux I__8349 (
            .O(N__39516),
            .I(n21538_cascade_));
    InMux I__8348 (
            .O(N__39513),
            .I(N__39510));
    LocalMux I__8347 (
            .O(N__39510),
            .I(n1_adj_1591));
    CascadeMux I__8346 (
            .O(N__39507),
            .I(n22369_cascade_));
    InMux I__8345 (
            .O(N__39504),
            .I(N__39501));
    LocalMux I__8344 (
            .O(N__39501),
            .I(n2_adj_1592));
    InMux I__8343 (
            .O(N__39498),
            .I(N__39495));
    LocalMux I__8342 (
            .O(N__39495),
            .I(n4_adj_1593));
    SRMux I__8341 (
            .O(N__39492),
            .I(N__39489));
    LocalMux I__8340 (
            .O(N__39489),
            .I(N__39486));
    Odrv4 I__8339 (
            .O(N__39486),
            .I(\comm_spi.data_tx_7__N_783 ));
    InMux I__8338 (
            .O(N__39483),
            .I(N__39480));
    LocalMux I__8337 (
            .O(N__39480),
            .I(N__39477));
    Span4Mux_v I__8336 (
            .O(N__39477),
            .I(N__39472));
    InMux I__8335 (
            .O(N__39476),
            .I(N__39467));
    InMux I__8334 (
            .O(N__39475),
            .I(N__39467));
    Odrv4 I__8333 (
            .O(N__39472),
            .I(comm_tx_buf_4));
    LocalMux I__8332 (
            .O(N__39467),
            .I(comm_tx_buf_4));
    SRMux I__8331 (
            .O(N__39462),
            .I(N__39459));
    LocalMux I__8330 (
            .O(N__39459),
            .I(N__39456));
    Span4Mux_v I__8329 (
            .O(N__39456),
            .I(N__39453));
    Sp12to4 I__8328 (
            .O(N__39453),
            .I(N__39450));
    Odrv12 I__8327 (
            .O(N__39450),
            .I(\comm_spi.data_tx_7__N_769 ));
    CEMux I__8326 (
            .O(N__39447),
            .I(N__39444));
    LocalMux I__8325 (
            .O(N__39444),
            .I(N__39441));
    Odrv12 I__8324 (
            .O(N__39441),
            .I(n11741));
    InMux I__8323 (
            .O(N__39438),
            .I(N__39435));
    LocalMux I__8322 (
            .O(N__39435),
            .I(n20992));
    CascadeMux I__8321 (
            .O(N__39432),
            .I(n9255_cascade_));
    SRMux I__8320 (
            .O(N__39429),
            .I(N__39426));
    LocalMux I__8319 (
            .O(N__39426),
            .I(N__39423));
    Span4Mux_h I__8318 (
            .O(N__39423),
            .I(N__39420));
    Odrv4 I__8317 (
            .O(N__39420),
            .I(n14737));
    SRMux I__8316 (
            .O(N__39417),
            .I(N__39414));
    LocalMux I__8315 (
            .O(N__39414),
            .I(N__39410));
    SRMux I__8314 (
            .O(N__39413),
            .I(N__39407));
    Span4Mux_v I__8313 (
            .O(N__39410),
            .I(N__39404));
    LocalMux I__8312 (
            .O(N__39407),
            .I(N__39401));
    Span4Mux_h I__8311 (
            .O(N__39404),
            .I(N__39398));
    Span12Mux_v I__8310 (
            .O(N__39401),
            .I(N__39395));
    Odrv4 I__8309 (
            .O(N__39398),
            .I(flagcntwd));
    Odrv12 I__8308 (
            .O(N__39395),
            .I(flagcntwd));
    CEMux I__8307 (
            .O(N__39390),
            .I(N__39387));
    LocalMux I__8306 (
            .O(N__39387),
            .I(N__39384));
    Span4Mux_h I__8305 (
            .O(N__39384),
            .I(N__39381));
    Odrv4 I__8304 (
            .O(N__39381),
            .I(n11390));
    CascadeMux I__8303 (
            .O(N__39378),
            .I(n12336_cascade_));
    SRMux I__8302 (
            .O(N__39375),
            .I(N__39372));
    LocalMux I__8301 (
            .O(N__39372),
            .I(N__39369));
    Span4Mux_h I__8300 (
            .O(N__39369),
            .I(N__39366));
    Odrv4 I__8299 (
            .O(N__39366),
            .I(\comm_spi.data_tx_7__N_772 ));
    SRMux I__8298 (
            .O(N__39363),
            .I(N__39360));
    LocalMux I__8297 (
            .O(N__39360),
            .I(N__39357));
    Span4Mux_h I__8296 (
            .O(N__39357),
            .I(N__39354));
    Odrv4 I__8295 (
            .O(N__39354),
            .I(\comm_spi.data_tx_7__N_792 ));
    InMux I__8294 (
            .O(N__39351),
            .I(N__39348));
    LocalMux I__8293 (
            .O(N__39348),
            .I(N__39345));
    Sp12to4 I__8292 (
            .O(N__39345),
            .I(N__39341));
    InMux I__8291 (
            .O(N__39344),
            .I(N__39338));
    Span12Mux_v I__8290 (
            .O(N__39341),
            .I(N__39334));
    LocalMux I__8289 (
            .O(N__39338),
            .I(N__39331));
    InMux I__8288 (
            .O(N__39337),
            .I(N__39328));
    Odrv12 I__8287 (
            .O(N__39334),
            .I(\comm_spi.n22881 ));
    Odrv4 I__8286 (
            .O(N__39331),
            .I(\comm_spi.n22881 ));
    LocalMux I__8285 (
            .O(N__39328),
            .I(\comm_spi.n22881 ));
    SRMux I__8284 (
            .O(N__39321),
            .I(N__39318));
    LocalMux I__8283 (
            .O(N__39318),
            .I(N__39315));
    Span12Mux_s9_v I__8282 (
            .O(N__39315),
            .I(N__39312));
    Odrv12 I__8281 (
            .O(N__39312),
            .I(\comm_spi.data_tx_7__N_789 ));
    SRMux I__8280 (
            .O(N__39309),
            .I(N__39306));
    LocalMux I__8279 (
            .O(N__39306),
            .I(N__39303));
    Span4Mux_v I__8278 (
            .O(N__39303),
            .I(N__39300));
    Span4Mux_v I__8277 (
            .O(N__39300),
            .I(N__39297));
    Span4Mux_v I__8276 (
            .O(N__39297),
            .I(N__39294));
    Odrv4 I__8275 (
            .O(N__39294),
            .I(\comm_spi.data_tx_7__N_771 ));
    InMux I__8274 (
            .O(N__39291),
            .I(N__39288));
    LocalMux I__8273 (
            .O(N__39288),
            .I(N__39284));
    InMux I__8272 (
            .O(N__39287),
            .I(N__39281));
    Span4Mux_v I__8271 (
            .O(N__39284),
            .I(N__39276));
    LocalMux I__8270 (
            .O(N__39281),
            .I(N__39276));
    Span4Mux_v I__8269 (
            .O(N__39276),
            .I(N__39272));
    InMux I__8268 (
            .O(N__39275),
            .I(N__39269));
    Odrv4 I__8267 (
            .O(N__39272),
            .I(\comm_spi.n22878 ));
    LocalMux I__8266 (
            .O(N__39269),
            .I(\comm_spi.n22878 ));
    CascadeMux I__8265 (
            .O(N__39264),
            .I(N__39261));
    InMux I__8264 (
            .O(N__39261),
            .I(N__39256));
    InMux I__8263 (
            .O(N__39260),
            .I(N__39251));
    InMux I__8262 (
            .O(N__39259),
            .I(N__39251));
    LocalMux I__8261 (
            .O(N__39256),
            .I(wdtick_cnt_2));
    LocalMux I__8260 (
            .O(N__39251),
            .I(wdtick_cnt_2));
    CascadeMux I__8259 (
            .O(N__39246),
            .I(N__39242));
    InMux I__8258 (
            .O(N__39245),
            .I(N__39237));
    InMux I__8257 (
            .O(N__39242),
            .I(N__39230));
    InMux I__8256 (
            .O(N__39241),
            .I(N__39230));
    InMux I__8255 (
            .O(N__39240),
            .I(N__39230));
    LocalMux I__8254 (
            .O(N__39237),
            .I(wdtick_cnt_0));
    LocalMux I__8253 (
            .O(N__39230),
            .I(wdtick_cnt_0));
    InMux I__8252 (
            .O(N__39225),
            .I(N__39219));
    InMux I__8251 (
            .O(N__39224),
            .I(N__39212));
    InMux I__8250 (
            .O(N__39223),
            .I(N__39212));
    InMux I__8249 (
            .O(N__39222),
            .I(N__39212));
    LocalMux I__8248 (
            .O(N__39219),
            .I(wdtick_cnt_1));
    LocalMux I__8247 (
            .O(N__39212),
            .I(wdtick_cnt_1));
    IoInMux I__8246 (
            .O(N__39207),
            .I(N__39202));
    ClkMux I__8245 (
            .O(N__39206),
            .I(N__39199));
    ClkMux I__8244 (
            .O(N__39205),
            .I(N__39196));
    LocalMux I__8243 (
            .O(N__39202),
            .I(N__39193));
    LocalMux I__8242 (
            .O(N__39199),
            .I(N__39190));
    LocalMux I__8241 (
            .O(N__39196),
            .I(N__39187));
    Span4Mux_s3_v I__8240 (
            .O(N__39193),
            .I(N__39184));
    Span4Mux_v I__8239 (
            .O(N__39190),
            .I(N__39181));
    Span4Mux_v I__8238 (
            .O(N__39187),
            .I(N__39178));
    Sp12to4 I__8237 (
            .O(N__39184),
            .I(N__39175));
    Span4Mux_h I__8236 (
            .O(N__39181),
            .I(N__39172));
    Span4Mux_h I__8235 (
            .O(N__39178),
            .I(N__39169));
    Span12Mux_s10_h I__8234 (
            .O(N__39175),
            .I(N__39165));
    Span4Mux_h I__8233 (
            .O(N__39172),
            .I(N__39162));
    Span4Mux_v I__8232 (
            .O(N__39169),
            .I(N__39159));
    InMux I__8231 (
            .O(N__39168),
            .I(N__39156));
    Odrv12 I__8230 (
            .O(N__39165),
            .I(TEST_LED));
    Odrv4 I__8229 (
            .O(N__39162),
            .I(TEST_LED));
    Odrv4 I__8228 (
            .O(N__39159),
            .I(TEST_LED));
    LocalMux I__8227 (
            .O(N__39156),
            .I(TEST_LED));
    InMux I__8226 (
            .O(N__39147),
            .I(N__39143));
    InMux I__8225 (
            .O(N__39146),
            .I(N__39140));
    LocalMux I__8224 (
            .O(N__39143),
            .I(\comm_spi.n14627 ));
    LocalMux I__8223 (
            .O(N__39140),
            .I(\comm_spi.n14627 ));
    InMux I__8222 (
            .O(N__39135),
            .I(N__39132));
    LocalMux I__8221 (
            .O(N__39132),
            .I(N__39128));
    InMux I__8220 (
            .O(N__39131),
            .I(N__39125));
    Span4Mux_v I__8219 (
            .O(N__39128),
            .I(N__39122));
    LocalMux I__8218 (
            .O(N__39125),
            .I(N__39119));
    Span4Mux_v I__8217 (
            .O(N__39122),
            .I(N__39115));
    Span4Mux_v I__8216 (
            .O(N__39119),
            .I(N__39112));
    InMux I__8215 (
            .O(N__39118),
            .I(N__39109));
    Odrv4 I__8214 (
            .O(N__39115),
            .I(\comm_spi.n22875 ));
    Odrv4 I__8213 (
            .O(N__39112),
            .I(\comm_spi.n22875 ));
    LocalMux I__8212 (
            .O(N__39109),
            .I(\comm_spi.n22875 ));
    InMux I__8211 (
            .O(N__39102),
            .I(N__39099));
    LocalMux I__8210 (
            .O(N__39099),
            .I(N__39096));
    Span4Mux_h I__8209 (
            .O(N__39096),
            .I(N__39092));
    InMux I__8208 (
            .O(N__39095),
            .I(N__39089));
    Span4Mux_v I__8207 (
            .O(N__39092),
            .I(N__39086));
    LocalMux I__8206 (
            .O(N__39089),
            .I(N__39083));
    Odrv4 I__8205 (
            .O(N__39086),
            .I(\comm_spi.n14626 ));
    Odrv12 I__8204 (
            .O(N__39083),
            .I(\comm_spi.n14626 ));
    InMux I__8203 (
            .O(N__39078),
            .I(N__39073));
    InMux I__8202 (
            .O(N__39077),
            .I(N__39070));
    InMux I__8201 (
            .O(N__39076),
            .I(N__39067));
    LocalMux I__8200 (
            .O(N__39073),
            .I(data_index_9));
    LocalMux I__8199 (
            .O(N__39070),
            .I(data_index_9));
    LocalMux I__8198 (
            .O(N__39067),
            .I(data_index_9));
    InMux I__8197 (
            .O(N__39060),
            .I(N__39057));
    LocalMux I__8196 (
            .O(N__39057),
            .I(n8_adj_1559));
    InMux I__8195 (
            .O(N__39054),
            .I(N__39050));
    InMux I__8194 (
            .O(N__39053),
            .I(N__39047));
    LocalMux I__8193 (
            .O(N__39050),
            .I(n7_adj_1558));
    LocalMux I__8192 (
            .O(N__39047),
            .I(n7_adj_1558));
    CascadeMux I__8191 (
            .O(N__39042),
            .I(n8_adj_1559_cascade_));
    CascadeMux I__8190 (
            .O(N__39039),
            .I(N__39036));
    CascadeBuf I__8189 (
            .O(N__39036),
            .I(N__39033));
    CascadeMux I__8188 (
            .O(N__39033),
            .I(N__39030));
    CascadeBuf I__8187 (
            .O(N__39030),
            .I(N__39027));
    CascadeMux I__8186 (
            .O(N__39027),
            .I(N__39024));
    CascadeBuf I__8185 (
            .O(N__39024),
            .I(N__39021));
    CascadeMux I__8184 (
            .O(N__39021),
            .I(N__39018));
    CascadeBuf I__8183 (
            .O(N__39018),
            .I(N__39015));
    CascadeMux I__8182 (
            .O(N__39015),
            .I(N__39012));
    CascadeBuf I__8181 (
            .O(N__39012),
            .I(N__39009));
    CascadeMux I__8180 (
            .O(N__39009),
            .I(N__39006));
    CascadeBuf I__8179 (
            .O(N__39006),
            .I(N__39003));
    CascadeMux I__8178 (
            .O(N__39003),
            .I(N__39000));
    CascadeBuf I__8177 (
            .O(N__39000),
            .I(N__38996));
    CascadeMux I__8176 (
            .O(N__38999),
            .I(N__38993));
    CascadeMux I__8175 (
            .O(N__38996),
            .I(N__38990));
    CascadeBuf I__8174 (
            .O(N__38993),
            .I(N__38987));
    CascadeBuf I__8173 (
            .O(N__38990),
            .I(N__38984));
    CascadeMux I__8172 (
            .O(N__38987),
            .I(N__38981));
    CascadeMux I__8171 (
            .O(N__38984),
            .I(N__38978));
    InMux I__8170 (
            .O(N__38981),
            .I(N__38975));
    CascadeBuf I__8169 (
            .O(N__38978),
            .I(N__38972));
    LocalMux I__8168 (
            .O(N__38975),
            .I(N__38969));
    CascadeMux I__8167 (
            .O(N__38972),
            .I(N__38966));
    Span12Mux_h I__8166 (
            .O(N__38969),
            .I(N__38963));
    InMux I__8165 (
            .O(N__38966),
            .I(N__38960));
    Span12Mux_v I__8164 (
            .O(N__38963),
            .I(N__38955));
    LocalMux I__8163 (
            .O(N__38960),
            .I(N__38955));
    Odrv12 I__8162 (
            .O(N__38955),
            .I(data_index_9_N_216_9));
    InMux I__8161 (
            .O(N__38952),
            .I(N__38948));
    InMux I__8160 (
            .O(N__38951),
            .I(N__38945));
    LocalMux I__8159 (
            .O(N__38948),
            .I(n7_adj_1560));
    LocalMux I__8158 (
            .O(N__38945),
            .I(n7_adj_1560));
    CascadeMux I__8157 (
            .O(N__38940),
            .I(N__38937));
    CascadeBuf I__8156 (
            .O(N__38937),
            .I(N__38934));
    CascadeMux I__8155 (
            .O(N__38934),
            .I(N__38931));
    CascadeBuf I__8154 (
            .O(N__38931),
            .I(N__38928));
    CascadeMux I__8153 (
            .O(N__38928),
            .I(N__38925));
    CascadeBuf I__8152 (
            .O(N__38925),
            .I(N__38922));
    CascadeMux I__8151 (
            .O(N__38922),
            .I(N__38919));
    CascadeBuf I__8150 (
            .O(N__38919),
            .I(N__38916));
    CascadeMux I__8149 (
            .O(N__38916),
            .I(N__38913));
    CascadeBuf I__8148 (
            .O(N__38913),
            .I(N__38910));
    CascadeMux I__8147 (
            .O(N__38910),
            .I(N__38907));
    CascadeBuf I__8146 (
            .O(N__38907),
            .I(N__38904));
    CascadeMux I__8145 (
            .O(N__38904),
            .I(N__38901));
    CascadeBuf I__8144 (
            .O(N__38901),
            .I(N__38897));
    CascadeMux I__8143 (
            .O(N__38900),
            .I(N__38894));
    CascadeMux I__8142 (
            .O(N__38897),
            .I(N__38891));
    CascadeBuf I__8141 (
            .O(N__38894),
            .I(N__38888));
    CascadeBuf I__8140 (
            .O(N__38891),
            .I(N__38885));
    CascadeMux I__8139 (
            .O(N__38888),
            .I(N__38882));
    CascadeMux I__8138 (
            .O(N__38885),
            .I(N__38879));
    InMux I__8137 (
            .O(N__38882),
            .I(N__38876));
    CascadeBuf I__8136 (
            .O(N__38879),
            .I(N__38873));
    LocalMux I__8135 (
            .O(N__38876),
            .I(N__38870));
    CascadeMux I__8134 (
            .O(N__38873),
            .I(N__38867));
    Span12Mux_h I__8133 (
            .O(N__38870),
            .I(N__38864));
    InMux I__8132 (
            .O(N__38867),
            .I(N__38861));
    Span12Mux_v I__8131 (
            .O(N__38864),
            .I(N__38856));
    LocalMux I__8130 (
            .O(N__38861),
            .I(N__38856));
    Odrv12 I__8129 (
            .O(N__38856),
            .I(data_index_9_N_216_8));
    CascadeMux I__8128 (
            .O(N__38853),
            .I(N__38850));
    CascadeBuf I__8127 (
            .O(N__38850),
            .I(N__38847));
    CascadeMux I__8126 (
            .O(N__38847),
            .I(N__38844));
    CascadeBuf I__8125 (
            .O(N__38844),
            .I(N__38841));
    CascadeMux I__8124 (
            .O(N__38841),
            .I(N__38838));
    CascadeBuf I__8123 (
            .O(N__38838),
            .I(N__38835));
    CascadeMux I__8122 (
            .O(N__38835),
            .I(N__38832));
    CascadeBuf I__8121 (
            .O(N__38832),
            .I(N__38829));
    CascadeMux I__8120 (
            .O(N__38829),
            .I(N__38826));
    CascadeBuf I__8119 (
            .O(N__38826),
            .I(N__38823));
    CascadeMux I__8118 (
            .O(N__38823),
            .I(N__38820));
    CascadeBuf I__8117 (
            .O(N__38820),
            .I(N__38817));
    CascadeMux I__8116 (
            .O(N__38817),
            .I(N__38814));
    CascadeBuf I__8115 (
            .O(N__38814),
            .I(N__38810));
    CascadeMux I__8114 (
            .O(N__38813),
            .I(N__38807));
    CascadeMux I__8113 (
            .O(N__38810),
            .I(N__38804));
    CascadeBuf I__8112 (
            .O(N__38807),
            .I(N__38801));
    CascadeBuf I__8111 (
            .O(N__38804),
            .I(N__38798));
    CascadeMux I__8110 (
            .O(N__38801),
            .I(N__38795));
    CascadeMux I__8109 (
            .O(N__38798),
            .I(N__38792));
    InMux I__8108 (
            .O(N__38795),
            .I(N__38789));
    CascadeBuf I__8107 (
            .O(N__38792),
            .I(N__38786));
    LocalMux I__8106 (
            .O(N__38789),
            .I(N__38783));
    CascadeMux I__8105 (
            .O(N__38786),
            .I(N__38780));
    Span12Mux_h I__8104 (
            .O(N__38783),
            .I(N__38777));
    InMux I__8103 (
            .O(N__38780),
            .I(N__38774));
    Span12Mux_v I__8102 (
            .O(N__38777),
            .I(N__38769));
    LocalMux I__8101 (
            .O(N__38774),
            .I(N__38769));
    Odrv12 I__8100 (
            .O(N__38769),
            .I(data_index_9_N_216_7));
    InMux I__8099 (
            .O(N__38766),
            .I(N__38762));
    InMux I__8098 (
            .O(N__38765),
            .I(N__38759));
    LocalMux I__8097 (
            .O(N__38762),
            .I(N__38756));
    LocalMux I__8096 (
            .O(N__38759),
            .I(N__38742));
    Glb2LocalMux I__8095 (
            .O(N__38756),
            .I(N__38706));
    ClkMux I__8094 (
            .O(N__38755),
            .I(N__38706));
    ClkMux I__8093 (
            .O(N__38754),
            .I(N__38706));
    ClkMux I__8092 (
            .O(N__38753),
            .I(N__38706));
    ClkMux I__8091 (
            .O(N__38752),
            .I(N__38706));
    ClkMux I__8090 (
            .O(N__38751),
            .I(N__38706));
    ClkMux I__8089 (
            .O(N__38750),
            .I(N__38706));
    ClkMux I__8088 (
            .O(N__38749),
            .I(N__38706));
    ClkMux I__8087 (
            .O(N__38748),
            .I(N__38706));
    ClkMux I__8086 (
            .O(N__38747),
            .I(N__38706));
    ClkMux I__8085 (
            .O(N__38746),
            .I(N__38706));
    ClkMux I__8084 (
            .O(N__38745),
            .I(N__38706));
    Glb2LocalMux I__8083 (
            .O(N__38742),
            .I(N__38706));
    ClkMux I__8082 (
            .O(N__38741),
            .I(N__38706));
    ClkMux I__8081 (
            .O(N__38740),
            .I(N__38706));
    ClkMux I__8080 (
            .O(N__38739),
            .I(N__38706));
    GlobalMux I__8079 (
            .O(N__38706),
            .I(clk_16MHz));
    InMux I__8078 (
            .O(N__38703),
            .I(N__38700));
    LocalMux I__8077 (
            .O(N__38700),
            .I(N__38697));
    Span4Mux_v I__8076 (
            .O(N__38697),
            .I(N__38694));
    Span4Mux_v I__8075 (
            .O(N__38694),
            .I(N__38691));
    Span4Mux_v I__8074 (
            .O(N__38691),
            .I(N__38687));
    InMux I__8073 (
            .O(N__38690),
            .I(N__38684));
    Odrv4 I__8072 (
            .O(N__38687),
            .I(dds0_mclk));
    LocalMux I__8071 (
            .O(N__38684),
            .I(dds0_mclk));
    InMux I__8070 (
            .O(N__38679),
            .I(N__38676));
    LocalMux I__8069 (
            .O(N__38676),
            .I(N__38671));
    CascadeMux I__8068 (
            .O(N__38675),
            .I(N__38668));
    InMux I__8067 (
            .O(N__38674),
            .I(N__38665));
    Span4Mux_v I__8066 (
            .O(N__38671),
            .I(N__38662));
    InMux I__8065 (
            .O(N__38668),
            .I(N__38659));
    LocalMux I__8064 (
            .O(N__38665),
            .I(N__38656));
    Odrv4 I__8063 (
            .O(N__38662),
            .I(buf_control_6));
    LocalMux I__8062 (
            .O(N__38659),
            .I(buf_control_6));
    Odrv4 I__8061 (
            .O(N__38656),
            .I(buf_control_6));
    IoInMux I__8060 (
            .O(N__38649),
            .I(N__38646));
    LocalMux I__8059 (
            .O(N__38646),
            .I(N__38643));
    Span4Mux_s2_v I__8058 (
            .O(N__38643),
            .I(N__38640));
    Span4Mux_h I__8057 (
            .O(N__38640),
            .I(N__38637));
    Span4Mux_h I__8056 (
            .O(N__38637),
            .I(N__38634));
    Span4Mux_v I__8055 (
            .O(N__38634),
            .I(N__38631));
    Odrv4 I__8054 (
            .O(N__38631),
            .I(DDS_MCLK));
    InMux I__8053 (
            .O(N__38628),
            .I(N__38625));
    LocalMux I__8052 (
            .O(N__38625),
            .I(N__38622));
    Span4Mux_v I__8051 (
            .O(N__38622),
            .I(N__38619));
    Span4Mux_v I__8050 (
            .O(N__38619),
            .I(N__38615));
    InMux I__8049 (
            .O(N__38618),
            .I(N__38612));
    Odrv4 I__8048 (
            .O(N__38615),
            .I(\comm_spi.n14619 ));
    LocalMux I__8047 (
            .O(N__38612),
            .I(\comm_spi.n14619 ));
    InMux I__8046 (
            .O(N__38607),
            .I(N__38603));
    InMux I__8045 (
            .O(N__38606),
            .I(N__38600));
    LocalMux I__8044 (
            .O(N__38603),
            .I(\comm_spi.n22884 ));
    LocalMux I__8043 (
            .O(N__38600),
            .I(\comm_spi.n22884 ));
    CascadeMux I__8042 (
            .O(N__38595),
            .I(\comm_spi.n22884_cascade_ ));
    InMux I__8041 (
            .O(N__38592),
            .I(N__38588));
    InMux I__8040 (
            .O(N__38591),
            .I(N__38585));
    LocalMux I__8039 (
            .O(N__38588),
            .I(\comm_spi.n14593 ));
    LocalMux I__8038 (
            .O(N__38585),
            .I(\comm_spi.n14593 ));
    InMux I__8037 (
            .O(N__38580),
            .I(N__38577));
    LocalMux I__8036 (
            .O(N__38577),
            .I(N__38574));
    Span4Mux_v I__8035 (
            .O(N__38574),
            .I(N__38570));
    InMux I__8034 (
            .O(N__38573),
            .I(N__38567));
    Span4Mux_v I__8033 (
            .O(N__38570),
            .I(N__38562));
    LocalMux I__8032 (
            .O(N__38567),
            .I(N__38562));
    Odrv4 I__8031 (
            .O(N__38562),
            .I(\comm_spi.n14618 ));
    CEMux I__8030 (
            .O(N__38559),
            .I(N__38553));
    CEMux I__8029 (
            .O(N__38558),
            .I(N__38549));
    CEMux I__8028 (
            .O(N__38557),
            .I(N__38546));
    InMux I__8027 (
            .O(N__38556),
            .I(N__38543));
    LocalMux I__8026 (
            .O(N__38553),
            .I(N__38540));
    CEMux I__8025 (
            .O(N__38552),
            .I(N__38537));
    LocalMux I__8024 (
            .O(N__38549),
            .I(N__38534));
    LocalMux I__8023 (
            .O(N__38546),
            .I(N__38531));
    LocalMux I__8022 (
            .O(N__38543),
            .I(N__38528));
    Span4Mux_v I__8021 (
            .O(N__38540),
            .I(N__38525));
    LocalMux I__8020 (
            .O(N__38537),
            .I(N__38522));
    Span4Mux_h I__8019 (
            .O(N__38534),
            .I(N__38519));
    Span4Mux_h I__8018 (
            .O(N__38531),
            .I(N__38516));
    Span4Mux_h I__8017 (
            .O(N__38528),
            .I(N__38513));
    Span4Mux_h I__8016 (
            .O(N__38525),
            .I(N__38508));
    Span4Mux_v I__8015 (
            .O(N__38522),
            .I(N__38508));
    Span4Mux_v I__8014 (
            .O(N__38519),
            .I(N__38501));
    Span4Mux_v I__8013 (
            .O(N__38516),
            .I(N__38501));
    Span4Mux_v I__8012 (
            .O(N__38513),
            .I(N__38501));
    Odrv4 I__8011 (
            .O(N__38508),
            .I(n13457));
    Odrv4 I__8010 (
            .O(N__38501),
            .I(n13457));
    SRMux I__8009 (
            .O(N__38496),
            .I(N__38493));
    LocalMux I__8008 (
            .O(N__38493),
            .I(N__38490));
    Span4Mux_v I__8007 (
            .O(N__38490),
            .I(N__38486));
    SRMux I__8006 (
            .O(N__38489),
            .I(N__38483));
    Span4Mux_h I__8005 (
            .O(N__38486),
            .I(N__38476));
    LocalMux I__8004 (
            .O(N__38483),
            .I(N__38476));
    SRMux I__8003 (
            .O(N__38482),
            .I(N__38473));
    SRMux I__8002 (
            .O(N__38481),
            .I(N__38470));
    Span4Mux_v I__8001 (
            .O(N__38476),
            .I(N__38465));
    LocalMux I__8000 (
            .O(N__38473),
            .I(N__38465));
    LocalMux I__7999 (
            .O(N__38470),
            .I(N__38462));
    Span4Mux_h I__7998 (
            .O(N__38465),
            .I(N__38459));
    Span4Mux_v I__7997 (
            .O(N__38462),
            .I(N__38456));
    Odrv4 I__7996 (
            .O(N__38459),
            .I(n14647));
    Odrv4 I__7995 (
            .O(N__38456),
            .I(n14647));
    CascadeMux I__7994 (
            .O(N__38451),
            .I(N__38447));
    InMux I__7993 (
            .O(N__38450),
            .I(N__38444));
    InMux I__7992 (
            .O(N__38447),
            .I(N__38441));
    LocalMux I__7991 (
            .O(N__38444),
            .I(N__38438));
    LocalMux I__7990 (
            .O(N__38441),
            .I(acadc_skipcnt_0));
    Odrv12 I__7989 (
            .O(N__38438),
            .I(acadc_skipcnt_0));
    CascadeMux I__7988 (
            .O(N__38433),
            .I(N__38430));
    InMux I__7987 (
            .O(N__38430),
            .I(N__38427));
    LocalMux I__7986 (
            .O(N__38427),
            .I(N__38423));
    InMux I__7985 (
            .O(N__38426),
            .I(N__38420));
    Span4Mux_h I__7984 (
            .O(N__38423),
            .I(N__38417));
    LocalMux I__7983 (
            .O(N__38420),
            .I(acadc_skipcnt_6));
    Odrv4 I__7982 (
            .O(N__38417),
            .I(acadc_skipcnt_6));
    InMux I__7981 (
            .O(N__38412),
            .I(N__38409));
    LocalMux I__7980 (
            .O(N__38409),
            .I(N__38406));
    Span4Mux_v I__7979 (
            .O(N__38406),
            .I(N__38403));
    Span4Mux_h I__7978 (
            .O(N__38403),
            .I(N__38400));
    Odrv4 I__7977 (
            .O(N__38400),
            .I(n17));
    CascadeMux I__7976 (
            .O(N__38397),
            .I(n8_adj_1565_cascade_));
    InMux I__7975 (
            .O(N__38394),
            .I(N__38389));
    InMux I__7974 (
            .O(N__38393),
            .I(N__38386));
    InMux I__7973 (
            .O(N__38392),
            .I(N__38383));
    LocalMux I__7972 (
            .O(N__38389),
            .I(data_index_6));
    LocalMux I__7971 (
            .O(N__38386),
            .I(data_index_6));
    LocalMux I__7970 (
            .O(N__38383),
            .I(data_index_6));
    CascadeMux I__7969 (
            .O(N__38376),
            .I(N__38373));
    CascadeBuf I__7968 (
            .O(N__38373),
            .I(N__38370));
    CascadeMux I__7967 (
            .O(N__38370),
            .I(N__38367));
    CascadeBuf I__7966 (
            .O(N__38367),
            .I(N__38364));
    CascadeMux I__7965 (
            .O(N__38364),
            .I(N__38361));
    CascadeBuf I__7964 (
            .O(N__38361),
            .I(N__38358));
    CascadeMux I__7963 (
            .O(N__38358),
            .I(N__38355));
    CascadeBuf I__7962 (
            .O(N__38355),
            .I(N__38352));
    CascadeMux I__7961 (
            .O(N__38352),
            .I(N__38349));
    CascadeBuf I__7960 (
            .O(N__38349),
            .I(N__38346));
    CascadeMux I__7959 (
            .O(N__38346),
            .I(N__38343));
    CascadeBuf I__7958 (
            .O(N__38343),
            .I(N__38340));
    CascadeMux I__7957 (
            .O(N__38340),
            .I(N__38337));
    CascadeBuf I__7956 (
            .O(N__38337),
            .I(N__38334));
    CascadeMux I__7955 (
            .O(N__38334),
            .I(N__38331));
    CascadeBuf I__7954 (
            .O(N__38331),
            .I(N__38327));
    CascadeMux I__7953 (
            .O(N__38330),
            .I(N__38324));
    CascadeMux I__7952 (
            .O(N__38327),
            .I(N__38321));
    CascadeBuf I__7951 (
            .O(N__38324),
            .I(N__38318));
    CascadeBuf I__7950 (
            .O(N__38321),
            .I(N__38315));
    CascadeMux I__7949 (
            .O(N__38318),
            .I(N__38312));
    CascadeMux I__7948 (
            .O(N__38315),
            .I(N__38309));
    InMux I__7947 (
            .O(N__38312),
            .I(N__38306));
    InMux I__7946 (
            .O(N__38309),
            .I(N__38303));
    LocalMux I__7945 (
            .O(N__38306),
            .I(N__38300));
    LocalMux I__7944 (
            .O(N__38303),
            .I(N__38297));
    Sp12to4 I__7943 (
            .O(N__38300),
            .I(N__38294));
    Span4Mux_h I__7942 (
            .O(N__38297),
            .I(N__38291));
    Span12Mux_v I__7941 (
            .O(N__38294),
            .I(N__38288));
    Span4Mux_h I__7940 (
            .O(N__38291),
            .I(N__38285));
    Odrv12 I__7939 (
            .O(N__38288),
            .I(data_index_9_N_216_3));
    Odrv4 I__7938 (
            .O(N__38285),
            .I(data_index_9_N_216_3));
    CascadeMux I__7937 (
            .O(N__38280),
            .I(N__38277));
    InMux I__7936 (
            .O(N__38277),
            .I(N__38274));
    LocalMux I__7935 (
            .O(N__38274),
            .I(N__38271));
    Odrv4 I__7934 (
            .O(N__38271),
            .I(n8_adj_1565));
    InMux I__7933 (
            .O(N__38268),
            .I(N__38264));
    InMux I__7932 (
            .O(N__38267),
            .I(N__38261));
    LocalMux I__7931 (
            .O(N__38264),
            .I(n7_adj_1564));
    LocalMux I__7930 (
            .O(N__38261),
            .I(n7_adj_1564));
    CascadeMux I__7929 (
            .O(N__38256),
            .I(N__38253));
    CascadeBuf I__7928 (
            .O(N__38253),
            .I(N__38250));
    CascadeMux I__7927 (
            .O(N__38250),
            .I(N__38247));
    CascadeBuf I__7926 (
            .O(N__38247),
            .I(N__38244));
    CascadeMux I__7925 (
            .O(N__38244),
            .I(N__38241));
    CascadeBuf I__7924 (
            .O(N__38241),
            .I(N__38238));
    CascadeMux I__7923 (
            .O(N__38238),
            .I(N__38235));
    CascadeBuf I__7922 (
            .O(N__38235),
            .I(N__38232));
    CascadeMux I__7921 (
            .O(N__38232),
            .I(N__38229));
    CascadeBuf I__7920 (
            .O(N__38229),
            .I(N__38226));
    CascadeMux I__7919 (
            .O(N__38226),
            .I(N__38223));
    CascadeBuf I__7918 (
            .O(N__38223),
            .I(N__38220));
    CascadeMux I__7917 (
            .O(N__38220),
            .I(N__38217));
    CascadeBuf I__7916 (
            .O(N__38217),
            .I(N__38214));
    CascadeMux I__7915 (
            .O(N__38214),
            .I(N__38210));
    CascadeMux I__7914 (
            .O(N__38213),
            .I(N__38207));
    CascadeBuf I__7913 (
            .O(N__38210),
            .I(N__38204));
    CascadeBuf I__7912 (
            .O(N__38207),
            .I(N__38201));
    CascadeMux I__7911 (
            .O(N__38204),
            .I(N__38198));
    CascadeMux I__7910 (
            .O(N__38201),
            .I(N__38195));
    CascadeBuf I__7909 (
            .O(N__38198),
            .I(N__38192));
    InMux I__7908 (
            .O(N__38195),
            .I(N__38189));
    CascadeMux I__7907 (
            .O(N__38192),
            .I(N__38186));
    LocalMux I__7906 (
            .O(N__38189),
            .I(N__38183));
    InMux I__7905 (
            .O(N__38186),
            .I(N__38180));
    Span12Mux_h I__7904 (
            .O(N__38183),
            .I(N__38177));
    LocalMux I__7903 (
            .O(N__38180),
            .I(N__38174));
    Span12Mux_v I__7902 (
            .O(N__38177),
            .I(N__38171));
    Span4Mux_h I__7901 (
            .O(N__38174),
            .I(N__38168));
    Odrv12 I__7900 (
            .O(N__38171),
            .I(data_index_9_N_216_6));
    Odrv4 I__7899 (
            .O(N__38168),
            .I(data_index_9_N_216_6));
    InMux I__7898 (
            .O(N__38163),
            .I(n19601));
    InMux I__7897 (
            .O(N__38160),
            .I(bfn_15_17_0_));
    InMux I__7896 (
            .O(N__38157),
            .I(n19603));
    InMux I__7895 (
            .O(N__38154),
            .I(n19604));
    InMux I__7894 (
            .O(N__38151),
            .I(n19605));
    InMux I__7893 (
            .O(N__38148),
            .I(N__38145));
    LocalMux I__7892 (
            .O(N__38145),
            .I(N__38141));
    InMux I__7891 (
            .O(N__38144),
            .I(N__38138));
    Span4Mux_h I__7890 (
            .O(N__38141),
            .I(N__38135));
    LocalMux I__7889 (
            .O(N__38138),
            .I(data_cntvec_12));
    Odrv4 I__7888 (
            .O(N__38135),
            .I(data_cntvec_12));
    InMux I__7887 (
            .O(N__38130),
            .I(n19606));
    InMux I__7886 (
            .O(N__38127),
            .I(N__38124));
    LocalMux I__7885 (
            .O(N__38124),
            .I(N__38120));
    InMux I__7884 (
            .O(N__38123),
            .I(N__38117));
    Span4Mux_v I__7883 (
            .O(N__38120),
            .I(N__38114));
    LocalMux I__7882 (
            .O(N__38117),
            .I(data_cntvec_13));
    Odrv4 I__7881 (
            .O(N__38114),
            .I(data_cntvec_13));
    InMux I__7880 (
            .O(N__38109),
            .I(n19607));
    InMux I__7879 (
            .O(N__38106),
            .I(N__38102));
    InMux I__7878 (
            .O(N__38105),
            .I(N__38099));
    LocalMux I__7877 (
            .O(N__38102),
            .I(data_cntvec_14));
    LocalMux I__7876 (
            .O(N__38099),
            .I(data_cntvec_14));
    InMux I__7875 (
            .O(N__38094),
            .I(n19608));
    InMux I__7874 (
            .O(N__38091),
            .I(n19609));
    InMux I__7873 (
            .O(N__38088),
            .I(N__38085));
    LocalMux I__7872 (
            .O(N__38085),
            .I(N__38081));
    InMux I__7871 (
            .O(N__38084),
            .I(N__38078));
    Span4Mux_h I__7870 (
            .O(N__38081),
            .I(N__38075));
    LocalMux I__7869 (
            .O(N__38078),
            .I(data_cntvec_15));
    Odrv4 I__7868 (
            .O(N__38075),
            .I(data_cntvec_15));
    InMux I__7867 (
            .O(N__38070),
            .I(N__38066));
    InMux I__7866 (
            .O(N__38069),
            .I(N__38063));
    LocalMux I__7865 (
            .O(N__38066),
            .I(N__38058));
    LocalMux I__7864 (
            .O(N__38063),
            .I(N__38058));
    Span4Mux_h I__7863 (
            .O(N__38058),
            .I(N__38055));
    Span4Mux_v I__7862 (
            .O(N__38055),
            .I(N__38052));
    Odrv4 I__7861 (
            .O(N__38052),
            .I(n14_adj_1576));
    CascadeMux I__7860 (
            .O(N__38049),
            .I(N__38045));
    InMux I__7859 (
            .O(N__38048),
            .I(N__38042));
    InMux I__7858 (
            .O(N__38045),
            .I(N__38039));
    LocalMux I__7857 (
            .O(N__38042),
            .I(N__38036));
    LocalMux I__7856 (
            .O(N__38039),
            .I(data_idxvec_14));
    Odrv12 I__7855 (
            .O(N__38036),
            .I(data_idxvec_14));
    InMux I__7854 (
            .O(N__38031),
            .I(n19647));
    InMux I__7853 (
            .O(N__38028),
            .I(N__38025));
    LocalMux I__7852 (
            .O(N__38025),
            .I(N__38022));
    Span4Mux_v I__7851 (
            .O(N__38022),
            .I(N__38019));
    Span4Mux_h I__7850 (
            .O(N__38019),
            .I(N__38015));
    InMux I__7849 (
            .O(N__38018),
            .I(N__38012));
    Odrv4 I__7848 (
            .O(N__38015),
            .I(n14_adj_1549));
    LocalMux I__7847 (
            .O(N__38012),
            .I(n14_adj_1549));
    InMux I__7846 (
            .O(N__38007),
            .I(n19648));
    InMux I__7845 (
            .O(N__38004),
            .I(N__38001));
    LocalMux I__7844 (
            .O(N__38001),
            .I(N__37997));
    InMux I__7843 (
            .O(N__38000),
            .I(N__37994));
    Span4Mux_h I__7842 (
            .O(N__37997),
            .I(N__37991));
    LocalMux I__7841 (
            .O(N__37994),
            .I(data_idxvec_15));
    Odrv4 I__7840 (
            .O(N__37991),
            .I(data_idxvec_15));
    CEMux I__7839 (
            .O(N__37986),
            .I(N__37983));
    LocalMux I__7838 (
            .O(N__37983),
            .I(N__37979));
    CEMux I__7837 (
            .O(N__37982),
            .I(N__37976));
    Span4Mux_v I__7836 (
            .O(N__37979),
            .I(N__37971));
    LocalMux I__7835 (
            .O(N__37976),
            .I(N__37971));
    Span4Mux_v I__7834 (
            .O(N__37971),
            .I(N__37968));
    Span4Mux_v I__7833 (
            .O(N__37968),
            .I(N__37965));
    Odrv4 I__7832 (
            .O(N__37965),
            .I(n12280));
    CascadeMux I__7831 (
            .O(N__37962),
            .I(N__37959));
    InMux I__7830 (
            .O(N__37959),
            .I(N__37955));
    InMux I__7829 (
            .O(N__37958),
            .I(N__37950));
    LocalMux I__7828 (
            .O(N__37955),
            .I(N__37947));
    InMux I__7827 (
            .O(N__37954),
            .I(N__37944));
    InMux I__7826 (
            .O(N__37953),
            .I(N__37941));
    LocalMux I__7825 (
            .O(N__37950),
            .I(N__37934));
    Span4Mux_h I__7824 (
            .O(N__37947),
            .I(N__37934));
    LocalMux I__7823 (
            .O(N__37944),
            .I(N__37934));
    LocalMux I__7822 (
            .O(N__37941),
            .I(N__37931));
    Span4Mux_v I__7821 (
            .O(N__37934),
            .I(N__37928));
    Odrv4 I__7820 (
            .O(N__37931),
            .I(iac_raw_buf_N_736));
    Odrv4 I__7819 (
            .O(N__37928),
            .I(iac_raw_buf_N_736));
    InMux I__7818 (
            .O(N__37923),
            .I(N__37920));
    LocalMux I__7817 (
            .O(N__37920),
            .I(N__37915));
    InMux I__7816 (
            .O(N__37919),
            .I(N__37912));
    InMux I__7815 (
            .O(N__37918),
            .I(N__37909));
    Span4Mux_v I__7814 (
            .O(N__37915),
            .I(N__37906));
    LocalMux I__7813 (
            .O(N__37912),
            .I(data_cntvec_1));
    LocalMux I__7812 (
            .O(N__37909),
            .I(data_cntvec_1));
    Odrv4 I__7811 (
            .O(N__37906),
            .I(data_cntvec_1));
    InMux I__7810 (
            .O(N__37899),
            .I(n19595));
    InMux I__7809 (
            .O(N__37896),
            .I(n19596));
    InMux I__7808 (
            .O(N__37893),
            .I(n19597));
    InMux I__7807 (
            .O(N__37890),
            .I(n19598));
    InMux I__7806 (
            .O(N__37887),
            .I(n19599));
    InMux I__7805 (
            .O(N__37884),
            .I(n19600));
    InMux I__7804 (
            .O(N__37881),
            .I(n19639));
    InMux I__7803 (
            .O(N__37878),
            .I(N__37874));
    InMux I__7802 (
            .O(N__37877),
            .I(N__37871));
    LocalMux I__7801 (
            .O(N__37874),
            .I(N__37866));
    LocalMux I__7800 (
            .O(N__37871),
            .I(N__37866));
    Span4Mux_v I__7799 (
            .O(N__37866),
            .I(N__37863));
    Span4Mux_h I__7798 (
            .O(N__37863),
            .I(N__37860));
    Span4Mux_h I__7797 (
            .O(N__37860),
            .I(N__37857));
    Odrv4 I__7796 (
            .O(N__37857),
            .I(n14_adj_1551));
    InMux I__7795 (
            .O(N__37854),
            .I(n19640));
    InMux I__7794 (
            .O(N__37851),
            .I(N__37848));
    LocalMux I__7793 (
            .O(N__37848),
            .I(N__37844));
    InMux I__7792 (
            .O(N__37847),
            .I(N__37841));
    Span4Mux_h I__7791 (
            .O(N__37844),
            .I(N__37836));
    LocalMux I__7790 (
            .O(N__37841),
            .I(N__37836));
    Span4Mux_v I__7789 (
            .O(N__37836),
            .I(N__37833));
    Odrv4 I__7788 (
            .O(N__37833),
            .I(n14_adj_1550));
    InMux I__7787 (
            .O(N__37830),
            .I(bfn_15_15_0_));
    InMux I__7786 (
            .O(N__37827),
            .I(N__37824));
    LocalMux I__7785 (
            .O(N__37824),
            .I(N__37820));
    InMux I__7784 (
            .O(N__37823),
            .I(N__37817));
    Span4Mux_v I__7783 (
            .O(N__37820),
            .I(N__37814));
    LocalMux I__7782 (
            .O(N__37817),
            .I(N__37811));
    Span4Mux_v I__7781 (
            .O(N__37814),
            .I(N__37808));
    Sp12to4 I__7780 (
            .O(N__37811),
            .I(N__37805));
    Sp12to4 I__7779 (
            .O(N__37808),
            .I(N__37800));
    Span12Mux_v I__7778 (
            .O(N__37805),
            .I(N__37800));
    Odrv12 I__7777 (
            .O(N__37800),
            .I(n14_adj_1580));
    InMux I__7776 (
            .O(N__37797),
            .I(n19642));
    InMux I__7775 (
            .O(N__37794),
            .I(N__37791));
    LocalMux I__7774 (
            .O(N__37791),
            .I(N__37787));
    InMux I__7773 (
            .O(N__37790),
            .I(N__37784));
    Span4Mux_v I__7772 (
            .O(N__37787),
            .I(N__37781));
    LocalMux I__7771 (
            .O(N__37784),
            .I(n14_adj_1579));
    Odrv4 I__7770 (
            .O(N__37781),
            .I(n14_adj_1579));
    InMux I__7769 (
            .O(N__37776),
            .I(n19643));
    InMux I__7768 (
            .O(N__37773),
            .I(n19644));
    InMux I__7767 (
            .O(N__37770),
            .I(N__37766));
    InMux I__7766 (
            .O(N__37769),
            .I(N__37763));
    LocalMux I__7765 (
            .O(N__37766),
            .I(N__37760));
    LocalMux I__7764 (
            .O(N__37763),
            .I(N__37757));
    Span4Mux_h I__7763 (
            .O(N__37760),
            .I(N__37754));
    Odrv4 I__7762 (
            .O(N__37757),
            .I(n14_adj_1577));
    Odrv4 I__7761 (
            .O(N__37754),
            .I(n14_adj_1577));
    CascadeMux I__7760 (
            .O(N__37749),
            .I(N__37745));
    InMux I__7759 (
            .O(N__37748),
            .I(N__37742));
    InMux I__7758 (
            .O(N__37745),
            .I(N__37739));
    LocalMux I__7757 (
            .O(N__37742),
            .I(N__37736));
    LocalMux I__7756 (
            .O(N__37739),
            .I(data_idxvec_12));
    Odrv4 I__7755 (
            .O(N__37736),
            .I(data_idxvec_12));
    InMux I__7754 (
            .O(N__37731),
            .I(n19645));
    InMux I__7753 (
            .O(N__37728),
            .I(N__37724));
    InMux I__7752 (
            .O(N__37727),
            .I(N__37721));
    LocalMux I__7751 (
            .O(N__37724),
            .I(N__37718));
    LocalMux I__7750 (
            .O(N__37721),
            .I(N__37714));
    Span4Mux_v I__7749 (
            .O(N__37718),
            .I(N__37711));
    InMux I__7748 (
            .O(N__37717),
            .I(N__37708));
    Span4Mux_h I__7747 (
            .O(N__37714),
            .I(N__37705));
    Odrv4 I__7746 (
            .O(N__37711),
            .I(n14_adj_1583));
    LocalMux I__7745 (
            .O(N__37708),
            .I(n14_adj_1583));
    Odrv4 I__7744 (
            .O(N__37705),
            .I(n14_adj_1583));
    CascadeMux I__7743 (
            .O(N__37698),
            .I(N__37695));
    InMux I__7742 (
            .O(N__37695),
            .I(N__37691));
    CascadeMux I__7741 (
            .O(N__37694),
            .I(N__37688));
    LocalMux I__7740 (
            .O(N__37691),
            .I(N__37685));
    InMux I__7739 (
            .O(N__37688),
            .I(N__37682));
    Span4Mux_h I__7738 (
            .O(N__37685),
            .I(N__37679));
    LocalMux I__7737 (
            .O(N__37682),
            .I(data_idxvec_13));
    Odrv4 I__7736 (
            .O(N__37679),
            .I(data_idxvec_13));
    InMux I__7735 (
            .O(N__37674),
            .I(n19646));
    CascadeMux I__7734 (
            .O(N__37671),
            .I(N__37668));
    InMux I__7733 (
            .O(N__37668),
            .I(N__37665));
    LocalMux I__7732 (
            .O(N__37665),
            .I(N__37662));
    Span4Mux_h I__7731 (
            .O(N__37662),
            .I(N__37659));
    Odrv4 I__7730 (
            .O(N__37659),
            .I(n26_adj_1644));
    InMux I__7729 (
            .O(N__37656),
            .I(N__37653));
    LocalMux I__7728 (
            .O(N__37653),
            .I(N__37649));
    InMux I__7727 (
            .O(N__37652),
            .I(N__37646));
    Span4Mux_h I__7726 (
            .O(N__37649),
            .I(N__37639));
    LocalMux I__7725 (
            .O(N__37646),
            .I(N__37639));
    InMux I__7724 (
            .O(N__37645),
            .I(N__37636));
    InMux I__7723 (
            .O(N__37644),
            .I(N__37633));
    Odrv4 I__7722 (
            .O(N__37639),
            .I(n20893));
    LocalMux I__7721 (
            .O(N__37636),
            .I(n20893));
    LocalMux I__7720 (
            .O(N__37633),
            .I(n20893));
    InMux I__7719 (
            .O(N__37626),
            .I(N__37623));
    LocalMux I__7718 (
            .O(N__37623),
            .I(N__37620));
    Span4Mux_v I__7717 (
            .O(N__37620),
            .I(N__37617));
    Odrv4 I__7716 (
            .O(N__37617),
            .I(n21521));
    InMux I__7715 (
            .O(N__37614),
            .I(N__37610));
    InMux I__7714 (
            .O(N__37613),
            .I(N__37607));
    LocalMux I__7713 (
            .O(N__37610),
            .I(n14_adj_1533));
    LocalMux I__7712 (
            .O(N__37607),
            .I(n14_adj_1533));
    InMux I__7711 (
            .O(N__37602),
            .I(bfn_15_14_0_));
    InMux I__7710 (
            .O(N__37599),
            .I(N__37596));
    LocalMux I__7709 (
            .O(N__37596),
            .I(N__37593));
    Span4Mux_v I__7708 (
            .O(N__37593),
            .I(N__37590));
    Span4Mux_h I__7707 (
            .O(N__37590),
            .I(N__37586));
    InMux I__7706 (
            .O(N__37589),
            .I(N__37583));
    Span4Mux_v I__7705 (
            .O(N__37586),
            .I(N__37580));
    LocalMux I__7704 (
            .O(N__37583),
            .I(n14_adj_1556));
    Odrv4 I__7703 (
            .O(N__37580),
            .I(n14_adj_1556));
    CascadeMux I__7702 (
            .O(N__37575),
            .I(N__37571));
    CascadeMux I__7701 (
            .O(N__37574),
            .I(N__37568));
    InMux I__7700 (
            .O(N__37571),
            .I(N__37565));
    InMux I__7699 (
            .O(N__37568),
            .I(N__37562));
    LocalMux I__7698 (
            .O(N__37565),
            .I(N__37559));
    LocalMux I__7697 (
            .O(N__37562),
            .I(data_idxvec_1));
    Odrv4 I__7696 (
            .O(N__37559),
            .I(data_idxvec_1));
    InMux I__7695 (
            .O(N__37554),
            .I(n19634));
    InMux I__7694 (
            .O(N__37551),
            .I(N__37548));
    LocalMux I__7693 (
            .O(N__37548),
            .I(N__37544));
    InMux I__7692 (
            .O(N__37547),
            .I(N__37541));
    Span4Mux_h I__7691 (
            .O(N__37544),
            .I(N__37538));
    LocalMux I__7690 (
            .O(N__37541),
            .I(n14_adj_1555));
    Odrv4 I__7689 (
            .O(N__37538),
            .I(n14_adj_1555));
    InMux I__7688 (
            .O(N__37533),
            .I(n19635));
    InMux I__7687 (
            .O(N__37530),
            .I(n19636));
    InMux I__7686 (
            .O(N__37527),
            .I(N__37523));
    InMux I__7685 (
            .O(N__37526),
            .I(N__37520));
    LocalMux I__7684 (
            .O(N__37523),
            .I(N__37517));
    LocalMux I__7683 (
            .O(N__37520),
            .I(N__37514));
    Span4Mux_h I__7682 (
            .O(N__37517),
            .I(N__37511));
    Span12Mux_h I__7681 (
            .O(N__37514),
            .I(N__37508));
    Span4Mux_h I__7680 (
            .O(N__37511),
            .I(N__37505));
    Odrv12 I__7679 (
            .O(N__37508),
            .I(n14_adj_1553));
    Odrv4 I__7678 (
            .O(N__37505),
            .I(n14_adj_1553));
    InMux I__7677 (
            .O(N__37500),
            .I(n19637));
    InMux I__7676 (
            .O(N__37497),
            .I(N__37493));
    CascadeMux I__7675 (
            .O(N__37496),
            .I(N__37490));
    LocalMux I__7674 (
            .O(N__37493),
            .I(N__37487));
    InMux I__7673 (
            .O(N__37490),
            .I(N__37483));
    Span4Mux_v I__7672 (
            .O(N__37487),
            .I(N__37480));
    InMux I__7671 (
            .O(N__37486),
            .I(N__37477));
    LocalMux I__7670 (
            .O(N__37483),
            .I(n14_adj_1584));
    Odrv4 I__7669 (
            .O(N__37480),
            .I(n14_adj_1584));
    LocalMux I__7668 (
            .O(N__37477),
            .I(n14_adj_1584));
    InMux I__7667 (
            .O(N__37470),
            .I(n19638));
    InMux I__7666 (
            .O(N__37467),
            .I(N__37464));
    LocalMux I__7665 (
            .O(N__37464),
            .I(n22264));
    CascadeMux I__7664 (
            .O(N__37461),
            .I(n22414_cascade_));
    CascadeMux I__7663 (
            .O(N__37458),
            .I(n30_adj_1524_cascade_));
    CascadeMux I__7662 (
            .O(N__37455),
            .I(N__37452));
    InMux I__7661 (
            .O(N__37452),
            .I(N__37449));
    LocalMux I__7660 (
            .O(N__37449),
            .I(N__37444));
    InMux I__7659 (
            .O(N__37448),
            .I(N__37441));
    InMux I__7658 (
            .O(N__37447),
            .I(N__37437));
    Span4Mux_v I__7657 (
            .O(N__37444),
            .I(N__37432));
    LocalMux I__7656 (
            .O(N__37441),
            .I(N__37432));
    InMux I__7655 (
            .O(N__37440),
            .I(N__37428));
    LocalMux I__7654 (
            .O(N__37437),
            .I(N__37425));
    Span4Mux_v I__7653 (
            .O(N__37432),
            .I(N__37421));
    InMux I__7652 (
            .O(N__37431),
            .I(N__37418));
    LocalMux I__7651 (
            .O(N__37428),
            .I(N__37413));
    Span4Mux_v I__7650 (
            .O(N__37425),
            .I(N__37413));
    InMux I__7649 (
            .O(N__37424),
            .I(N__37410));
    Sp12to4 I__7648 (
            .O(N__37421),
            .I(N__37405));
    LocalMux I__7647 (
            .O(N__37418),
            .I(N__37405));
    Sp12to4 I__7646 (
            .O(N__37413),
            .I(N__37400));
    LocalMux I__7645 (
            .O(N__37410),
            .I(N__37400));
    Span12Mux_h I__7644 (
            .O(N__37405),
            .I(N__37397));
    Span12Mux_v I__7643 (
            .O(N__37400),
            .I(N__37394));
    Odrv12 I__7642 (
            .O(N__37397),
            .I(comm_buf_1_1));
    Odrv12 I__7641 (
            .O(N__37394),
            .I(comm_buf_1_1));
    InMux I__7640 (
            .O(N__37389),
            .I(N__37386));
    LocalMux I__7639 (
            .O(N__37386),
            .I(N__37382));
    InMux I__7638 (
            .O(N__37385),
            .I(N__37379));
    Span12Mux_v I__7637 (
            .O(N__37382),
            .I(N__37374));
    LocalMux I__7636 (
            .O(N__37379),
            .I(N__37374));
    Odrv12 I__7635 (
            .O(N__37374),
            .I(\comm_spi.n14623 ));
    SRMux I__7634 (
            .O(N__37371),
            .I(N__37368));
    LocalMux I__7633 (
            .O(N__37368),
            .I(N__37365));
    Span4Mux_h I__7632 (
            .O(N__37365),
            .I(N__37362));
    Odrv4 I__7631 (
            .O(N__37362),
            .I(\comm_spi.data_tx_7__N_770 ));
    InMux I__7630 (
            .O(N__37359),
            .I(N__37356));
    LocalMux I__7629 (
            .O(N__37356),
            .I(N__37352));
    InMux I__7628 (
            .O(N__37355),
            .I(N__37349));
    Odrv12 I__7627 (
            .O(N__37352),
            .I(\comm_spi.n14622 ));
    LocalMux I__7626 (
            .O(N__37349),
            .I(\comm_spi.n14622 ));
    InMux I__7625 (
            .O(N__37344),
            .I(N__37340));
    InMux I__7624 (
            .O(N__37343),
            .I(N__37337));
    LocalMux I__7623 (
            .O(N__37340),
            .I(N__37332));
    LocalMux I__7622 (
            .O(N__37337),
            .I(N__37332));
    Span4Mux_h I__7621 (
            .O(N__37332),
            .I(N__37329));
    Span4Mux_v I__7620 (
            .O(N__37329),
            .I(N__37325));
    InMux I__7619 (
            .O(N__37328),
            .I(N__37322));
    Odrv4 I__7618 (
            .O(N__37325),
            .I(\comm_spi.n22857 ));
    LocalMux I__7617 (
            .O(N__37322),
            .I(\comm_spi.n22857 ));
    InMux I__7616 (
            .O(N__37317),
            .I(N__37313));
    InMux I__7615 (
            .O(N__37316),
            .I(N__37310));
    LocalMux I__7614 (
            .O(N__37313),
            .I(N__37304));
    LocalMux I__7613 (
            .O(N__37310),
            .I(N__37301));
    CascadeMux I__7612 (
            .O(N__37309),
            .I(N__37294));
    InMux I__7611 (
            .O(N__37308),
            .I(N__37288));
    InMux I__7610 (
            .O(N__37307),
            .I(N__37285));
    Span4Mux_h I__7609 (
            .O(N__37304),
            .I(N__37282));
    Span4Mux_h I__7608 (
            .O(N__37301),
            .I(N__37279));
    CascadeMux I__7607 (
            .O(N__37300),
            .I(N__37276));
    CascadeMux I__7606 (
            .O(N__37299),
            .I(N__37273));
    CascadeMux I__7605 (
            .O(N__37298),
            .I(N__37269));
    InMux I__7604 (
            .O(N__37297),
            .I(N__37266));
    InMux I__7603 (
            .O(N__37294),
            .I(N__37263));
    InMux I__7602 (
            .O(N__37293),
            .I(N__37258));
    InMux I__7601 (
            .O(N__37292),
            .I(N__37258));
    InMux I__7600 (
            .O(N__37291),
            .I(N__37255));
    LocalMux I__7599 (
            .O(N__37288),
            .I(N__37250));
    LocalMux I__7598 (
            .O(N__37285),
            .I(N__37250));
    Span4Mux_v I__7597 (
            .O(N__37282),
            .I(N__37247));
    Span4Mux_v I__7596 (
            .O(N__37279),
            .I(N__37244));
    InMux I__7595 (
            .O(N__37276),
            .I(N__37235));
    InMux I__7594 (
            .O(N__37273),
            .I(N__37235));
    InMux I__7593 (
            .O(N__37272),
            .I(N__37235));
    InMux I__7592 (
            .O(N__37269),
            .I(N__37235));
    LocalMux I__7591 (
            .O(N__37266),
            .I(eis_state_1));
    LocalMux I__7590 (
            .O(N__37263),
            .I(eis_state_1));
    LocalMux I__7589 (
            .O(N__37258),
            .I(eis_state_1));
    LocalMux I__7588 (
            .O(N__37255),
            .I(eis_state_1));
    Odrv4 I__7587 (
            .O(N__37250),
            .I(eis_state_1));
    Odrv4 I__7586 (
            .O(N__37247),
            .I(eis_state_1));
    Odrv4 I__7585 (
            .O(N__37244),
            .I(eis_state_1));
    LocalMux I__7584 (
            .O(N__37235),
            .I(eis_state_1));
    CascadeMux I__7583 (
            .O(N__37218),
            .I(n20937_cascade_));
    InMux I__7582 (
            .O(N__37215),
            .I(N__37212));
    LocalMux I__7581 (
            .O(N__37212),
            .I(n20939));
    InMux I__7580 (
            .O(N__37209),
            .I(N__37206));
    LocalMux I__7579 (
            .O(N__37206),
            .I(n19_adj_1522));
    CascadeMux I__7578 (
            .O(N__37203),
            .I(N__37200));
    InMux I__7577 (
            .O(N__37200),
            .I(N__37197));
    LocalMux I__7576 (
            .O(N__37197),
            .I(N__37194));
    Span4Mux_h I__7575 (
            .O(N__37194),
            .I(N__37190));
    CascadeMux I__7574 (
            .O(N__37193),
            .I(N__37187));
    Span4Mux_h I__7573 (
            .O(N__37190),
            .I(N__37184));
    InMux I__7572 (
            .O(N__37187),
            .I(N__37181));
    Odrv4 I__7571 (
            .O(N__37184),
            .I(buf_readRTD_1));
    LocalMux I__7570 (
            .O(N__37181),
            .I(buf_readRTD_1));
    InMux I__7569 (
            .O(N__37176),
            .I(N__37173));
    LocalMux I__7568 (
            .O(N__37173),
            .I(N__37169));
    InMux I__7567 (
            .O(N__37172),
            .I(N__37166));
    Span4Mux_v I__7566 (
            .O(N__37169),
            .I(N__37163));
    LocalMux I__7565 (
            .O(N__37166),
            .I(N__37160));
    Span4Mux_h I__7564 (
            .O(N__37163),
            .I(N__37156));
    Sp12to4 I__7563 (
            .O(N__37160),
            .I(N__37153));
    InMux I__7562 (
            .O(N__37159),
            .I(N__37150));
    Sp12to4 I__7561 (
            .O(N__37156),
            .I(N__37145));
    Span12Mux_v I__7560 (
            .O(N__37153),
            .I(N__37145));
    LocalMux I__7559 (
            .O(N__37150),
            .I(buf_adcdata_iac_9));
    Odrv12 I__7558 (
            .O(N__37145),
            .I(buf_adcdata_iac_9));
    CascadeMux I__7557 (
            .O(N__37140),
            .I(n22261_cascade_));
    InMux I__7556 (
            .O(N__37137),
            .I(N__37134));
    LocalMux I__7555 (
            .O(N__37134),
            .I(N__37131));
    Span4Mux_v I__7554 (
            .O(N__37131),
            .I(N__37128));
    Odrv4 I__7553 (
            .O(N__37128),
            .I(n16_adj_1521));
    CascadeMux I__7552 (
            .O(N__37125),
            .I(n26_adj_1523_cascade_));
    InMux I__7551 (
            .O(N__37122),
            .I(N__37119));
    LocalMux I__7550 (
            .O(N__37119),
            .I(N__37116));
    Span4Mux_v I__7549 (
            .O(N__37116),
            .I(N__37112));
    InMux I__7548 (
            .O(N__37115),
            .I(N__37108));
    Span4Mux_h I__7547 (
            .O(N__37112),
            .I(N__37105));
    InMux I__7546 (
            .O(N__37111),
            .I(N__37102));
    LocalMux I__7545 (
            .O(N__37108),
            .I(acadc_skipCount_1));
    Odrv4 I__7544 (
            .O(N__37105),
            .I(acadc_skipCount_1));
    LocalMux I__7543 (
            .O(N__37102),
            .I(acadc_skipCount_1));
    CascadeMux I__7542 (
            .O(N__37095),
            .I(n22411_cascade_));
    InMux I__7541 (
            .O(N__37092),
            .I(N__37089));
    LocalMux I__7540 (
            .O(N__37089),
            .I(N__37086));
    Span4Mux_v I__7539 (
            .O(N__37086),
            .I(N__37082));
    InMux I__7538 (
            .O(N__37085),
            .I(N__37078));
    Span4Mux_v I__7537 (
            .O(N__37082),
            .I(N__37075));
    InMux I__7536 (
            .O(N__37081),
            .I(N__37072));
    LocalMux I__7535 (
            .O(N__37078),
            .I(req_data_cnt_1));
    Odrv4 I__7534 (
            .O(N__37075),
            .I(req_data_cnt_1));
    LocalMux I__7533 (
            .O(N__37072),
            .I(req_data_cnt_1));
    CascadeMux I__7532 (
            .O(N__37065),
            .I(n21370_cascade_));
    InMux I__7531 (
            .O(N__37062),
            .I(N__37059));
    LocalMux I__7530 (
            .O(N__37059),
            .I(n21369));
    InMux I__7529 (
            .O(N__37056),
            .I(N__37053));
    LocalMux I__7528 (
            .O(N__37053),
            .I(n22426));
    CEMux I__7527 (
            .O(N__37050),
            .I(N__37047));
    LocalMux I__7526 (
            .O(N__37047),
            .I(N__37044));
    Sp12to4 I__7525 (
            .O(N__37044),
            .I(N__37041));
    Odrv12 I__7524 (
            .O(N__37041),
            .I(n14));
    CascadeMux I__7523 (
            .O(N__37038),
            .I(n1264_cascade_));
    InMux I__7522 (
            .O(N__37035),
            .I(N__37032));
    LocalMux I__7521 (
            .O(N__37032),
            .I(n4_adj_1643));
    InMux I__7520 (
            .O(N__37029),
            .I(N__37025));
    InMux I__7519 (
            .O(N__37028),
            .I(N__37022));
    LocalMux I__7518 (
            .O(N__37025),
            .I(n1264));
    LocalMux I__7517 (
            .O(N__37022),
            .I(n1264));
    InMux I__7516 (
            .O(N__37017),
            .I(N__37014));
    LocalMux I__7515 (
            .O(N__37014),
            .I(n8_adj_1582));
    CascadeMux I__7514 (
            .O(N__37011),
            .I(N__37008));
    InMux I__7513 (
            .O(N__37008),
            .I(N__37005));
    LocalMux I__7512 (
            .O(N__37005),
            .I(comm_state_3_N_420_3));
    CascadeMux I__7511 (
            .O(N__37002),
            .I(comm_state_3_N_420_3_cascade_));
    CascadeMux I__7510 (
            .O(N__36999),
            .I(n21435_cascade_));
    CEMux I__7509 (
            .O(N__36996),
            .I(N__36993));
    LocalMux I__7508 (
            .O(N__36993),
            .I(N__36990));
    Span4Mux_h I__7507 (
            .O(N__36990),
            .I(N__36987));
    Odrv4 I__7506 (
            .O(N__36987),
            .I(n20829));
    CascadeMux I__7505 (
            .O(N__36984),
            .I(n20944_cascade_));
    CEMux I__7504 (
            .O(N__36981),
            .I(N__36978));
    LocalMux I__7503 (
            .O(N__36978),
            .I(n20964));
    InMux I__7502 (
            .O(N__36975),
            .I(N__36972));
    LocalMux I__7501 (
            .O(N__36972),
            .I(n20962));
    InMux I__7500 (
            .O(N__36969),
            .I(N__36963));
    InMux I__7499 (
            .O(N__36968),
            .I(N__36963));
    LocalMux I__7498 (
            .O(N__36963),
            .I(N__36960));
    Span12Mux_v I__7497 (
            .O(N__36960),
            .I(N__36957));
    Odrv12 I__7496 (
            .O(N__36957),
            .I(n3));
    InMux I__7495 (
            .O(N__36954),
            .I(N__36951));
    LocalMux I__7494 (
            .O(N__36951),
            .I(n20801));
    InMux I__7493 (
            .O(N__36948),
            .I(N__36945));
    LocalMux I__7492 (
            .O(N__36945),
            .I(n4_adj_1586));
    CascadeMux I__7491 (
            .O(N__36942),
            .I(n20801_cascade_));
    InMux I__7490 (
            .O(N__36939),
            .I(N__36936));
    LocalMux I__7489 (
            .O(N__36936),
            .I(n19902));
    InMux I__7488 (
            .O(N__36933),
            .I(N__36930));
    LocalMux I__7487 (
            .O(N__36930),
            .I(N__36927));
    Odrv4 I__7486 (
            .O(N__36927),
            .I(n22423));
    CascadeMux I__7485 (
            .O(N__36924),
            .I(n2_adj_1581_cascade_));
    InMux I__7484 (
            .O(N__36921),
            .I(N__36914));
    InMux I__7483 (
            .O(N__36920),
            .I(N__36914));
    InMux I__7482 (
            .O(N__36919),
            .I(N__36909));
    LocalMux I__7481 (
            .O(N__36914),
            .I(N__36906));
    InMux I__7480 (
            .O(N__36913),
            .I(N__36903));
    InMux I__7479 (
            .O(N__36912),
            .I(N__36900));
    LocalMux I__7478 (
            .O(N__36909),
            .I(N__36897));
    Span4Mux_h I__7477 (
            .O(N__36906),
            .I(N__36894));
    LocalMux I__7476 (
            .O(N__36903),
            .I(\ADC_VDC.bit_cnt_4 ));
    LocalMux I__7475 (
            .O(N__36900),
            .I(\ADC_VDC.bit_cnt_4 ));
    Odrv4 I__7474 (
            .O(N__36897),
            .I(\ADC_VDC.bit_cnt_4 ));
    Odrv4 I__7473 (
            .O(N__36894),
            .I(\ADC_VDC.bit_cnt_4 ));
    InMux I__7472 (
            .O(N__36885),
            .I(\ADC_VDC.n19775 ));
    CascadeMux I__7471 (
            .O(N__36882),
            .I(N__36876));
    InMux I__7470 (
            .O(N__36881),
            .I(N__36873));
    InMux I__7469 (
            .O(N__36880),
            .I(N__36868));
    InMux I__7468 (
            .O(N__36879),
            .I(N__36868));
    InMux I__7467 (
            .O(N__36876),
            .I(N__36865));
    LocalMux I__7466 (
            .O(N__36873),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__7465 (
            .O(N__36868),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__7464 (
            .O(N__36865),
            .I(\ADC_VDC.bit_cnt_5 ));
    InMux I__7463 (
            .O(N__36858),
            .I(\ADC_VDC.n19776 ));
    InMux I__7462 (
            .O(N__36855),
            .I(N__36849));
    InMux I__7461 (
            .O(N__36854),
            .I(N__36844));
    InMux I__7460 (
            .O(N__36853),
            .I(N__36844));
    InMux I__7459 (
            .O(N__36852),
            .I(N__36841));
    LocalMux I__7458 (
            .O(N__36849),
            .I(\ADC_VDC.bit_cnt_6 ));
    LocalMux I__7457 (
            .O(N__36844),
            .I(\ADC_VDC.bit_cnt_6 ));
    LocalMux I__7456 (
            .O(N__36841),
            .I(\ADC_VDC.bit_cnt_6 ));
    InMux I__7455 (
            .O(N__36834),
            .I(\ADC_VDC.n19777 ));
    InMux I__7454 (
            .O(N__36831),
            .I(\ADC_VDC.n19778 ));
    InMux I__7453 (
            .O(N__36828),
            .I(N__36822));
    InMux I__7452 (
            .O(N__36827),
            .I(N__36819));
    InMux I__7451 (
            .O(N__36826),
            .I(N__36816));
    InMux I__7450 (
            .O(N__36825),
            .I(N__36813));
    LocalMux I__7449 (
            .O(N__36822),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__7448 (
            .O(N__36819),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__7447 (
            .O(N__36816),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__7446 (
            .O(N__36813),
            .I(\ADC_VDC.bit_cnt_7 ));
    SRMux I__7445 (
            .O(N__36804),
            .I(N__36801));
    LocalMux I__7444 (
            .O(N__36801),
            .I(N__36798));
    Odrv4 I__7443 (
            .O(N__36798),
            .I(\ADC_VDC.n18550 ));
    SRMux I__7442 (
            .O(N__36795),
            .I(N__36792));
    LocalMux I__7441 (
            .O(N__36792),
            .I(N__36789));
    Span4Mux_h I__7440 (
            .O(N__36789),
            .I(N__36786));
    Span4Mux_v I__7439 (
            .O(N__36786),
            .I(N__36783));
    Odrv4 I__7438 (
            .O(N__36783),
            .I(\comm_spi.data_tx_7__N_786 ));
    InMux I__7437 (
            .O(N__36780),
            .I(N__36777));
    LocalMux I__7436 (
            .O(N__36777),
            .I(N__36774));
    Span4Mux_v I__7435 (
            .O(N__36774),
            .I(N__36770));
    InMux I__7434 (
            .O(N__36773),
            .I(N__36767));
    Odrv4 I__7433 (
            .O(N__36770),
            .I(tmp_buf_15));
    LocalMux I__7432 (
            .O(N__36767),
            .I(tmp_buf_15));
    IoInMux I__7431 (
            .O(N__36762),
            .I(N__36759));
    LocalMux I__7430 (
            .O(N__36759),
            .I(N__36756));
    Span12Mux_s1_v I__7429 (
            .O(N__36756),
            .I(N__36753));
    Span12Mux_h I__7428 (
            .O(N__36753),
            .I(N__36749));
    InMux I__7427 (
            .O(N__36752),
            .I(N__36746));
    Odrv12 I__7426 (
            .O(N__36749),
            .I(DDS_MOSI));
    LocalMux I__7425 (
            .O(N__36746),
            .I(DDS_MOSI));
    IoInMux I__7424 (
            .O(N__36741),
            .I(N__36738));
    LocalMux I__7423 (
            .O(N__36738),
            .I(N__36735));
    Span4Mux_s2_v I__7422 (
            .O(N__36735),
            .I(N__36732));
    Span4Mux_h I__7421 (
            .O(N__36732),
            .I(N__36729));
    Span4Mux_v I__7420 (
            .O(N__36729),
            .I(N__36726));
    Sp12to4 I__7419 (
            .O(N__36726),
            .I(N__36723));
    Odrv12 I__7418 (
            .O(N__36723),
            .I(DDS_CS));
    CEMux I__7417 (
            .O(N__36720),
            .I(N__36717));
    LocalMux I__7416 (
            .O(N__36717),
            .I(\SIG_DDS.n9_adj_1393 ));
    SRMux I__7415 (
            .O(N__36714),
            .I(N__36711));
    LocalMux I__7414 (
            .O(N__36711),
            .I(\comm_spi.data_tx_7__N_795 ));
    InMux I__7413 (
            .O(N__36708),
            .I(N__36701));
    CascadeMux I__7412 (
            .O(N__36707),
            .I(N__36698));
    CascadeMux I__7411 (
            .O(N__36706),
            .I(N__36695));
    InMux I__7410 (
            .O(N__36705),
            .I(N__36692));
    InMux I__7409 (
            .O(N__36704),
            .I(N__36689));
    LocalMux I__7408 (
            .O(N__36701),
            .I(N__36686));
    InMux I__7407 (
            .O(N__36698),
            .I(N__36681));
    InMux I__7406 (
            .O(N__36695),
            .I(N__36681));
    LocalMux I__7405 (
            .O(N__36692),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__7404 (
            .O(N__36689),
            .I(\ADC_VDC.bit_cnt_0 ));
    Odrv4 I__7403 (
            .O(N__36686),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__7402 (
            .O(N__36681),
            .I(\ADC_VDC.bit_cnt_0 ));
    InMux I__7401 (
            .O(N__36672),
            .I(bfn_15_4_0_));
    InMux I__7400 (
            .O(N__36669),
            .I(N__36663));
    InMux I__7399 (
            .O(N__36668),
            .I(N__36658));
    InMux I__7398 (
            .O(N__36667),
            .I(N__36658));
    InMux I__7397 (
            .O(N__36666),
            .I(N__36655));
    LocalMux I__7396 (
            .O(N__36663),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__7395 (
            .O(N__36658),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__7394 (
            .O(N__36655),
            .I(\ADC_VDC.bit_cnt_1 ));
    InMux I__7393 (
            .O(N__36648),
            .I(\ADC_VDC.n19772 ));
    InMux I__7392 (
            .O(N__36645),
            .I(N__36641));
    InMux I__7391 (
            .O(N__36644),
            .I(N__36635));
    LocalMux I__7390 (
            .O(N__36641),
            .I(N__36632));
    InMux I__7389 (
            .O(N__36640),
            .I(N__36629));
    InMux I__7388 (
            .O(N__36639),
            .I(N__36624));
    InMux I__7387 (
            .O(N__36638),
            .I(N__36624));
    LocalMux I__7386 (
            .O(N__36635),
            .I(\ADC_VDC.bit_cnt_2 ));
    Odrv4 I__7385 (
            .O(N__36632),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__7384 (
            .O(N__36629),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__7383 (
            .O(N__36624),
            .I(\ADC_VDC.bit_cnt_2 ));
    InMux I__7382 (
            .O(N__36615),
            .I(\ADC_VDC.n19773 ));
    InMux I__7381 (
            .O(N__36612),
            .I(N__36605));
    InMux I__7380 (
            .O(N__36611),
            .I(N__36605));
    InMux I__7379 (
            .O(N__36610),
            .I(N__36600));
    LocalMux I__7378 (
            .O(N__36605),
            .I(N__36597));
    InMux I__7377 (
            .O(N__36604),
            .I(N__36594));
    InMux I__7376 (
            .O(N__36603),
            .I(N__36591));
    LocalMux I__7375 (
            .O(N__36600),
            .I(\ADC_VDC.bit_cnt_3 ));
    Odrv4 I__7374 (
            .O(N__36597),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__7373 (
            .O(N__36594),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__7372 (
            .O(N__36591),
            .I(\ADC_VDC.bit_cnt_3 ));
    InMux I__7371 (
            .O(N__36582),
            .I(\ADC_VDC.n19774 ));
    InMux I__7370 (
            .O(N__36579),
            .I(n19629));
    InMux I__7369 (
            .O(N__36576),
            .I(n19630));
    InMux I__7368 (
            .O(N__36573),
            .I(n19631));
    InMux I__7367 (
            .O(N__36570),
            .I(bfn_14_19_0_));
    CascadeMux I__7366 (
            .O(N__36567),
            .I(N__36563));
    CascadeMux I__7365 (
            .O(N__36566),
            .I(N__36555));
    InMux I__7364 (
            .O(N__36563),
            .I(N__36552));
    CascadeMux I__7363 (
            .O(N__36562),
            .I(N__36549));
    CascadeMux I__7362 (
            .O(N__36561),
            .I(N__36546));
    CascadeMux I__7361 (
            .O(N__36560),
            .I(N__36543));
    CascadeMux I__7360 (
            .O(N__36559),
            .I(N__36540));
    CascadeMux I__7359 (
            .O(N__36558),
            .I(N__36533));
    InMux I__7358 (
            .O(N__36555),
            .I(N__36530));
    LocalMux I__7357 (
            .O(N__36552),
            .I(N__36527));
    InMux I__7356 (
            .O(N__36549),
            .I(N__36518));
    InMux I__7355 (
            .O(N__36546),
            .I(N__36518));
    InMux I__7354 (
            .O(N__36543),
            .I(N__36518));
    InMux I__7353 (
            .O(N__36540),
            .I(N__36518));
    CascadeMux I__7352 (
            .O(N__36539),
            .I(N__36515));
    CascadeMux I__7351 (
            .O(N__36538),
            .I(N__36512));
    CascadeMux I__7350 (
            .O(N__36537),
            .I(N__36509));
    CascadeMux I__7349 (
            .O(N__36536),
            .I(N__36506));
    InMux I__7348 (
            .O(N__36533),
            .I(N__36503));
    LocalMux I__7347 (
            .O(N__36530),
            .I(N__36496));
    Span4Mux_h I__7346 (
            .O(N__36527),
            .I(N__36496));
    LocalMux I__7345 (
            .O(N__36518),
            .I(N__36496));
    InMux I__7344 (
            .O(N__36515),
            .I(N__36487));
    InMux I__7343 (
            .O(N__36512),
            .I(N__36487));
    InMux I__7342 (
            .O(N__36509),
            .I(N__36487));
    InMux I__7341 (
            .O(N__36506),
            .I(N__36487));
    LocalMux I__7340 (
            .O(N__36503),
            .I(n10598));
    Odrv4 I__7339 (
            .O(N__36496),
            .I(n10598));
    LocalMux I__7338 (
            .O(N__36487),
            .I(n10598));
    InMux I__7337 (
            .O(N__36480),
            .I(n19633));
    InMux I__7336 (
            .O(N__36477),
            .I(N__36473));
    InMux I__7335 (
            .O(N__36476),
            .I(N__36470));
    LocalMux I__7334 (
            .O(N__36473),
            .I(n7_adj_1572));
    LocalMux I__7333 (
            .O(N__36470),
            .I(n7_adj_1572));
    InMux I__7332 (
            .O(N__36465),
            .I(N__36462));
    LocalMux I__7331 (
            .O(N__36462),
            .I(n8_adj_1573));
    CascadeMux I__7330 (
            .O(N__36459),
            .I(N__36456));
    CascadeBuf I__7329 (
            .O(N__36456),
            .I(N__36453));
    CascadeMux I__7328 (
            .O(N__36453),
            .I(N__36450));
    CascadeBuf I__7327 (
            .O(N__36450),
            .I(N__36447));
    CascadeMux I__7326 (
            .O(N__36447),
            .I(N__36444));
    CascadeBuf I__7325 (
            .O(N__36444),
            .I(N__36441));
    CascadeMux I__7324 (
            .O(N__36441),
            .I(N__36438));
    CascadeBuf I__7323 (
            .O(N__36438),
            .I(N__36435));
    CascadeMux I__7322 (
            .O(N__36435),
            .I(N__36432));
    CascadeBuf I__7321 (
            .O(N__36432),
            .I(N__36429));
    CascadeMux I__7320 (
            .O(N__36429),
            .I(N__36426));
    CascadeBuf I__7319 (
            .O(N__36426),
            .I(N__36423));
    CascadeMux I__7318 (
            .O(N__36423),
            .I(N__36420));
    CascadeBuf I__7317 (
            .O(N__36420),
            .I(N__36417));
    CascadeMux I__7316 (
            .O(N__36417),
            .I(N__36413));
    CascadeMux I__7315 (
            .O(N__36416),
            .I(N__36410));
    CascadeBuf I__7314 (
            .O(N__36413),
            .I(N__36407));
    CascadeBuf I__7313 (
            .O(N__36410),
            .I(N__36404));
    CascadeMux I__7312 (
            .O(N__36407),
            .I(N__36401));
    CascadeMux I__7311 (
            .O(N__36404),
            .I(N__36398));
    CascadeBuf I__7310 (
            .O(N__36401),
            .I(N__36395));
    InMux I__7309 (
            .O(N__36398),
            .I(N__36392));
    CascadeMux I__7308 (
            .O(N__36395),
            .I(N__36389));
    LocalMux I__7307 (
            .O(N__36392),
            .I(N__36386));
    InMux I__7306 (
            .O(N__36389),
            .I(N__36383));
    Span12Mux_h I__7305 (
            .O(N__36386),
            .I(N__36380));
    LocalMux I__7304 (
            .O(N__36383),
            .I(N__36377));
    Span12Mux_v I__7303 (
            .O(N__36380),
            .I(N__36374));
    Span4Mux_h I__7302 (
            .O(N__36377),
            .I(N__36371));
    Odrv12 I__7301 (
            .O(N__36374),
            .I(data_index_9_N_216_1));
    Odrv4 I__7300 (
            .O(N__36371),
            .I(data_index_9_N_216_1));
    CascadeMux I__7299 (
            .O(N__36366),
            .I(N__36362));
    IoInMux I__7298 (
            .O(N__36365),
            .I(N__36359));
    InMux I__7297 (
            .O(N__36362),
            .I(N__36356));
    LocalMux I__7296 (
            .O(N__36359),
            .I(N__36353));
    LocalMux I__7295 (
            .O(N__36356),
            .I(N__36349));
    Span12Mux_s7_v I__7294 (
            .O(N__36353),
            .I(N__36346));
    InMux I__7293 (
            .O(N__36352),
            .I(N__36343));
    Span4Mux_h I__7292 (
            .O(N__36349),
            .I(N__36340));
    Odrv12 I__7291 (
            .O(N__36346),
            .I(DDS_RNG_0));
    LocalMux I__7290 (
            .O(N__36343),
            .I(DDS_RNG_0));
    Odrv4 I__7289 (
            .O(N__36340),
            .I(DDS_RNG_0));
    InMux I__7288 (
            .O(N__36333),
            .I(N__36330));
    LocalMux I__7287 (
            .O(N__36330),
            .I(n11338));
    CascadeMux I__7286 (
            .O(N__36327),
            .I(n11338_cascade_));
    CascadeMux I__7285 (
            .O(N__36324),
            .I(n8813_cascade_));
    InMux I__7284 (
            .O(N__36321),
            .I(N__36316));
    InMux I__7283 (
            .O(N__36320),
            .I(N__36313));
    InMux I__7282 (
            .O(N__36319),
            .I(N__36310));
    LocalMux I__7281 (
            .O(N__36316),
            .I(data_index_0));
    LocalMux I__7280 (
            .O(N__36313),
            .I(data_index_0));
    LocalMux I__7279 (
            .O(N__36310),
            .I(data_index_0));
    InMux I__7278 (
            .O(N__36303),
            .I(N__36297));
    InMux I__7277 (
            .O(N__36302),
            .I(N__36297));
    LocalMux I__7276 (
            .O(N__36297),
            .I(N__36294));
    Odrv12 I__7275 (
            .O(N__36294),
            .I(n7));
    InMux I__7274 (
            .O(N__36291),
            .I(bfn_14_18_0_));
    InMux I__7273 (
            .O(N__36288),
            .I(N__36283));
    InMux I__7272 (
            .O(N__36287),
            .I(N__36280));
    InMux I__7271 (
            .O(N__36286),
            .I(N__36277));
    LocalMux I__7270 (
            .O(N__36283),
            .I(data_index_1));
    LocalMux I__7269 (
            .O(N__36280),
            .I(data_index_1));
    LocalMux I__7268 (
            .O(N__36277),
            .I(data_index_1));
    InMux I__7267 (
            .O(N__36270),
            .I(n19625));
    InMux I__7266 (
            .O(N__36267),
            .I(n19626));
    InMux I__7265 (
            .O(N__36264),
            .I(n19627));
    InMux I__7264 (
            .O(N__36261),
            .I(n19628));
    InMux I__7263 (
            .O(N__36258),
            .I(N__36255));
    LocalMux I__7262 (
            .O(N__36255),
            .I(N__36251));
    InMux I__7261 (
            .O(N__36254),
            .I(N__36248));
    Span4Mux_v I__7260 (
            .O(N__36251),
            .I(N__36244));
    LocalMux I__7259 (
            .O(N__36248),
            .I(N__36241));
    InMux I__7258 (
            .O(N__36247),
            .I(N__36238));
    Odrv4 I__7257 (
            .O(N__36244),
            .I(n10520));
    Odrv12 I__7256 (
            .O(N__36241),
            .I(n10520));
    LocalMux I__7255 (
            .O(N__36238),
            .I(n10520));
    InMux I__7254 (
            .O(N__36231),
            .I(N__36227));
    CascadeMux I__7253 (
            .O(N__36230),
            .I(N__36224));
    LocalMux I__7252 (
            .O(N__36227),
            .I(N__36220));
    InMux I__7251 (
            .O(N__36224),
            .I(N__36217));
    InMux I__7250 (
            .O(N__36223),
            .I(N__36214));
    Span4Mux_h I__7249 (
            .O(N__36220),
            .I(N__36209));
    LocalMux I__7248 (
            .O(N__36217),
            .I(N__36209));
    LocalMux I__7247 (
            .O(N__36214),
            .I(req_data_cnt_15));
    Odrv4 I__7246 (
            .O(N__36209),
            .I(req_data_cnt_15));
    CascadeMux I__7245 (
            .O(N__36204),
            .I(n8_adj_1532_cascade_));
    CascadeMux I__7244 (
            .O(N__36201),
            .I(N__36198));
    CascadeBuf I__7243 (
            .O(N__36198),
            .I(N__36195));
    CascadeMux I__7242 (
            .O(N__36195),
            .I(N__36192));
    CascadeBuf I__7241 (
            .O(N__36192),
            .I(N__36189));
    CascadeMux I__7240 (
            .O(N__36189),
            .I(N__36186));
    CascadeBuf I__7239 (
            .O(N__36186),
            .I(N__36183));
    CascadeMux I__7238 (
            .O(N__36183),
            .I(N__36180));
    CascadeBuf I__7237 (
            .O(N__36180),
            .I(N__36177));
    CascadeMux I__7236 (
            .O(N__36177),
            .I(N__36174));
    CascadeBuf I__7235 (
            .O(N__36174),
            .I(N__36171));
    CascadeMux I__7234 (
            .O(N__36171),
            .I(N__36168));
    CascadeBuf I__7233 (
            .O(N__36168),
            .I(N__36165));
    CascadeMux I__7232 (
            .O(N__36165),
            .I(N__36162));
    CascadeBuf I__7231 (
            .O(N__36162),
            .I(N__36159));
    CascadeMux I__7230 (
            .O(N__36159),
            .I(N__36155));
    CascadeMux I__7229 (
            .O(N__36158),
            .I(N__36152));
    CascadeBuf I__7228 (
            .O(N__36155),
            .I(N__36149));
    CascadeBuf I__7227 (
            .O(N__36152),
            .I(N__36146));
    CascadeMux I__7226 (
            .O(N__36149),
            .I(N__36143));
    CascadeMux I__7225 (
            .O(N__36146),
            .I(N__36140));
    CascadeBuf I__7224 (
            .O(N__36143),
            .I(N__36137));
    InMux I__7223 (
            .O(N__36140),
            .I(N__36134));
    CascadeMux I__7222 (
            .O(N__36137),
            .I(N__36131));
    LocalMux I__7221 (
            .O(N__36134),
            .I(N__36128));
    InMux I__7220 (
            .O(N__36131),
            .I(N__36125));
    Span4Mux_h I__7219 (
            .O(N__36128),
            .I(N__36122));
    LocalMux I__7218 (
            .O(N__36125),
            .I(N__36119));
    Sp12to4 I__7217 (
            .O(N__36122),
            .I(N__36116));
    Span4Mux_v I__7216 (
            .O(N__36119),
            .I(N__36113));
    Span12Mux_v I__7215 (
            .O(N__36116),
            .I(N__36110));
    Span4Mux_h I__7214 (
            .O(N__36113),
            .I(N__36107));
    Odrv12 I__7213 (
            .O(N__36110),
            .I(data_index_9_N_216_0));
    Odrv4 I__7212 (
            .O(N__36107),
            .I(data_index_9_N_216_0));
    InMux I__7211 (
            .O(N__36102),
            .I(N__36099));
    LocalMux I__7210 (
            .O(N__36099),
            .I(n8_adj_1532));
    CEMux I__7209 (
            .O(N__36096),
            .I(N__36093));
    LocalMux I__7208 (
            .O(N__36093),
            .I(N__36089));
    CEMux I__7207 (
            .O(N__36092),
            .I(N__36086));
    Span4Mux_v I__7206 (
            .O(N__36089),
            .I(N__36083));
    LocalMux I__7205 (
            .O(N__36086),
            .I(N__36080));
    Span4Mux_h I__7204 (
            .O(N__36083),
            .I(N__36075));
    Span4Mux_h I__7203 (
            .O(N__36080),
            .I(N__36075));
    Odrv4 I__7202 (
            .O(N__36075),
            .I(\SIG_DDS.n9 ));
    InMux I__7201 (
            .O(N__36072),
            .I(N__36069));
    LocalMux I__7200 (
            .O(N__36069),
            .I(n22_adj_1499));
    InMux I__7199 (
            .O(N__36066),
            .I(N__36063));
    LocalMux I__7198 (
            .O(N__36063),
            .I(n18));
    CascadeMux I__7197 (
            .O(N__36060),
            .I(N__36057));
    InMux I__7196 (
            .O(N__36057),
            .I(N__36052));
    InMux I__7195 (
            .O(N__36056),
            .I(N__36047));
    InMux I__7194 (
            .O(N__36055),
            .I(N__36047));
    LocalMux I__7193 (
            .O(N__36052),
            .I(N__36044));
    LocalMux I__7192 (
            .O(N__36047),
            .I(req_data_cnt_14));
    Odrv4 I__7191 (
            .O(N__36044),
            .I(req_data_cnt_14));
    InMux I__7190 (
            .O(N__36039),
            .I(N__36036));
    LocalMux I__7189 (
            .O(N__36036),
            .I(n23_adj_1614));
    CascadeMux I__7188 (
            .O(N__36033),
            .I(n10_adj_1554_cascade_));
    CEMux I__7187 (
            .O(N__36030),
            .I(N__36027));
    LocalMux I__7186 (
            .O(N__36027),
            .I(N__36024));
    Span4Mux_v I__7185 (
            .O(N__36024),
            .I(N__36021));
    Odrv4 I__7184 (
            .O(N__36021),
            .I(n11850));
    CascadeMux I__7183 (
            .O(N__36018),
            .I(n20914_cascade_));
    InMux I__7182 (
            .O(N__36015),
            .I(N__36012));
    LocalMux I__7181 (
            .O(N__36012),
            .I(n21014));
    CascadeMux I__7180 (
            .O(N__36009),
            .I(N__36006));
    InMux I__7179 (
            .O(N__36006),
            .I(N__36003));
    LocalMux I__7178 (
            .O(N__36003),
            .I(n17_adj_1489));
    CascadeMux I__7177 (
            .O(N__36000),
            .I(n16891_cascade_));
    InMux I__7176 (
            .O(N__35997),
            .I(N__35994));
    LocalMux I__7175 (
            .O(N__35994),
            .I(N__35991));
    Span4Mux_v I__7174 (
            .O(N__35991),
            .I(N__35988));
    Span4Mux_h I__7173 (
            .O(N__35988),
            .I(N__35985));
    Odrv4 I__7172 (
            .O(N__35985),
            .I(\SIG_DDS.n21571 ));
    InMux I__7171 (
            .O(N__35982),
            .I(N__35979));
    LocalMux I__7170 (
            .O(N__35979),
            .I(N__35976));
    Span4Mux_v I__7169 (
            .O(N__35976),
            .I(N__35973));
    Span4Mux_v I__7168 (
            .O(N__35973),
            .I(N__35969));
    InMux I__7167 (
            .O(N__35972),
            .I(N__35966));
    Odrv4 I__7166 (
            .O(N__35969),
            .I(buf_adcdata_vdc_10));
    LocalMux I__7165 (
            .O(N__35966),
            .I(buf_adcdata_vdc_10));
    InMux I__7164 (
            .O(N__35961),
            .I(N__35958));
    LocalMux I__7163 (
            .O(N__35958),
            .I(N__35955));
    Span4Mux_v I__7162 (
            .O(N__35955),
            .I(N__35951));
    CascadeMux I__7161 (
            .O(N__35954),
            .I(N__35948));
    Span4Mux_h I__7160 (
            .O(N__35951),
            .I(N__35944));
    InMux I__7159 (
            .O(N__35948),
            .I(N__35941));
    InMux I__7158 (
            .O(N__35947),
            .I(N__35938));
    Span4Mux_h I__7157 (
            .O(N__35944),
            .I(N__35935));
    LocalMux I__7156 (
            .O(N__35941),
            .I(buf_adcdata_vac_10));
    LocalMux I__7155 (
            .O(N__35938),
            .I(buf_adcdata_vac_10));
    Odrv4 I__7154 (
            .O(N__35935),
            .I(buf_adcdata_vac_10));
    IoInMux I__7153 (
            .O(N__35928),
            .I(N__35925));
    LocalMux I__7152 (
            .O(N__35925),
            .I(N__35922));
    Span4Mux_s2_h I__7151 (
            .O(N__35922),
            .I(N__35919));
    Sp12to4 I__7150 (
            .O(N__35919),
            .I(N__35916));
    Span12Mux_v I__7149 (
            .O(N__35916),
            .I(N__35913));
    Span12Mux_h I__7148 (
            .O(N__35913),
            .I(N__35910));
    Odrv12 I__7147 (
            .O(N__35910),
            .I(ICE_GPMI_0));
    CEMux I__7146 (
            .O(N__35907),
            .I(N__35904));
    LocalMux I__7145 (
            .O(N__35904),
            .I(N__35901));
    Odrv4 I__7144 (
            .O(N__35901),
            .I(n11385));
    InMux I__7143 (
            .O(N__35898),
            .I(N__35895));
    LocalMux I__7142 (
            .O(N__35895),
            .I(N__35885));
    InMux I__7141 (
            .O(N__35894),
            .I(N__35869));
    InMux I__7140 (
            .O(N__35893),
            .I(N__35869));
    InMux I__7139 (
            .O(N__35892),
            .I(N__35869));
    InMux I__7138 (
            .O(N__35891),
            .I(N__35869));
    InMux I__7137 (
            .O(N__35890),
            .I(N__35869));
    InMux I__7136 (
            .O(N__35889),
            .I(N__35869));
    InMux I__7135 (
            .O(N__35888),
            .I(N__35869));
    Span4Mux_v I__7134 (
            .O(N__35885),
            .I(N__35866));
    InMux I__7133 (
            .O(N__35884),
            .I(N__35863));
    LocalMux I__7132 (
            .O(N__35869),
            .I(N__35860));
    Odrv4 I__7131 (
            .O(N__35866),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__7130 (
            .O(N__35863),
            .I(\comm_spi.bit_cnt_3 ));
    Odrv4 I__7129 (
            .O(N__35860),
            .I(\comm_spi.bit_cnt_3 ));
    InMux I__7128 (
            .O(N__35853),
            .I(N__35850));
    LocalMux I__7127 (
            .O(N__35850),
            .I(N__35847));
    Span4Mux_v I__7126 (
            .O(N__35847),
            .I(N__35837));
    InMux I__7125 (
            .O(N__35846),
            .I(N__35822));
    InMux I__7124 (
            .O(N__35845),
            .I(N__35822));
    InMux I__7123 (
            .O(N__35844),
            .I(N__35822));
    InMux I__7122 (
            .O(N__35843),
            .I(N__35822));
    InMux I__7121 (
            .O(N__35842),
            .I(N__35822));
    InMux I__7120 (
            .O(N__35841),
            .I(N__35822));
    InMux I__7119 (
            .O(N__35840),
            .I(N__35822));
    Odrv4 I__7118 (
            .O(N__35837),
            .I(\comm_spi.n17036 ));
    LocalMux I__7117 (
            .O(N__35822),
            .I(\comm_spi.n17036 ));
    CascadeMux I__7116 (
            .O(N__35817),
            .I(N__35812));
    CascadeMux I__7115 (
            .O(N__35816),
            .I(N__35809));
    InMux I__7114 (
            .O(N__35815),
            .I(N__35799));
    InMux I__7113 (
            .O(N__35812),
            .I(N__35792));
    InMux I__7112 (
            .O(N__35809),
            .I(N__35792));
    InMux I__7111 (
            .O(N__35808),
            .I(N__35789));
    InMux I__7110 (
            .O(N__35807),
            .I(N__35786));
    InMux I__7109 (
            .O(N__35806),
            .I(N__35783));
    InMux I__7108 (
            .O(N__35805),
            .I(N__35780));
    InMux I__7107 (
            .O(N__35804),
            .I(N__35771));
    InMux I__7106 (
            .O(N__35803),
            .I(N__35771));
    InMux I__7105 (
            .O(N__35802),
            .I(N__35768));
    LocalMux I__7104 (
            .O(N__35799),
            .I(N__35765));
    InMux I__7103 (
            .O(N__35798),
            .I(N__35760));
    InMux I__7102 (
            .O(N__35797),
            .I(N__35760));
    LocalMux I__7101 (
            .O(N__35792),
            .I(N__35751));
    LocalMux I__7100 (
            .O(N__35789),
            .I(N__35751));
    LocalMux I__7099 (
            .O(N__35786),
            .I(N__35748));
    LocalMux I__7098 (
            .O(N__35783),
            .I(N__35743));
    LocalMux I__7097 (
            .O(N__35780),
            .I(N__35743));
    InMux I__7096 (
            .O(N__35779),
            .I(N__35735));
    InMux I__7095 (
            .O(N__35778),
            .I(N__35735));
    InMux I__7094 (
            .O(N__35777),
            .I(N__35735));
    InMux I__7093 (
            .O(N__35776),
            .I(N__35732));
    LocalMux I__7092 (
            .O(N__35771),
            .I(N__35729));
    LocalMux I__7091 (
            .O(N__35768),
            .I(N__35726));
    Span4Mux_v I__7090 (
            .O(N__35765),
            .I(N__35723));
    LocalMux I__7089 (
            .O(N__35760),
            .I(N__35720));
    InMux I__7088 (
            .O(N__35759),
            .I(N__35712));
    InMux I__7087 (
            .O(N__35758),
            .I(N__35712));
    InMux I__7086 (
            .O(N__35757),
            .I(N__35712));
    InMux I__7085 (
            .O(N__35756),
            .I(N__35709));
    Span4Mux_v I__7084 (
            .O(N__35751),
            .I(N__35706));
    Span4Mux_v I__7083 (
            .O(N__35748),
            .I(N__35703));
    Span4Mux_h I__7082 (
            .O(N__35743),
            .I(N__35698));
    InMux I__7081 (
            .O(N__35742),
            .I(N__35695));
    LocalMux I__7080 (
            .O(N__35735),
            .I(N__35688));
    LocalMux I__7079 (
            .O(N__35732),
            .I(N__35688));
    Span4Mux_h I__7078 (
            .O(N__35729),
            .I(N__35688));
    Span4Mux_v I__7077 (
            .O(N__35726),
            .I(N__35681));
    Span4Mux_h I__7076 (
            .O(N__35723),
            .I(N__35681));
    Span4Mux_v I__7075 (
            .O(N__35720),
            .I(N__35681));
    InMux I__7074 (
            .O(N__35719),
            .I(N__35678));
    LocalMux I__7073 (
            .O(N__35712),
            .I(N__35675));
    LocalMux I__7072 (
            .O(N__35709),
            .I(N__35668));
    Span4Mux_v I__7071 (
            .O(N__35706),
            .I(N__35668));
    Span4Mux_h I__7070 (
            .O(N__35703),
            .I(N__35668));
    InMux I__7069 (
            .O(N__35702),
            .I(N__35663));
    InMux I__7068 (
            .O(N__35701),
            .I(N__35663));
    Span4Mux_h I__7067 (
            .O(N__35698),
            .I(N__35660));
    LocalMux I__7066 (
            .O(N__35695),
            .I(N__35653));
    Span4Mux_h I__7065 (
            .O(N__35688),
            .I(N__35653));
    Span4Mux_v I__7064 (
            .O(N__35681),
            .I(N__35653));
    LocalMux I__7063 (
            .O(N__35678),
            .I(N__35646));
    Span4Mux_h I__7062 (
            .O(N__35675),
            .I(N__35646));
    Span4Mux_h I__7061 (
            .O(N__35668),
            .I(N__35646));
    LocalMux I__7060 (
            .O(N__35663),
            .I(n20858));
    Odrv4 I__7059 (
            .O(N__35660),
            .I(n20858));
    Odrv4 I__7058 (
            .O(N__35653),
            .I(n20858));
    Odrv4 I__7057 (
            .O(N__35646),
            .I(n20858));
    InMux I__7056 (
            .O(N__35637),
            .I(N__35613));
    InMux I__7055 (
            .O(N__35636),
            .I(N__35608));
    InMux I__7054 (
            .O(N__35635),
            .I(N__35608));
    InMux I__7053 (
            .O(N__35634),
            .I(N__35599));
    InMux I__7052 (
            .O(N__35633),
            .I(N__35599));
    InMux I__7051 (
            .O(N__35632),
            .I(N__35599));
    InMux I__7050 (
            .O(N__35631),
            .I(N__35599));
    InMux I__7049 (
            .O(N__35630),
            .I(N__35595));
    InMux I__7048 (
            .O(N__35629),
            .I(N__35586));
    InMux I__7047 (
            .O(N__35628),
            .I(N__35586));
    InMux I__7046 (
            .O(N__35627),
            .I(N__35586));
    InMux I__7045 (
            .O(N__35626),
            .I(N__35586));
    InMux I__7044 (
            .O(N__35625),
            .I(N__35580));
    InMux I__7043 (
            .O(N__35624),
            .I(N__35580));
    InMux I__7042 (
            .O(N__35623),
            .I(N__35574));
    InMux I__7041 (
            .O(N__35622),
            .I(N__35574));
    CascadeMux I__7040 (
            .O(N__35621),
            .I(N__35571));
    InMux I__7039 (
            .O(N__35620),
            .I(N__35560));
    InMux I__7038 (
            .O(N__35619),
            .I(N__35560));
    InMux I__7037 (
            .O(N__35618),
            .I(N__35560));
    InMux I__7036 (
            .O(N__35617),
            .I(N__35560));
    InMux I__7035 (
            .O(N__35616),
            .I(N__35548));
    LocalMux I__7034 (
            .O(N__35613),
            .I(N__35545));
    LocalMux I__7033 (
            .O(N__35608),
            .I(N__35542));
    LocalMux I__7032 (
            .O(N__35599),
            .I(N__35539));
    CascadeMux I__7031 (
            .O(N__35598),
            .I(N__35532));
    LocalMux I__7030 (
            .O(N__35595),
            .I(N__35521));
    LocalMux I__7029 (
            .O(N__35586),
            .I(N__35521));
    CascadeMux I__7028 (
            .O(N__35585),
            .I(N__35517));
    LocalMux I__7027 (
            .O(N__35580),
            .I(N__35514));
    InMux I__7026 (
            .O(N__35579),
            .I(N__35511));
    LocalMux I__7025 (
            .O(N__35574),
            .I(N__35508));
    InMux I__7024 (
            .O(N__35571),
            .I(N__35503));
    InMux I__7023 (
            .O(N__35570),
            .I(N__35503));
    InMux I__7022 (
            .O(N__35569),
            .I(N__35500));
    LocalMux I__7021 (
            .O(N__35560),
            .I(N__35497));
    InMux I__7020 (
            .O(N__35559),
            .I(N__35487));
    InMux I__7019 (
            .O(N__35558),
            .I(N__35487));
    InMux I__7018 (
            .O(N__35557),
            .I(N__35478));
    InMux I__7017 (
            .O(N__35556),
            .I(N__35478));
    InMux I__7016 (
            .O(N__35555),
            .I(N__35478));
    InMux I__7015 (
            .O(N__35554),
            .I(N__35478));
    InMux I__7014 (
            .O(N__35553),
            .I(N__35473));
    InMux I__7013 (
            .O(N__35552),
            .I(N__35473));
    InMux I__7012 (
            .O(N__35551),
            .I(N__35470));
    LocalMux I__7011 (
            .O(N__35548),
            .I(N__35465));
    Span4Mux_h I__7010 (
            .O(N__35545),
            .I(N__35465));
    Span4Mux_h I__7009 (
            .O(N__35542),
            .I(N__35460));
    Span4Mux_h I__7008 (
            .O(N__35539),
            .I(N__35460));
    InMux I__7007 (
            .O(N__35538),
            .I(N__35449));
    InMux I__7006 (
            .O(N__35537),
            .I(N__35449));
    InMux I__7005 (
            .O(N__35536),
            .I(N__35449));
    InMux I__7004 (
            .O(N__35535),
            .I(N__35449));
    InMux I__7003 (
            .O(N__35532),
            .I(N__35446));
    InMux I__7002 (
            .O(N__35531),
            .I(N__35443));
    InMux I__7001 (
            .O(N__35530),
            .I(N__35432));
    InMux I__7000 (
            .O(N__35529),
            .I(N__35432));
    InMux I__6999 (
            .O(N__35528),
            .I(N__35432));
    InMux I__6998 (
            .O(N__35527),
            .I(N__35432));
    InMux I__6997 (
            .O(N__35526),
            .I(N__35432));
    Span4Mux_v I__6996 (
            .O(N__35521),
            .I(N__35429));
    InMux I__6995 (
            .O(N__35520),
            .I(N__35426));
    InMux I__6994 (
            .O(N__35517),
            .I(N__35423));
    Span4Mux_h I__6993 (
            .O(N__35514),
            .I(N__35420));
    LocalMux I__6992 (
            .O(N__35511),
            .I(N__35417));
    Span4Mux_v I__6991 (
            .O(N__35508),
            .I(N__35412));
    LocalMux I__6990 (
            .O(N__35503),
            .I(N__35412));
    LocalMux I__6989 (
            .O(N__35500),
            .I(N__35398));
    Span4Mux_h I__6988 (
            .O(N__35497),
            .I(N__35395));
    InMux I__6987 (
            .O(N__35496),
            .I(N__35383));
    InMux I__6986 (
            .O(N__35495),
            .I(N__35383));
    InMux I__6985 (
            .O(N__35494),
            .I(N__35383));
    InMux I__6984 (
            .O(N__35493),
            .I(N__35383));
    InMux I__6983 (
            .O(N__35492),
            .I(N__35383));
    LocalMux I__6982 (
            .O(N__35487),
            .I(N__35380));
    LocalMux I__6981 (
            .O(N__35478),
            .I(N__35369));
    LocalMux I__6980 (
            .O(N__35473),
            .I(N__35369));
    LocalMux I__6979 (
            .O(N__35470),
            .I(N__35369));
    Span4Mux_h I__6978 (
            .O(N__35465),
            .I(N__35369));
    Span4Mux_v I__6977 (
            .O(N__35460),
            .I(N__35369));
    InMux I__6976 (
            .O(N__35459),
            .I(N__35366));
    InMux I__6975 (
            .O(N__35458),
            .I(N__35363));
    LocalMux I__6974 (
            .O(N__35449),
            .I(N__35360));
    LocalMux I__6973 (
            .O(N__35446),
            .I(N__35353));
    LocalMux I__6972 (
            .O(N__35443),
            .I(N__35353));
    LocalMux I__6971 (
            .O(N__35432),
            .I(N__35353));
    Span4Mux_v I__6970 (
            .O(N__35429),
            .I(N__35350));
    LocalMux I__6969 (
            .O(N__35426),
            .I(N__35339));
    LocalMux I__6968 (
            .O(N__35423),
            .I(N__35339));
    Span4Mux_v I__6967 (
            .O(N__35420),
            .I(N__35339));
    Span4Mux_h I__6966 (
            .O(N__35417),
            .I(N__35339));
    Span4Mux_h I__6965 (
            .O(N__35412),
            .I(N__35339));
    InMux I__6964 (
            .O(N__35411),
            .I(N__35326));
    InMux I__6963 (
            .O(N__35410),
            .I(N__35326));
    InMux I__6962 (
            .O(N__35409),
            .I(N__35326));
    InMux I__6961 (
            .O(N__35408),
            .I(N__35326));
    InMux I__6960 (
            .O(N__35407),
            .I(N__35326));
    InMux I__6959 (
            .O(N__35406),
            .I(N__35326));
    InMux I__6958 (
            .O(N__35405),
            .I(N__35321));
    InMux I__6957 (
            .O(N__35404),
            .I(N__35318));
    InMux I__6956 (
            .O(N__35403),
            .I(N__35315));
    InMux I__6955 (
            .O(N__35402),
            .I(N__35312));
    InMux I__6954 (
            .O(N__35401),
            .I(N__35309));
    Span4Mux_h I__6953 (
            .O(N__35398),
            .I(N__35304));
    Span4Mux_v I__6952 (
            .O(N__35395),
            .I(N__35304));
    InMux I__6951 (
            .O(N__35394),
            .I(N__35301));
    LocalMux I__6950 (
            .O(N__35383),
            .I(N__35294));
    Span4Mux_h I__6949 (
            .O(N__35380),
            .I(N__35294));
    Span4Mux_v I__6948 (
            .O(N__35369),
            .I(N__35294));
    LocalMux I__6947 (
            .O(N__35366),
            .I(N__35281));
    LocalMux I__6946 (
            .O(N__35363),
            .I(N__35281));
    Span4Mux_h I__6945 (
            .O(N__35360),
            .I(N__35281));
    Span4Mux_h I__6944 (
            .O(N__35353),
            .I(N__35281));
    Span4Mux_h I__6943 (
            .O(N__35350),
            .I(N__35281));
    Span4Mux_v I__6942 (
            .O(N__35339),
            .I(N__35281));
    LocalMux I__6941 (
            .O(N__35326),
            .I(N__35278));
    InMux I__6940 (
            .O(N__35325),
            .I(N__35273));
    InMux I__6939 (
            .O(N__35324),
            .I(N__35273));
    LocalMux I__6938 (
            .O(N__35321),
            .I(adc_state_0));
    LocalMux I__6937 (
            .O(N__35318),
            .I(adc_state_0));
    LocalMux I__6936 (
            .O(N__35315),
            .I(adc_state_0));
    LocalMux I__6935 (
            .O(N__35312),
            .I(adc_state_0));
    LocalMux I__6934 (
            .O(N__35309),
            .I(adc_state_0));
    Odrv4 I__6933 (
            .O(N__35304),
            .I(adc_state_0));
    LocalMux I__6932 (
            .O(N__35301),
            .I(adc_state_0));
    Odrv4 I__6931 (
            .O(N__35294),
            .I(adc_state_0));
    Odrv4 I__6930 (
            .O(N__35281),
            .I(adc_state_0));
    Odrv4 I__6929 (
            .O(N__35278),
            .I(adc_state_0));
    LocalMux I__6928 (
            .O(N__35273),
            .I(adc_state_0));
    CascadeMux I__6927 (
            .O(N__35250),
            .I(N__35247));
    InMux I__6926 (
            .O(N__35247),
            .I(N__35244));
    LocalMux I__6925 (
            .O(N__35244),
            .I(N__35241));
    Span4Mux_v I__6924 (
            .O(N__35241),
            .I(N__35237));
    InMux I__6923 (
            .O(N__35240),
            .I(N__35234));
    Span4Mux_h I__6922 (
            .O(N__35237),
            .I(N__35228));
    LocalMux I__6921 (
            .O(N__35234),
            .I(N__35228));
    CascadeMux I__6920 (
            .O(N__35233),
            .I(N__35225));
    Span4Mux_h I__6919 (
            .O(N__35228),
            .I(N__35222));
    InMux I__6918 (
            .O(N__35225),
            .I(N__35219));
    Odrv4 I__6917 (
            .O(N__35222),
            .I(cmd_rdadctmp_21));
    LocalMux I__6916 (
            .O(N__35219),
            .I(cmd_rdadctmp_21));
    InMux I__6915 (
            .O(N__35214),
            .I(N__35211));
    LocalMux I__6914 (
            .O(N__35211),
            .I(N__35208));
    Span4Mux_v I__6913 (
            .O(N__35208),
            .I(N__35205));
    Span4Mux_h I__6912 (
            .O(N__35205),
            .I(N__35202));
    Span4Mux_v I__6911 (
            .O(N__35202),
            .I(N__35199));
    Odrv4 I__6910 (
            .O(N__35199),
            .I(buf_data_iac_21));
    CascadeMux I__6909 (
            .O(N__35196),
            .I(N__35193));
    InMux I__6908 (
            .O(N__35193),
            .I(N__35190));
    LocalMux I__6907 (
            .O(N__35190),
            .I(N__35187));
    Span4Mux_v I__6906 (
            .O(N__35187),
            .I(N__35184));
    Span4Mux_h I__6905 (
            .O(N__35184),
            .I(N__35181));
    Odrv4 I__6904 (
            .O(N__35181),
            .I(n21124));
    InMux I__6903 (
            .O(N__35178),
            .I(N__35173));
    InMux I__6902 (
            .O(N__35177),
            .I(N__35169));
    InMux I__6901 (
            .O(N__35176),
            .I(N__35166));
    LocalMux I__6900 (
            .O(N__35173),
            .I(N__35162));
    InMux I__6899 (
            .O(N__35172),
            .I(N__35159));
    LocalMux I__6898 (
            .O(N__35169),
            .I(N__35156));
    LocalMux I__6897 (
            .O(N__35166),
            .I(N__35153));
    InMux I__6896 (
            .O(N__35165),
            .I(N__35150));
    Span4Mux_h I__6895 (
            .O(N__35162),
            .I(N__35147));
    LocalMux I__6894 (
            .O(N__35159),
            .I(N__35143));
    Span4Mux_h I__6893 (
            .O(N__35156),
            .I(N__35140));
    Span4Mux_h I__6892 (
            .O(N__35153),
            .I(N__35137));
    LocalMux I__6891 (
            .O(N__35150),
            .I(N__35134));
    Span4Mux_v I__6890 (
            .O(N__35147),
            .I(N__35131));
    InMux I__6889 (
            .O(N__35146),
            .I(N__35128));
    Span4Mux_h I__6888 (
            .O(N__35143),
            .I(N__35125));
    Span4Mux_h I__6887 (
            .O(N__35140),
            .I(N__35120));
    Span4Mux_v I__6886 (
            .O(N__35137),
            .I(N__35120));
    Odrv12 I__6885 (
            .O(N__35134),
            .I(\comm_spi.n14603 ));
    Odrv4 I__6884 (
            .O(N__35131),
            .I(\comm_spi.n14603 ));
    LocalMux I__6883 (
            .O(N__35128),
            .I(\comm_spi.n14603 ));
    Odrv4 I__6882 (
            .O(N__35125),
            .I(\comm_spi.n14603 ));
    Odrv4 I__6881 (
            .O(N__35120),
            .I(\comm_spi.n14603 ));
    SRMux I__6880 (
            .O(N__35109),
            .I(N__35104));
    SRMux I__6879 (
            .O(N__35108),
            .I(N__35101));
    SRMux I__6878 (
            .O(N__35107),
            .I(N__35098));
    LocalMux I__6877 (
            .O(N__35104),
            .I(N__35095));
    LocalMux I__6876 (
            .O(N__35101),
            .I(N__35092));
    LocalMux I__6875 (
            .O(N__35098),
            .I(N__35089));
    Span4Mux_h I__6874 (
            .O(N__35095),
            .I(N__35086));
    Span4Mux_v I__6873 (
            .O(N__35092),
            .I(N__35083));
    Span4Mux_h I__6872 (
            .O(N__35089),
            .I(N__35080));
    Span4Mux_v I__6871 (
            .O(N__35086),
            .I(N__35077));
    Span4Mux_h I__6870 (
            .O(N__35083),
            .I(N__35072));
    Span4Mux_v I__6869 (
            .O(N__35080),
            .I(N__35072));
    Odrv4 I__6868 (
            .O(N__35077),
            .I(\comm_spi.data_tx_7__N_774 ));
    Odrv4 I__6867 (
            .O(N__35072),
            .I(\comm_spi.data_tx_7__N_774 ));
    InMux I__6866 (
            .O(N__35067),
            .I(N__35062));
    InMux I__6865 (
            .O(N__35066),
            .I(N__35057));
    InMux I__6864 (
            .O(N__35065),
            .I(N__35057));
    LocalMux I__6863 (
            .O(N__35062),
            .I(N__35052));
    LocalMux I__6862 (
            .O(N__35057),
            .I(N__35052));
    Odrv4 I__6861 (
            .O(N__35052),
            .I(comm_tx_buf_7));
    SRMux I__6860 (
            .O(N__35049),
            .I(N__35046));
    LocalMux I__6859 (
            .O(N__35046),
            .I(N__35041));
    SRMux I__6858 (
            .O(N__35045),
            .I(N__35038));
    SRMux I__6857 (
            .O(N__35044),
            .I(N__35035));
    Span4Mux_v I__6856 (
            .O(N__35041),
            .I(N__35032));
    LocalMux I__6855 (
            .O(N__35038),
            .I(N__35029));
    LocalMux I__6854 (
            .O(N__35035),
            .I(N__35026));
    Span4Mux_v I__6853 (
            .O(N__35032),
            .I(N__35023));
    Span4Mux_h I__6852 (
            .O(N__35029),
            .I(N__35020));
    Span4Mux_v I__6851 (
            .O(N__35026),
            .I(N__35017));
    Span4Mux_v I__6850 (
            .O(N__35023),
            .I(N__35014));
    Span4Mux_h I__6849 (
            .O(N__35020),
            .I(N__35011));
    Odrv4 I__6848 (
            .O(N__35017),
            .I(\comm_spi.data_tx_7__N_766 ));
    Odrv4 I__6847 (
            .O(N__35014),
            .I(\comm_spi.data_tx_7__N_766 ));
    Odrv4 I__6846 (
            .O(N__35011),
            .I(\comm_spi.data_tx_7__N_766 ));
    InMux I__6845 (
            .O(N__35004),
            .I(N__34998));
    InMux I__6844 (
            .O(N__35003),
            .I(N__34998));
    LocalMux I__6843 (
            .O(N__34998),
            .I(N__34990));
    InMux I__6842 (
            .O(N__34997),
            .I(N__34987));
    InMux I__6841 (
            .O(N__34996),
            .I(N__34980));
    InMux I__6840 (
            .O(N__34995),
            .I(N__34980));
    InMux I__6839 (
            .O(N__34994),
            .I(N__34980));
    InMux I__6838 (
            .O(N__34993),
            .I(N__34977));
    Odrv4 I__6837 (
            .O(N__34990),
            .I(n12228));
    LocalMux I__6836 (
            .O(N__34987),
            .I(n12228));
    LocalMux I__6835 (
            .O(N__34980),
            .I(n12228));
    LocalMux I__6834 (
            .O(N__34977),
            .I(n12228));
    InMux I__6833 (
            .O(N__34968),
            .I(N__34965));
    LocalMux I__6832 (
            .O(N__34965),
            .I(N__34962));
    Span4Mux_v I__6831 (
            .O(N__34962),
            .I(N__34959));
    Span4Mux_v I__6830 (
            .O(N__34959),
            .I(N__34955));
    CascadeMux I__6829 (
            .O(N__34958),
            .I(N__34952));
    Span4Mux_h I__6828 (
            .O(N__34955),
            .I(N__34949));
    InMux I__6827 (
            .O(N__34952),
            .I(N__34946));
    Odrv4 I__6826 (
            .O(N__34949),
            .I(buf_adcdata_vdc_9));
    LocalMux I__6825 (
            .O(N__34946),
            .I(buf_adcdata_vdc_9));
    InMux I__6824 (
            .O(N__34941),
            .I(N__34938));
    LocalMux I__6823 (
            .O(N__34938),
            .I(N__34934));
    InMux I__6822 (
            .O(N__34937),
            .I(N__34930));
    Span4Mux_h I__6821 (
            .O(N__34934),
            .I(N__34927));
    CascadeMux I__6820 (
            .O(N__34933),
            .I(N__34924));
    LocalMux I__6819 (
            .O(N__34930),
            .I(N__34921));
    Sp12to4 I__6818 (
            .O(N__34927),
            .I(N__34918));
    InMux I__6817 (
            .O(N__34924),
            .I(N__34915));
    Span4Mux_v I__6816 (
            .O(N__34921),
            .I(N__34912));
    Span12Mux_v I__6815 (
            .O(N__34918),
            .I(N__34909));
    LocalMux I__6814 (
            .O(N__34915),
            .I(buf_adcdata_vac_9));
    Odrv4 I__6813 (
            .O(N__34912),
            .I(buf_adcdata_vac_9));
    Odrv12 I__6812 (
            .O(N__34909),
            .I(buf_adcdata_vac_9));
    InMux I__6811 (
            .O(N__34902),
            .I(N__34898));
    InMux I__6810 (
            .O(N__34901),
            .I(N__34894));
    LocalMux I__6809 (
            .O(N__34898),
            .I(N__34891));
    InMux I__6808 (
            .O(N__34897),
            .I(N__34888));
    LocalMux I__6807 (
            .O(N__34894),
            .I(N__34881));
    Span4Mux_h I__6806 (
            .O(N__34891),
            .I(N__34881));
    LocalMux I__6805 (
            .O(N__34888),
            .I(N__34881));
    Odrv4 I__6804 (
            .O(N__34881),
            .I(comm_tx_buf_3));
    CascadeMux I__6803 (
            .O(N__34878),
            .I(n21122_cascade_));
    CascadeMux I__6802 (
            .O(N__34875),
            .I(N__34872));
    InMux I__6801 (
            .O(N__34872),
            .I(N__34869));
    LocalMux I__6800 (
            .O(N__34869),
            .I(n21120));
    CEMux I__6799 (
            .O(N__34866),
            .I(N__34863));
    LocalMux I__6798 (
            .O(N__34863),
            .I(N__34860));
    Odrv4 I__6797 (
            .O(N__34860),
            .I(n11361));
    CascadeMux I__6796 (
            .O(N__34857),
            .I(n7_adj_1616_cascade_));
    CascadeMux I__6795 (
            .O(N__34854),
            .I(N__34851));
    InMux I__6794 (
            .O(N__34851),
            .I(N__34848));
    LocalMux I__6793 (
            .O(N__34848),
            .I(\ADC_VDC.n17509 ));
    InMux I__6792 (
            .O(N__34845),
            .I(N__34842));
    LocalMux I__6791 (
            .O(N__34842),
            .I(\ADC_VDC.n11265 ));
    InMux I__6790 (
            .O(N__34839),
            .I(N__34836));
    LocalMux I__6789 (
            .O(N__34836),
            .I(\ADC_VDC.n6 ));
    CascadeMux I__6788 (
            .O(N__34833),
            .I(\ADC_VDC.n11265_cascade_ ));
    InMux I__6787 (
            .O(N__34830),
            .I(N__34827));
    LocalMux I__6786 (
            .O(N__34827),
            .I(N__34823));
    InMux I__6785 (
            .O(N__34826),
            .I(N__34820));
    Span4Mux_h I__6784 (
            .O(N__34823),
            .I(N__34817));
    LocalMux I__6783 (
            .O(N__34820),
            .I(N__34814));
    Odrv4 I__6782 (
            .O(N__34817),
            .I(\ADC_VDC.n15 ));
    Odrv4 I__6781 (
            .O(N__34814),
            .I(\ADC_VDC.n15 ));
    CascadeMux I__6780 (
            .O(N__34809),
            .I(\ADC_VDC.n15_cascade_ ));
    InMux I__6779 (
            .O(N__34806),
            .I(N__34803));
    LocalMux I__6778 (
            .O(N__34803),
            .I(N__34800));
    Odrv4 I__6777 (
            .O(N__34800),
            .I(\ADC_VDC.n20996 ));
    CascadeMux I__6776 (
            .O(N__34797),
            .I(N__34777));
    InMux I__6775 (
            .O(N__34796),
            .I(N__34773));
    InMux I__6774 (
            .O(N__34795),
            .I(N__34768));
    InMux I__6773 (
            .O(N__34794),
            .I(N__34753));
    InMux I__6772 (
            .O(N__34793),
            .I(N__34753));
    InMux I__6771 (
            .O(N__34792),
            .I(N__34753));
    InMux I__6770 (
            .O(N__34791),
            .I(N__34753));
    InMux I__6769 (
            .O(N__34790),
            .I(N__34753));
    InMux I__6768 (
            .O(N__34789),
            .I(N__34753));
    InMux I__6767 (
            .O(N__34788),
            .I(N__34753));
    InMux I__6766 (
            .O(N__34787),
            .I(N__34732));
    InMux I__6765 (
            .O(N__34786),
            .I(N__34732));
    InMux I__6764 (
            .O(N__34785),
            .I(N__34732));
    InMux I__6763 (
            .O(N__34784),
            .I(N__34732));
    InMux I__6762 (
            .O(N__34783),
            .I(N__34732));
    InMux I__6761 (
            .O(N__34782),
            .I(N__34732));
    InMux I__6760 (
            .O(N__34781),
            .I(N__34732));
    InMux I__6759 (
            .O(N__34780),
            .I(N__34732));
    InMux I__6758 (
            .O(N__34777),
            .I(N__34727));
    InMux I__6757 (
            .O(N__34776),
            .I(N__34727));
    LocalMux I__6756 (
            .O(N__34773),
            .I(N__34724));
    SRMux I__6755 (
            .O(N__34772),
            .I(N__34721));
    InMux I__6754 (
            .O(N__34771),
            .I(N__34718));
    LocalMux I__6753 (
            .O(N__34768),
            .I(N__34715));
    LocalMux I__6752 (
            .O(N__34753),
            .I(N__34712));
    CascadeMux I__6751 (
            .O(N__34752),
            .I(N__34707));
    CEMux I__6750 (
            .O(N__34751),
            .I(N__34703));
    InMux I__6749 (
            .O(N__34750),
            .I(N__34700));
    InMux I__6748 (
            .O(N__34749),
            .I(N__34697));
    LocalMux I__6747 (
            .O(N__34732),
            .I(N__34692));
    LocalMux I__6746 (
            .O(N__34727),
            .I(N__34692));
    Span4Mux_v I__6745 (
            .O(N__34724),
            .I(N__34687));
    LocalMux I__6744 (
            .O(N__34721),
            .I(N__34687));
    LocalMux I__6743 (
            .O(N__34718),
            .I(N__34684));
    Span4Mux_v I__6742 (
            .O(N__34715),
            .I(N__34679));
    Span4Mux_v I__6741 (
            .O(N__34712),
            .I(N__34679));
    InMux I__6740 (
            .O(N__34711),
            .I(N__34676));
    InMux I__6739 (
            .O(N__34710),
            .I(N__34673));
    InMux I__6738 (
            .O(N__34707),
            .I(N__34670));
    InMux I__6737 (
            .O(N__34706),
            .I(N__34667));
    LocalMux I__6736 (
            .O(N__34703),
            .I(N__34664));
    LocalMux I__6735 (
            .O(N__34700),
            .I(N__34661));
    LocalMux I__6734 (
            .O(N__34697),
            .I(N__34656));
    Span4Mux_v I__6733 (
            .O(N__34692),
            .I(N__34656));
    Span4Mux_h I__6732 (
            .O(N__34687),
            .I(N__34651));
    Span4Mux_v I__6731 (
            .O(N__34684),
            .I(N__34651));
    Span4Mux_h I__6730 (
            .O(N__34679),
            .I(N__34646));
    LocalMux I__6729 (
            .O(N__34676),
            .I(N__34646));
    LocalMux I__6728 (
            .O(N__34673),
            .I(N__34643));
    LocalMux I__6727 (
            .O(N__34670),
            .I(N__34638));
    LocalMux I__6726 (
            .O(N__34667),
            .I(N__34638));
    Span4Mux_v I__6725 (
            .O(N__34664),
            .I(N__34629));
    Span4Mux_h I__6724 (
            .O(N__34661),
            .I(N__34629));
    Span4Mux_v I__6723 (
            .O(N__34656),
            .I(N__34629));
    Span4Mux_h I__6722 (
            .O(N__34651),
            .I(N__34629));
    Odrv4 I__6721 (
            .O(N__34646),
            .I(dds_state_1_adj_1453));
    Odrv4 I__6720 (
            .O(N__34643),
            .I(dds_state_1_adj_1453));
    Odrv12 I__6719 (
            .O(N__34638),
            .I(dds_state_1_adj_1453));
    Odrv4 I__6718 (
            .O(N__34629),
            .I(dds_state_1_adj_1453));
    InMux I__6717 (
            .O(N__34620),
            .I(N__34606));
    CascadeMux I__6716 (
            .O(N__34619),
            .I(N__34603));
    InMux I__6715 (
            .O(N__34618),
            .I(N__34577));
    InMux I__6714 (
            .O(N__34617),
            .I(N__34577));
    InMux I__6713 (
            .O(N__34616),
            .I(N__34577));
    InMux I__6712 (
            .O(N__34615),
            .I(N__34577));
    InMux I__6711 (
            .O(N__34614),
            .I(N__34577));
    InMux I__6710 (
            .O(N__34613),
            .I(N__34577));
    InMux I__6709 (
            .O(N__34612),
            .I(N__34577));
    InMux I__6708 (
            .O(N__34611),
            .I(N__34577));
    InMux I__6707 (
            .O(N__34610),
            .I(N__34574));
    InMux I__6706 (
            .O(N__34609),
            .I(N__34571));
    LocalMux I__6705 (
            .O(N__34606),
            .I(N__34568));
    InMux I__6704 (
            .O(N__34603),
            .I(N__34564));
    InMux I__6703 (
            .O(N__34602),
            .I(N__34549));
    InMux I__6702 (
            .O(N__34601),
            .I(N__34549));
    InMux I__6701 (
            .O(N__34600),
            .I(N__34549));
    InMux I__6700 (
            .O(N__34599),
            .I(N__34549));
    InMux I__6699 (
            .O(N__34598),
            .I(N__34549));
    InMux I__6698 (
            .O(N__34597),
            .I(N__34549));
    InMux I__6697 (
            .O(N__34596),
            .I(N__34549));
    InMux I__6696 (
            .O(N__34595),
            .I(N__34542));
    InMux I__6695 (
            .O(N__34594),
            .I(N__34542));
    LocalMux I__6694 (
            .O(N__34577),
            .I(N__34537));
    LocalMux I__6693 (
            .O(N__34574),
            .I(N__34537));
    LocalMux I__6692 (
            .O(N__34571),
            .I(N__34533));
    Span4Mux_h I__6691 (
            .O(N__34568),
            .I(N__34530));
    InMux I__6690 (
            .O(N__34567),
            .I(N__34526));
    LocalMux I__6689 (
            .O(N__34564),
            .I(N__34521));
    LocalMux I__6688 (
            .O(N__34549),
            .I(N__34521));
    InMux I__6687 (
            .O(N__34548),
            .I(N__34518));
    InMux I__6686 (
            .O(N__34547),
            .I(N__34515));
    LocalMux I__6685 (
            .O(N__34542),
            .I(N__34512));
    Span4Mux_v I__6684 (
            .O(N__34537),
            .I(N__34509));
    InMux I__6683 (
            .O(N__34536),
            .I(N__34506));
    Span4Mux_v I__6682 (
            .O(N__34533),
            .I(N__34501));
    Span4Mux_h I__6681 (
            .O(N__34530),
            .I(N__34501));
    InMux I__6680 (
            .O(N__34529),
            .I(N__34498));
    LocalMux I__6679 (
            .O(N__34526),
            .I(N__34495));
    Span12Mux_v I__6678 (
            .O(N__34521),
            .I(N__34492));
    LocalMux I__6677 (
            .O(N__34518),
            .I(N__34489));
    LocalMux I__6676 (
            .O(N__34515),
            .I(N__34484));
    Span4Mux_v I__6675 (
            .O(N__34512),
            .I(N__34484));
    Span4Mux_h I__6674 (
            .O(N__34509),
            .I(N__34477));
    LocalMux I__6673 (
            .O(N__34506),
            .I(N__34477));
    Span4Mux_h I__6672 (
            .O(N__34501),
            .I(N__34477));
    LocalMux I__6671 (
            .O(N__34498),
            .I(dds_state_2_adj_1452));
    Odrv4 I__6670 (
            .O(N__34495),
            .I(dds_state_2_adj_1452));
    Odrv12 I__6669 (
            .O(N__34492),
            .I(dds_state_2_adj_1452));
    Odrv4 I__6668 (
            .O(N__34489),
            .I(dds_state_2_adj_1452));
    Odrv4 I__6667 (
            .O(N__34484),
            .I(dds_state_2_adj_1452));
    Odrv4 I__6666 (
            .O(N__34477),
            .I(dds_state_2_adj_1452));
    InMux I__6665 (
            .O(N__34464),
            .I(N__34460));
    InMux I__6664 (
            .O(N__34463),
            .I(N__34454));
    LocalMux I__6663 (
            .O(N__34460),
            .I(N__34450));
    InMux I__6662 (
            .O(N__34459),
            .I(N__34447));
    InMux I__6661 (
            .O(N__34458),
            .I(N__34444));
    InMux I__6660 (
            .O(N__34457),
            .I(N__34441));
    LocalMux I__6659 (
            .O(N__34454),
            .I(N__34438));
    InMux I__6658 (
            .O(N__34453),
            .I(N__34434));
    Span4Mux_h I__6657 (
            .O(N__34450),
            .I(N__34431));
    LocalMux I__6656 (
            .O(N__34447),
            .I(N__34426));
    LocalMux I__6655 (
            .O(N__34444),
            .I(N__34426));
    LocalMux I__6654 (
            .O(N__34441),
            .I(N__34420));
    Span4Mux_h I__6653 (
            .O(N__34438),
            .I(N__34417));
    InMux I__6652 (
            .O(N__34437),
            .I(N__34414));
    LocalMux I__6651 (
            .O(N__34434),
            .I(N__34407));
    Span4Mux_h I__6650 (
            .O(N__34431),
            .I(N__34407));
    Span4Mux_v I__6649 (
            .O(N__34426),
            .I(N__34407));
    InMux I__6648 (
            .O(N__34425),
            .I(N__34404));
    InMux I__6647 (
            .O(N__34424),
            .I(N__34399));
    InMux I__6646 (
            .O(N__34423),
            .I(N__34399));
    Odrv4 I__6645 (
            .O(N__34420),
            .I(dds_state_0_adj_1454));
    Odrv4 I__6644 (
            .O(N__34417),
            .I(dds_state_0_adj_1454));
    LocalMux I__6643 (
            .O(N__34414),
            .I(dds_state_0_adj_1454));
    Odrv4 I__6642 (
            .O(N__34407),
            .I(dds_state_0_adj_1454));
    LocalMux I__6641 (
            .O(N__34404),
            .I(dds_state_0_adj_1454));
    LocalMux I__6640 (
            .O(N__34399),
            .I(dds_state_0_adj_1454));
    CEMux I__6639 (
            .O(N__34386),
            .I(N__34383));
    LocalMux I__6638 (
            .O(N__34383),
            .I(N__34379));
    CEMux I__6637 (
            .O(N__34382),
            .I(N__34376));
    Span4Mux_v I__6636 (
            .O(N__34379),
            .I(N__34373));
    LocalMux I__6635 (
            .O(N__34376),
            .I(N__34370));
    Span4Mux_h I__6634 (
            .O(N__34373),
            .I(N__34367));
    Span12Mux_v I__6633 (
            .O(N__34370),
            .I(N__34364));
    Odrv4 I__6632 (
            .O(N__34367),
            .I(\CLK_DDS.n12784 ));
    Odrv12 I__6631 (
            .O(N__34364),
            .I(\CLK_DDS.n12784 ));
    InMux I__6630 (
            .O(N__34359),
            .I(N__34356));
    LocalMux I__6629 (
            .O(N__34356),
            .I(N__34353));
    Span4Mux_v I__6628 (
            .O(N__34353),
            .I(N__34349));
    InMux I__6627 (
            .O(N__34352),
            .I(N__34346));
    Span4Mux_v I__6626 (
            .O(N__34349),
            .I(N__34341));
    LocalMux I__6625 (
            .O(N__34346),
            .I(N__34341));
    Odrv4 I__6624 (
            .O(N__34341),
            .I(\comm_spi.n14607 ));
    InMux I__6623 (
            .O(N__34338),
            .I(N__34335));
    LocalMux I__6622 (
            .O(N__34335),
            .I(\ADC_VDC.n19_adj_1401 ));
    CascadeMux I__6621 (
            .O(N__34332),
            .I(\ADC_VDC.n21323_cascade_ ));
    InMux I__6620 (
            .O(N__34329),
            .I(N__34326));
    LocalMux I__6619 (
            .O(N__34326),
            .I(\ADC_VDC.n21320 ));
    InMux I__6618 (
            .O(N__34323),
            .I(N__34320));
    LocalMux I__6617 (
            .O(N__34320),
            .I(N__34317));
    Odrv4 I__6616 (
            .O(N__34317),
            .I(\ADC_VDC.n20965 ));
    CascadeMux I__6615 (
            .O(N__34314),
            .I(\ADC_VDC.n10_cascade_ ));
    InMux I__6614 (
            .O(N__34311),
            .I(N__34308));
    LocalMux I__6613 (
            .O(N__34308),
            .I(\ADC_VDC.n20812 ));
    InMux I__6612 (
            .O(N__34305),
            .I(N__34302));
    LocalMux I__6611 (
            .O(N__34302),
            .I(\ADC_VDC.n20784 ));
    CascadeMux I__6610 (
            .O(N__34299),
            .I(n8_adj_1573_cascade_));
    InMux I__6609 (
            .O(N__34296),
            .I(N__34292));
    InMux I__6608 (
            .O(N__34295),
            .I(N__34289));
    LocalMux I__6607 (
            .O(N__34292),
            .I(N__34286));
    LocalMux I__6606 (
            .O(N__34289),
            .I(N__34281));
    Span4Mux_v I__6605 (
            .O(N__34286),
            .I(N__34278));
    InMux I__6604 (
            .O(N__34285),
            .I(N__34273));
    InMux I__6603 (
            .O(N__34284),
            .I(N__34273));
    Odrv4 I__6602 (
            .O(N__34281),
            .I(eis_stop));
    Odrv4 I__6601 (
            .O(N__34278),
            .I(eis_stop));
    LocalMux I__6600 (
            .O(N__34273),
            .I(eis_stop));
    InMux I__6599 (
            .O(N__34266),
            .I(N__34262));
    InMux I__6598 (
            .O(N__34265),
            .I(N__34258));
    LocalMux I__6597 (
            .O(N__34262),
            .I(N__34255));
    InMux I__6596 (
            .O(N__34261),
            .I(N__34252));
    LocalMux I__6595 (
            .O(N__34258),
            .I(req_data_cnt_9));
    Odrv4 I__6594 (
            .O(N__34255),
            .I(req_data_cnt_9));
    LocalMux I__6593 (
            .O(N__34252),
            .I(req_data_cnt_9));
    InMux I__6592 (
            .O(N__34245),
            .I(N__34242));
    LocalMux I__6591 (
            .O(N__34242),
            .I(n22375));
    CascadeMux I__6590 (
            .O(N__34239),
            .I(N__34236));
    InMux I__6589 (
            .O(N__34236),
            .I(N__34233));
    LocalMux I__6588 (
            .O(N__34233),
            .I(N__34230));
    Span4Mux_v I__6587 (
            .O(N__34230),
            .I(N__34227));
    Span4Mux_v I__6586 (
            .O(N__34227),
            .I(N__34224));
    Odrv4 I__6585 (
            .O(N__34224),
            .I(n22381));
    InMux I__6584 (
            .O(N__34221),
            .I(N__34218));
    LocalMux I__6583 (
            .O(N__34218),
            .I(N__34215));
    Span4Mux_v I__6582 (
            .O(N__34215),
            .I(N__34212));
    Span4Mux_v I__6581 (
            .O(N__34212),
            .I(N__34209));
    Odrv4 I__6580 (
            .O(N__34209),
            .I(n22384));
    InMux I__6579 (
            .O(N__34206),
            .I(N__34203));
    LocalMux I__6578 (
            .O(N__34203),
            .I(N__34200));
    Odrv4 I__6577 (
            .O(N__34200),
            .I(n11396));
    IoInMux I__6576 (
            .O(N__34197),
            .I(N__34194));
    LocalMux I__6575 (
            .O(N__34194),
            .I(N__34191));
    IoSpan4Mux I__6574 (
            .O(N__34191),
            .I(N__34188));
    IoSpan4Mux I__6573 (
            .O(N__34188),
            .I(N__34185));
    Span4Mux_s3_v I__6572 (
            .O(N__34185),
            .I(N__34182));
    Span4Mux_h I__6571 (
            .O(N__34182),
            .I(N__34179));
    Span4Mux_v I__6570 (
            .O(N__34179),
            .I(N__34175));
    InMux I__6569 (
            .O(N__34178),
            .I(N__34172));
    Odrv4 I__6568 (
            .O(N__34175),
            .I(DDS_SCK));
    LocalMux I__6567 (
            .O(N__34172),
            .I(DDS_SCK));
    InMux I__6566 (
            .O(N__34167),
            .I(N__34164));
    LocalMux I__6565 (
            .O(N__34164),
            .I(N__34161));
    Span4Mux_v I__6564 (
            .O(N__34161),
            .I(N__34158));
    Odrv4 I__6563 (
            .O(N__34158),
            .I(\comm_spi.n14605 ));
    InMux I__6562 (
            .O(N__34155),
            .I(N__34152));
    LocalMux I__6561 (
            .O(N__34152),
            .I(N__34149));
    Span4Mux_h I__6560 (
            .O(N__34149),
            .I(N__34146));
    Odrv4 I__6559 (
            .O(N__34146),
            .I(\comm_spi.n14604 ));
    IoInMux I__6558 (
            .O(N__34143),
            .I(N__34140));
    LocalMux I__6557 (
            .O(N__34140),
            .I(N__34137));
    IoSpan4Mux I__6556 (
            .O(N__34137),
            .I(N__34134));
    Span4Mux_s3_h I__6555 (
            .O(N__34134),
            .I(N__34131));
    Sp12to4 I__6554 (
            .O(N__34131),
            .I(N__34128));
    Span12Mux_h I__6553 (
            .O(N__34128),
            .I(N__34125));
    Odrv12 I__6552 (
            .O(N__34125),
            .I(ICE_SPI_MISO));
    InMux I__6551 (
            .O(N__34122),
            .I(N__34119));
    LocalMux I__6550 (
            .O(N__34119),
            .I(n20_adj_1617));
    InMux I__6549 (
            .O(N__34116),
            .I(N__34113));
    LocalMux I__6548 (
            .O(N__34113),
            .I(N__34108));
    InMux I__6547 (
            .O(N__34112),
            .I(N__34105));
    InMux I__6546 (
            .O(N__34111),
            .I(N__34102));
    Span4Mux_h I__6545 (
            .O(N__34108),
            .I(N__34099));
    LocalMux I__6544 (
            .O(N__34105),
            .I(N__34094));
    LocalMux I__6543 (
            .O(N__34102),
            .I(N__34094));
    Odrv4 I__6542 (
            .O(N__34099),
            .I(n10717));
    Odrv12 I__6541 (
            .O(N__34094),
            .I(n10717));
    InMux I__6540 (
            .O(N__34089),
            .I(N__34084));
    InMux I__6539 (
            .O(N__34088),
            .I(N__34079));
    InMux I__6538 (
            .O(N__34087),
            .I(N__34079));
    LocalMux I__6537 (
            .O(N__34084),
            .I(req_data_cnt_12));
    LocalMux I__6536 (
            .O(N__34079),
            .I(req_data_cnt_12));
    CascadeMux I__6535 (
            .O(N__34074),
            .I(N__34069));
    InMux I__6534 (
            .O(N__34073),
            .I(N__34066));
    InMux I__6533 (
            .O(N__34072),
            .I(N__34063));
    InMux I__6532 (
            .O(N__34069),
            .I(N__34060));
    LocalMux I__6531 (
            .O(N__34066),
            .I(acadc_skipCount_9));
    LocalMux I__6530 (
            .O(N__34063),
            .I(acadc_skipCount_9));
    LocalMux I__6529 (
            .O(N__34060),
            .I(acadc_skipCount_9));
    InMux I__6528 (
            .O(N__34053),
            .I(N__34050));
    LocalMux I__6527 (
            .O(N__34050),
            .I(N__34047));
    Odrv12 I__6526 (
            .O(N__34047),
            .I(n19_adj_1607));
    CascadeMux I__6525 (
            .O(N__34044),
            .I(n29_cascade_));
    CascadeMux I__6524 (
            .O(N__34041),
            .I(N__34038));
    InMux I__6523 (
            .O(N__34038),
            .I(N__34034));
    InMux I__6522 (
            .O(N__34037),
            .I(N__34031));
    LocalMux I__6521 (
            .O(N__34034),
            .I(N__34025));
    LocalMux I__6520 (
            .O(N__34031),
            .I(N__34025));
    InMux I__6519 (
            .O(N__34030),
            .I(N__34022));
    Span4Mux_v I__6518 (
            .O(N__34025),
            .I(N__34019));
    LocalMux I__6517 (
            .O(N__34022),
            .I(n16_adj_1603));
    Odrv4 I__6516 (
            .O(N__34019),
            .I(n16_adj_1603));
    InMux I__6515 (
            .O(N__34014),
            .I(N__34011));
    LocalMux I__6514 (
            .O(N__34011),
            .I(n24));
    CascadeMux I__6513 (
            .O(N__34008),
            .I(n21_adj_1492_cascade_));
    InMux I__6512 (
            .O(N__34005),
            .I(N__34002));
    LocalMux I__6511 (
            .O(N__34002),
            .I(n30_adj_1618));
    InMux I__6510 (
            .O(N__33999),
            .I(N__33996));
    LocalMux I__6509 (
            .O(N__33996),
            .I(N__33993));
    Span4Mux_v I__6508 (
            .O(N__33993),
            .I(N__33989));
    InMux I__6507 (
            .O(N__33992),
            .I(N__33985));
    Span4Mux_h I__6506 (
            .O(N__33989),
            .I(N__33982));
    InMux I__6505 (
            .O(N__33988),
            .I(N__33979));
    LocalMux I__6504 (
            .O(N__33985),
            .I(buf_dds1_4));
    Odrv4 I__6503 (
            .O(N__33982),
            .I(buf_dds1_4));
    LocalMux I__6502 (
            .O(N__33979),
            .I(buf_dds1_4));
    CascadeMux I__6501 (
            .O(N__33972),
            .I(N__33969));
    InMux I__6500 (
            .O(N__33969),
            .I(N__33964));
    InMux I__6499 (
            .O(N__33968),
            .I(N__33961));
    InMux I__6498 (
            .O(N__33967),
            .I(N__33958));
    LocalMux I__6497 (
            .O(N__33964),
            .I(N__33953));
    LocalMux I__6496 (
            .O(N__33961),
            .I(N__33953));
    LocalMux I__6495 (
            .O(N__33958),
            .I(buf_dds0_0));
    Odrv4 I__6494 (
            .O(N__33953),
            .I(buf_dds0_0));
    InMux I__6493 (
            .O(N__33948),
            .I(N__33945));
    LocalMux I__6492 (
            .O(N__33945),
            .I(N__33941));
    InMux I__6491 (
            .O(N__33944),
            .I(N__33937));
    Span4Mux_h I__6490 (
            .O(N__33941),
            .I(N__33934));
    InMux I__6489 (
            .O(N__33940),
            .I(N__33931));
    LocalMux I__6488 (
            .O(N__33937),
            .I(req_data_cnt_13));
    Odrv4 I__6487 (
            .O(N__33934),
            .I(req_data_cnt_13));
    LocalMux I__6486 (
            .O(N__33931),
            .I(req_data_cnt_13));
    InMux I__6485 (
            .O(N__33924),
            .I(N__33920));
    InMux I__6484 (
            .O(N__33923),
            .I(N__33916));
    LocalMux I__6483 (
            .O(N__33920),
            .I(N__33913));
    InMux I__6482 (
            .O(N__33919),
            .I(N__33910));
    LocalMux I__6481 (
            .O(N__33916),
            .I(buf_dds1_0));
    Odrv12 I__6480 (
            .O(N__33913),
            .I(buf_dds1_0));
    LocalMux I__6479 (
            .O(N__33910),
            .I(buf_dds1_0));
    InMux I__6478 (
            .O(N__33903),
            .I(N__33900));
    LocalMux I__6477 (
            .O(N__33900),
            .I(n22_adj_1615));
    CascadeMux I__6476 (
            .O(N__33897),
            .I(n10717_cascade_));
    InMux I__6475 (
            .O(N__33894),
            .I(N__33891));
    LocalMux I__6474 (
            .O(N__33891),
            .I(N__33888));
    Odrv4 I__6473 (
            .O(N__33888),
            .I(n21344));
    InMux I__6472 (
            .O(N__33885),
            .I(N__33880));
    InMux I__6471 (
            .O(N__33884),
            .I(N__33877));
    InMux I__6470 (
            .O(N__33883),
            .I(N__33874));
    LocalMux I__6469 (
            .O(N__33880),
            .I(N__33871));
    LocalMux I__6468 (
            .O(N__33877),
            .I(N__33868));
    LocalMux I__6467 (
            .O(N__33874),
            .I(N__33863));
    Span4Mux_v I__6466 (
            .O(N__33871),
            .I(N__33863));
    Span4Mux_h I__6465 (
            .O(N__33868),
            .I(N__33860));
    Odrv4 I__6464 (
            .O(N__33863),
            .I(buf_dds1_5));
    Odrv4 I__6463 (
            .O(N__33860),
            .I(buf_dds1_5));
    CascadeMux I__6462 (
            .O(N__33855),
            .I(N__33852));
    InMux I__6461 (
            .O(N__33852),
            .I(N__33849));
    LocalMux I__6460 (
            .O(N__33849),
            .I(N__33844));
    InMux I__6459 (
            .O(N__33848),
            .I(N__33841));
    InMux I__6458 (
            .O(N__33847),
            .I(N__33838));
    Span4Mux_v I__6457 (
            .O(N__33844),
            .I(N__33833));
    LocalMux I__6456 (
            .O(N__33841),
            .I(N__33833));
    LocalMux I__6455 (
            .O(N__33838),
            .I(buf_dds1_7));
    Odrv4 I__6454 (
            .O(N__33833),
            .I(buf_dds1_7));
    InMux I__6453 (
            .O(N__33828),
            .I(N__33825));
    LocalMux I__6452 (
            .O(N__33825),
            .I(N__33822));
    Span4Mux_v I__6451 (
            .O(N__33822),
            .I(N__33817));
    InMux I__6450 (
            .O(N__33821),
            .I(N__33812));
    InMux I__6449 (
            .O(N__33820),
            .I(N__33812));
    Odrv4 I__6448 (
            .O(N__33817),
            .I(acadc_skipCount_14));
    LocalMux I__6447 (
            .O(N__33812),
            .I(acadc_skipCount_14));
    InMux I__6446 (
            .O(N__33807),
            .I(N__33803));
    InMux I__6445 (
            .O(N__33806),
            .I(N__33799));
    LocalMux I__6444 (
            .O(N__33803),
            .I(N__33796));
    InMux I__6443 (
            .O(N__33802),
            .I(N__33793));
    LocalMux I__6442 (
            .O(N__33799),
            .I(N__33790));
    Span4Mux_h I__6441 (
            .O(N__33796),
            .I(N__33787));
    LocalMux I__6440 (
            .O(N__33793),
            .I(buf_dds0_4));
    Odrv4 I__6439 (
            .O(N__33790),
            .I(buf_dds0_4));
    Odrv4 I__6438 (
            .O(N__33787),
            .I(buf_dds0_4));
    InMux I__6437 (
            .O(N__33780),
            .I(N__33777));
    LocalMux I__6436 (
            .O(N__33777),
            .I(N__33773));
    InMux I__6435 (
            .O(N__33776),
            .I(N__33770));
    Span4Mux_v I__6434 (
            .O(N__33773),
            .I(N__33767));
    LocalMux I__6433 (
            .O(N__33770),
            .I(comm_buf_6_3));
    Odrv4 I__6432 (
            .O(N__33767),
            .I(comm_buf_6_3));
    CascadeMux I__6431 (
            .O(N__33762),
            .I(N__33759));
    InMux I__6430 (
            .O(N__33759),
            .I(N__33755));
    InMux I__6429 (
            .O(N__33758),
            .I(N__33751));
    LocalMux I__6428 (
            .O(N__33755),
            .I(N__33748));
    InMux I__6427 (
            .O(N__33754),
            .I(N__33745));
    LocalMux I__6426 (
            .O(N__33751),
            .I(buf_dds1_1));
    Odrv4 I__6425 (
            .O(N__33748),
            .I(buf_dds1_1));
    LocalMux I__6424 (
            .O(N__33745),
            .I(buf_dds1_1));
    InMux I__6423 (
            .O(N__33738),
            .I(N__33735));
    LocalMux I__6422 (
            .O(N__33735),
            .I(N__33730));
    InMux I__6421 (
            .O(N__33734),
            .I(N__33727));
    InMux I__6420 (
            .O(N__33733),
            .I(N__33724));
    Odrv12 I__6419 (
            .O(N__33730),
            .I(cmd_rdadctmp_9_adj_1441));
    LocalMux I__6418 (
            .O(N__33727),
            .I(cmd_rdadctmp_9_adj_1441));
    LocalMux I__6417 (
            .O(N__33724),
            .I(cmd_rdadctmp_9_adj_1441));
    InMux I__6416 (
            .O(N__33717),
            .I(N__33714));
    LocalMux I__6415 (
            .O(N__33714),
            .I(N__33710));
    InMux I__6414 (
            .O(N__33713),
            .I(N__33706));
    Span4Mux_v I__6413 (
            .O(N__33710),
            .I(N__33703));
    CascadeMux I__6412 (
            .O(N__33709),
            .I(N__33700));
    LocalMux I__6411 (
            .O(N__33706),
            .I(N__33697));
    Span4Mux_h I__6410 (
            .O(N__33703),
            .I(N__33694));
    InMux I__6409 (
            .O(N__33700),
            .I(N__33691));
    Span4Mux_v I__6408 (
            .O(N__33697),
            .I(N__33686));
    Span4Mux_h I__6407 (
            .O(N__33694),
            .I(N__33686));
    LocalMux I__6406 (
            .O(N__33691),
            .I(buf_adcdata_vac_1));
    Odrv4 I__6405 (
            .O(N__33686),
            .I(buf_adcdata_vac_1));
    InMux I__6404 (
            .O(N__33681),
            .I(N__33667));
    InMux I__6403 (
            .O(N__33680),
            .I(N__33664));
    CascadeMux I__6402 (
            .O(N__33679),
            .I(N__33659));
    InMux I__6401 (
            .O(N__33678),
            .I(N__33652));
    InMux I__6400 (
            .O(N__33677),
            .I(N__33652));
    InMux I__6399 (
            .O(N__33676),
            .I(N__33644));
    InMux I__6398 (
            .O(N__33675),
            .I(N__33641));
    CascadeMux I__6397 (
            .O(N__33674),
            .I(N__33638));
    InMux I__6396 (
            .O(N__33673),
            .I(N__33631));
    InMux I__6395 (
            .O(N__33672),
            .I(N__33631));
    InMux I__6394 (
            .O(N__33671),
            .I(N__33631));
    InMux I__6393 (
            .O(N__33670),
            .I(N__33628));
    LocalMux I__6392 (
            .O(N__33667),
            .I(N__33625));
    LocalMux I__6391 (
            .O(N__33664),
            .I(N__33622));
    InMux I__6390 (
            .O(N__33663),
            .I(N__33615));
    InMux I__6389 (
            .O(N__33662),
            .I(N__33615));
    InMux I__6388 (
            .O(N__33659),
            .I(N__33610));
    InMux I__6387 (
            .O(N__33658),
            .I(N__33610));
    InMux I__6386 (
            .O(N__33657),
            .I(N__33607));
    LocalMux I__6385 (
            .O(N__33652),
            .I(N__33604));
    InMux I__6384 (
            .O(N__33651),
            .I(N__33598));
    InMux I__6383 (
            .O(N__33650),
            .I(N__33598));
    InMux I__6382 (
            .O(N__33649),
            .I(N__33591));
    InMux I__6381 (
            .O(N__33648),
            .I(N__33591));
    InMux I__6380 (
            .O(N__33647),
            .I(N__33591));
    LocalMux I__6379 (
            .O(N__33644),
            .I(N__33588));
    LocalMux I__6378 (
            .O(N__33641),
            .I(N__33585));
    InMux I__6377 (
            .O(N__33638),
            .I(N__33582));
    LocalMux I__6376 (
            .O(N__33631),
            .I(N__33579));
    LocalMux I__6375 (
            .O(N__33628),
            .I(N__33576));
    Span4Mux_h I__6374 (
            .O(N__33625),
            .I(N__33571));
    Span4Mux_h I__6373 (
            .O(N__33622),
            .I(N__33571));
    InMux I__6372 (
            .O(N__33621),
            .I(N__33566));
    InMux I__6371 (
            .O(N__33620),
            .I(N__33566));
    LocalMux I__6370 (
            .O(N__33615),
            .I(N__33563));
    LocalMux I__6369 (
            .O(N__33610),
            .I(N__33556));
    LocalMux I__6368 (
            .O(N__33607),
            .I(N__33556));
    Span4Mux_h I__6367 (
            .O(N__33604),
            .I(N__33556));
    InMux I__6366 (
            .O(N__33603),
            .I(N__33553));
    LocalMux I__6365 (
            .O(N__33598),
            .I(N__33544));
    LocalMux I__6364 (
            .O(N__33591),
            .I(N__33544));
    Span4Mux_h I__6363 (
            .O(N__33588),
            .I(N__33544));
    Span4Mux_h I__6362 (
            .O(N__33585),
            .I(N__33544));
    LocalMux I__6361 (
            .O(N__33582),
            .I(N__33535));
    Span4Mux_v I__6360 (
            .O(N__33579),
            .I(N__33535));
    Span4Mux_h I__6359 (
            .O(N__33576),
            .I(N__33535));
    Span4Mux_v I__6358 (
            .O(N__33571),
            .I(N__33535));
    LocalMux I__6357 (
            .O(N__33566),
            .I(N__33530));
    Span4Mux_h I__6356 (
            .O(N__33563),
            .I(N__33530));
    Span4Mux_h I__6355 (
            .O(N__33556),
            .I(N__33527));
    LocalMux I__6354 (
            .O(N__33553),
            .I(N__33522));
    Span4Mux_v I__6353 (
            .O(N__33544),
            .I(N__33522));
    Span4Mux_v I__6352 (
            .O(N__33535),
            .I(N__33519));
    Span4Mux_v I__6351 (
            .O(N__33530),
            .I(N__33514));
    Span4Mux_h I__6350 (
            .O(N__33527),
            .I(N__33514));
    Odrv4 I__6349 (
            .O(N__33522),
            .I(n20853));
    Odrv4 I__6348 (
            .O(N__33519),
            .I(n20853));
    Odrv4 I__6347 (
            .O(N__33514),
            .I(n20853));
    CascadeMux I__6346 (
            .O(N__33507),
            .I(N__33498));
    CascadeMux I__6345 (
            .O(N__33506),
            .I(N__33495));
    InMux I__6344 (
            .O(N__33505),
            .I(N__33466));
    InMux I__6343 (
            .O(N__33504),
            .I(N__33466));
    InMux I__6342 (
            .O(N__33503),
            .I(N__33466));
    InMux I__6341 (
            .O(N__33502),
            .I(N__33466));
    InMux I__6340 (
            .O(N__33501),
            .I(N__33463));
    InMux I__6339 (
            .O(N__33498),
            .I(N__33460));
    InMux I__6338 (
            .O(N__33495),
            .I(N__33451));
    InMux I__6337 (
            .O(N__33494),
            .I(N__33451));
    InMux I__6336 (
            .O(N__33493),
            .I(N__33439));
    InMux I__6335 (
            .O(N__33492),
            .I(N__33439));
    InMux I__6334 (
            .O(N__33491),
            .I(N__33439));
    InMux I__6333 (
            .O(N__33490),
            .I(N__33439));
    InMux I__6332 (
            .O(N__33489),
            .I(N__33439));
    InMux I__6331 (
            .O(N__33488),
            .I(N__33432));
    InMux I__6330 (
            .O(N__33487),
            .I(N__33432));
    InMux I__6329 (
            .O(N__33486),
            .I(N__33432));
    InMux I__6328 (
            .O(N__33485),
            .I(N__33421));
    InMux I__6327 (
            .O(N__33484),
            .I(N__33421));
    InMux I__6326 (
            .O(N__33483),
            .I(N__33421));
    InMux I__6325 (
            .O(N__33482),
            .I(N__33421));
    InMux I__6324 (
            .O(N__33481),
            .I(N__33421));
    InMux I__6323 (
            .O(N__33480),
            .I(N__33410));
    InMux I__6322 (
            .O(N__33479),
            .I(N__33410));
    InMux I__6321 (
            .O(N__33478),
            .I(N__33410));
    InMux I__6320 (
            .O(N__33477),
            .I(N__33410));
    InMux I__6319 (
            .O(N__33476),
            .I(N__33410));
    InMux I__6318 (
            .O(N__33475),
            .I(N__33407));
    LocalMux I__6317 (
            .O(N__33466),
            .I(N__33404));
    LocalMux I__6316 (
            .O(N__33463),
            .I(N__33399));
    LocalMux I__6315 (
            .O(N__33460),
            .I(N__33399));
    InMux I__6314 (
            .O(N__33459),
            .I(N__33394));
    InMux I__6313 (
            .O(N__33458),
            .I(N__33394));
    CascadeMux I__6312 (
            .O(N__33457),
            .I(N__33391));
    InMux I__6311 (
            .O(N__33456),
            .I(N__33384));
    LocalMux I__6310 (
            .O(N__33451),
            .I(N__33381));
    InMux I__6309 (
            .O(N__33450),
            .I(N__33370));
    LocalMux I__6308 (
            .O(N__33439),
            .I(N__33367));
    LocalMux I__6307 (
            .O(N__33432),
            .I(N__33360));
    LocalMux I__6306 (
            .O(N__33421),
            .I(N__33360));
    LocalMux I__6305 (
            .O(N__33410),
            .I(N__33360));
    LocalMux I__6304 (
            .O(N__33407),
            .I(N__33357));
    Span4Mux_h I__6303 (
            .O(N__33404),
            .I(N__33354));
    Span4Mux_v I__6302 (
            .O(N__33399),
            .I(N__33351));
    LocalMux I__6301 (
            .O(N__33394),
            .I(N__33348));
    InMux I__6300 (
            .O(N__33391),
            .I(N__33340));
    InMux I__6299 (
            .O(N__33390),
            .I(N__33335));
    InMux I__6298 (
            .O(N__33389),
            .I(N__33335));
    InMux I__6297 (
            .O(N__33388),
            .I(N__33332));
    InMux I__6296 (
            .O(N__33387),
            .I(N__33329));
    LocalMux I__6295 (
            .O(N__33384),
            .I(N__33324));
    Span4Mux_v I__6294 (
            .O(N__33381),
            .I(N__33324));
    InMux I__6293 (
            .O(N__33380),
            .I(N__33313));
    InMux I__6292 (
            .O(N__33379),
            .I(N__33313));
    InMux I__6291 (
            .O(N__33378),
            .I(N__33313));
    InMux I__6290 (
            .O(N__33377),
            .I(N__33313));
    InMux I__6289 (
            .O(N__33376),
            .I(N__33313));
    CascadeMux I__6288 (
            .O(N__33375),
            .I(N__33310));
    InMux I__6287 (
            .O(N__33374),
            .I(N__33301));
    InMux I__6286 (
            .O(N__33373),
            .I(N__33301));
    LocalMux I__6285 (
            .O(N__33370),
            .I(N__33292));
    Span4Mux_h I__6284 (
            .O(N__33367),
            .I(N__33292));
    Span4Mux_h I__6283 (
            .O(N__33360),
            .I(N__33292));
    Span4Mux_v I__6282 (
            .O(N__33357),
            .I(N__33292));
    Span4Mux_v I__6281 (
            .O(N__33354),
            .I(N__33285));
    Span4Mux_v I__6280 (
            .O(N__33351),
            .I(N__33285));
    Span4Mux_h I__6279 (
            .O(N__33348),
            .I(N__33285));
    InMux I__6278 (
            .O(N__33347),
            .I(N__33278));
    InMux I__6277 (
            .O(N__33346),
            .I(N__33278));
    InMux I__6276 (
            .O(N__33345),
            .I(N__33278));
    InMux I__6275 (
            .O(N__33344),
            .I(N__33275));
    CascadeMux I__6274 (
            .O(N__33343),
            .I(N__33269));
    LocalMux I__6273 (
            .O(N__33340),
            .I(N__33261));
    LocalMux I__6272 (
            .O(N__33335),
            .I(N__33254));
    LocalMux I__6271 (
            .O(N__33332),
            .I(N__33254));
    LocalMux I__6270 (
            .O(N__33329),
            .I(N__33251));
    Span4Mux_h I__6269 (
            .O(N__33324),
            .I(N__33246));
    LocalMux I__6268 (
            .O(N__33313),
            .I(N__33246));
    InMux I__6267 (
            .O(N__33310),
            .I(N__33234));
    InMux I__6266 (
            .O(N__33309),
            .I(N__33234));
    InMux I__6265 (
            .O(N__33308),
            .I(N__33234));
    InMux I__6264 (
            .O(N__33307),
            .I(N__33234));
    InMux I__6263 (
            .O(N__33306),
            .I(N__33234));
    LocalMux I__6262 (
            .O(N__33301),
            .I(N__33227));
    Span4Mux_v I__6261 (
            .O(N__33292),
            .I(N__33227));
    Span4Mux_h I__6260 (
            .O(N__33285),
            .I(N__33227));
    LocalMux I__6259 (
            .O(N__33278),
            .I(N__33222));
    LocalMux I__6258 (
            .O(N__33275),
            .I(N__33222));
    InMux I__6257 (
            .O(N__33274),
            .I(N__33213));
    InMux I__6256 (
            .O(N__33273),
            .I(N__33213));
    InMux I__6255 (
            .O(N__33272),
            .I(N__33210));
    InMux I__6254 (
            .O(N__33269),
            .I(N__33207));
    InMux I__6253 (
            .O(N__33268),
            .I(N__33202));
    InMux I__6252 (
            .O(N__33267),
            .I(N__33202));
    InMux I__6251 (
            .O(N__33266),
            .I(N__33195));
    InMux I__6250 (
            .O(N__33265),
            .I(N__33195));
    InMux I__6249 (
            .O(N__33264),
            .I(N__33195));
    Span4Mux_h I__6248 (
            .O(N__33261),
            .I(N__33192));
    InMux I__6247 (
            .O(N__33260),
            .I(N__33189));
    InMux I__6246 (
            .O(N__33259),
            .I(N__33186));
    Span12Mux_v I__6245 (
            .O(N__33254),
            .I(N__33183));
    Span4Mux_h I__6244 (
            .O(N__33251),
            .I(N__33178));
    Span4Mux_v I__6243 (
            .O(N__33246),
            .I(N__33178));
    InMux I__6242 (
            .O(N__33245),
            .I(N__33175));
    LocalMux I__6241 (
            .O(N__33234),
            .I(N__33168));
    Sp12to4 I__6240 (
            .O(N__33227),
            .I(N__33168));
    Span12Mux_h I__6239 (
            .O(N__33222),
            .I(N__33168));
    InMux I__6238 (
            .O(N__33221),
            .I(N__33161));
    InMux I__6237 (
            .O(N__33220),
            .I(N__33161));
    InMux I__6236 (
            .O(N__33219),
            .I(N__33161));
    InMux I__6235 (
            .O(N__33218),
            .I(N__33158));
    LocalMux I__6234 (
            .O(N__33213),
            .I(adc_state_0_adj_1418));
    LocalMux I__6233 (
            .O(N__33210),
            .I(adc_state_0_adj_1418));
    LocalMux I__6232 (
            .O(N__33207),
            .I(adc_state_0_adj_1418));
    LocalMux I__6231 (
            .O(N__33202),
            .I(adc_state_0_adj_1418));
    LocalMux I__6230 (
            .O(N__33195),
            .I(adc_state_0_adj_1418));
    Odrv4 I__6229 (
            .O(N__33192),
            .I(adc_state_0_adj_1418));
    LocalMux I__6228 (
            .O(N__33189),
            .I(adc_state_0_adj_1418));
    LocalMux I__6227 (
            .O(N__33186),
            .I(adc_state_0_adj_1418));
    Odrv12 I__6226 (
            .O(N__33183),
            .I(adc_state_0_adj_1418));
    Odrv4 I__6225 (
            .O(N__33178),
            .I(adc_state_0_adj_1418));
    LocalMux I__6224 (
            .O(N__33175),
            .I(adc_state_0_adj_1418));
    Odrv12 I__6223 (
            .O(N__33168),
            .I(adc_state_0_adj_1418));
    LocalMux I__6222 (
            .O(N__33161),
            .I(adc_state_0_adj_1418));
    LocalMux I__6221 (
            .O(N__33158),
            .I(adc_state_0_adj_1418));
    CascadeMux I__6220 (
            .O(N__33129),
            .I(N__33124));
    InMux I__6219 (
            .O(N__33128),
            .I(N__33121));
    InMux I__6218 (
            .O(N__33127),
            .I(N__33116));
    InMux I__6217 (
            .O(N__33124),
            .I(N__33116));
    LocalMux I__6216 (
            .O(N__33121),
            .I(cmd_rdadctmp_18_adj_1432));
    LocalMux I__6215 (
            .O(N__33116),
            .I(cmd_rdadctmp_18_adj_1432));
    CascadeMux I__6214 (
            .O(N__33111),
            .I(N__33108));
    InMux I__6213 (
            .O(N__33108),
            .I(N__33105));
    LocalMux I__6212 (
            .O(N__33105),
            .I(N__33102));
    Span12Mux_h I__6211 (
            .O(N__33102),
            .I(N__33099));
    Odrv12 I__6210 (
            .O(N__33099),
            .I(n9_adj_1416));
    CascadeMux I__6209 (
            .O(N__33096),
            .I(n31_adj_1613_cascade_));
    CEMux I__6208 (
            .O(N__33093),
            .I(N__33089));
    CEMux I__6207 (
            .O(N__33092),
            .I(N__33086));
    LocalMux I__6206 (
            .O(N__33089),
            .I(N__33083));
    LocalMux I__6205 (
            .O(N__33086),
            .I(N__33080));
    Odrv4 I__6204 (
            .O(N__33083),
            .I(n12085));
    Odrv12 I__6203 (
            .O(N__33080),
            .I(n12085));
    CascadeMux I__6202 (
            .O(N__33075),
            .I(n12085_cascade_));
    SRMux I__6201 (
            .O(N__33072),
            .I(N__33068));
    SRMux I__6200 (
            .O(N__33071),
            .I(N__33065));
    LocalMux I__6199 (
            .O(N__33068),
            .I(N__33062));
    LocalMux I__6198 (
            .O(N__33065),
            .I(N__33059));
    Span4Mux_h I__6197 (
            .O(N__33062),
            .I(N__33056));
    Odrv4 I__6196 (
            .O(N__33059),
            .I(n14764));
    Odrv4 I__6195 (
            .O(N__33056),
            .I(n14764));
    CascadeMux I__6194 (
            .O(N__33051),
            .I(n12228_cascade_));
    InMux I__6193 (
            .O(N__33048),
            .I(N__33044));
    InMux I__6192 (
            .O(N__33047),
            .I(N__33041));
    LocalMux I__6191 (
            .O(N__33044),
            .I(comm_buf_6_7));
    LocalMux I__6190 (
            .O(N__33041),
            .I(comm_buf_6_7));
    InMux I__6189 (
            .O(N__33036),
            .I(N__33033));
    LocalMux I__6188 (
            .O(N__33033),
            .I(n20850));
    InMux I__6187 (
            .O(N__33030),
            .I(N__33027));
    LocalMux I__6186 (
            .O(N__33027),
            .I(n20852));
    InMux I__6185 (
            .O(N__33024),
            .I(N__33021));
    LocalMux I__6184 (
            .O(N__33021),
            .I(comm_buf_2_3));
    CascadeMux I__6183 (
            .O(N__33018),
            .I(n22387_cascade_));
    InMux I__6182 (
            .O(N__33015),
            .I(N__33012));
    LocalMux I__6181 (
            .O(N__33012),
            .I(n21193));
    CascadeMux I__6180 (
            .O(N__33009),
            .I(n22390_cascade_));
    CascadeMux I__6179 (
            .O(N__33006),
            .I(n4_adj_1587_cascade_));
    CascadeMux I__6178 (
            .O(N__33003),
            .I(n21175_cascade_));
    CascadeMux I__6177 (
            .O(N__33000),
            .I(n2358_cascade_));
    CascadeMux I__6176 (
            .O(N__32997),
            .I(n20850_cascade_));
    InMux I__6175 (
            .O(N__32994),
            .I(N__32991));
    LocalMux I__6174 (
            .O(N__32991),
            .I(N__32988));
    Span4Mux_v I__6173 (
            .O(N__32988),
            .I(N__32985));
    Odrv4 I__6172 (
            .O(N__32985),
            .I(n30_adj_1482));
    InMux I__6171 (
            .O(N__32982),
            .I(N__32979));
    LocalMux I__6170 (
            .O(N__32979),
            .I(N__32976));
    Span4Mux_h I__6169 (
            .O(N__32976),
            .I(N__32973));
    Span4Mux_h I__6168 (
            .O(N__32973),
            .I(N__32970));
    Odrv4 I__6167 (
            .O(N__32970),
            .I(n30_adj_1625));
    InMux I__6166 (
            .O(N__32967),
            .I(N__32964));
    LocalMux I__6165 (
            .O(N__32964),
            .I(comm_buf_2_7));
    InMux I__6164 (
            .O(N__32961),
            .I(N__32958));
    LocalMux I__6163 (
            .O(N__32958),
            .I(N__32955));
    Span4Mux_h I__6162 (
            .O(N__32955),
            .I(N__32952));
    Span4Mux_h I__6161 (
            .O(N__32952),
            .I(N__32949));
    Odrv4 I__6160 (
            .O(N__32949),
            .I(n30_adj_1628));
    InMux I__6159 (
            .O(N__32946),
            .I(N__32943));
    LocalMux I__6158 (
            .O(N__32943),
            .I(N__32940));
    Span4Mux_h I__6157 (
            .O(N__32940),
            .I(N__32937));
    Odrv4 I__6156 (
            .O(N__32937),
            .I(n30_adj_1631));
    InMux I__6155 (
            .O(N__32934),
            .I(N__32931));
    LocalMux I__6154 (
            .O(N__32931),
            .I(N__32928));
    Odrv12 I__6153 (
            .O(N__32928),
            .I(n30_adj_1634));
    InMux I__6152 (
            .O(N__32925),
            .I(N__32922));
    LocalMux I__6151 (
            .O(N__32922),
            .I(N__32919));
    Odrv4 I__6150 (
            .O(N__32919),
            .I(n30_adj_1638));
    InMux I__6149 (
            .O(N__32916),
            .I(N__32913));
    LocalMux I__6148 (
            .O(N__32913),
            .I(N__32910));
    Odrv4 I__6147 (
            .O(N__32910),
            .I(n30_adj_1641));
    CascadeMux I__6146 (
            .O(N__32907),
            .I(n4_adj_1594_cascade_));
    InMux I__6145 (
            .O(N__32904),
            .I(N__32901));
    LocalMux I__6144 (
            .O(N__32901),
            .I(\ADC_VDC.n21229 ));
    CEMux I__6143 (
            .O(N__32898),
            .I(N__32895));
    LocalMux I__6142 (
            .O(N__32895),
            .I(N__32892));
    Odrv12 I__6141 (
            .O(N__32892),
            .I(\ADC_VDC.n47 ));
    InMux I__6140 (
            .O(N__32889),
            .I(N__32886));
    LocalMux I__6139 (
            .O(N__32886),
            .I(N__32883));
    Span4Mux_v I__6138 (
            .O(N__32883),
            .I(N__32879));
    InMux I__6137 (
            .O(N__32882),
            .I(N__32876));
    Odrv4 I__6136 (
            .O(N__32879),
            .I(\comm_spi.n14608 ));
    LocalMux I__6135 (
            .O(N__32876),
            .I(\comm_spi.n14608 ));
    CascadeMux I__6134 (
            .O(N__32871),
            .I(N__32868));
    InMux I__6133 (
            .O(N__32868),
            .I(N__32865));
    LocalMux I__6132 (
            .O(N__32865),
            .I(N__32861));
    CascadeMux I__6131 (
            .O(N__32864),
            .I(N__32858));
    Span4Mux_v I__6130 (
            .O(N__32861),
            .I(N__32855));
    InMux I__6129 (
            .O(N__32858),
            .I(N__32852));
    Odrv4 I__6128 (
            .O(N__32855),
            .I(buf_adcdata_vdc_1));
    LocalMux I__6127 (
            .O(N__32852),
            .I(buf_adcdata_vdc_1));
    InMux I__6126 (
            .O(N__32847),
            .I(N__32843));
    InMux I__6125 (
            .O(N__32846),
            .I(N__32839));
    LocalMux I__6124 (
            .O(N__32843),
            .I(N__32836));
    InMux I__6123 (
            .O(N__32842),
            .I(N__32833));
    LocalMux I__6122 (
            .O(N__32839),
            .I(N__32828));
    Span12Mux_s9_h I__6121 (
            .O(N__32836),
            .I(N__32828));
    LocalMux I__6120 (
            .O(N__32833),
            .I(buf_adcdata_iac_1));
    Odrv12 I__6119 (
            .O(N__32828),
            .I(buf_adcdata_iac_1));
    CascadeMux I__6118 (
            .O(N__32823),
            .I(n19_adj_1491_cascade_));
    InMux I__6117 (
            .O(N__32820),
            .I(N__32817));
    LocalMux I__6116 (
            .O(N__32817),
            .I(N__32814));
    Span4Mux_h I__6115 (
            .O(N__32814),
            .I(N__32811));
    Span4Mux_h I__6114 (
            .O(N__32811),
            .I(N__32808));
    Odrv4 I__6113 (
            .O(N__32808),
            .I(buf_data_iac_1));
    CascadeMux I__6112 (
            .O(N__32805),
            .I(n22_adj_1488_cascade_));
    InMux I__6111 (
            .O(N__32802),
            .I(N__32799));
    LocalMux I__6110 (
            .O(N__32799),
            .I(n30_adj_1506));
    InMux I__6109 (
            .O(N__32796),
            .I(N__32793));
    LocalMux I__6108 (
            .O(N__32793),
            .I(comm_buf_2_1));
    CascadeMux I__6107 (
            .O(N__32790),
            .I(n22249_cascade_));
    CascadeMux I__6106 (
            .O(N__32787),
            .I(\ADC_VDC.n77_cascade_ ));
    InMux I__6105 (
            .O(N__32784),
            .I(N__32781));
    LocalMux I__6104 (
            .O(N__32781),
            .I(\ADC_VDC.n12 ));
    InMux I__6103 (
            .O(N__32778),
            .I(N__32775));
    LocalMux I__6102 (
            .O(N__32775),
            .I(\ADC_VDC.n20899 ));
    CascadeMux I__6101 (
            .O(N__32772),
            .I(\ADC_VDC.n72_cascade_ ));
    CascadeMux I__6100 (
            .O(N__32769),
            .I(\ADC_VDC.n31_cascade_ ));
    CascadeMux I__6099 (
            .O(N__32766),
            .I(\ADC_VDC.n22195_cascade_ ));
    CascadeMux I__6098 (
            .O(N__32763),
            .I(\ADC_VDC.n22198_cascade_ ));
    InMux I__6097 (
            .O(N__32760),
            .I(N__32757));
    LocalMux I__6096 (
            .O(N__32757),
            .I(N__32754));
    Span4Mux_h I__6095 (
            .O(N__32754),
            .I(N__32751));
    Span4Mux_h I__6094 (
            .O(N__32751),
            .I(N__32748));
    Odrv4 I__6093 (
            .O(N__32748),
            .I(\ADC_VDC.n18566 ));
    CEMux I__6092 (
            .O(N__32745),
            .I(N__32742));
    LocalMux I__6091 (
            .O(N__32742),
            .I(N__32739));
    Odrv4 I__6090 (
            .O(N__32739),
            .I(\ADC_VDC.n20811 ));
    CascadeMux I__6089 (
            .O(N__32736),
            .I(\ADC_VDC.n6_adj_1399_cascade_ ));
    InMux I__6088 (
            .O(N__32733),
            .I(N__32730));
    LocalMux I__6087 (
            .O(N__32730),
            .I(N__32727));
    Span4Mux_h I__6086 (
            .O(N__32727),
            .I(N__32723));
    InMux I__6085 (
            .O(N__32726),
            .I(N__32720));
    Odrv4 I__6084 (
            .O(N__32723),
            .I(\ADC_VDC.n10536 ));
    LocalMux I__6083 (
            .O(N__32720),
            .I(\ADC_VDC.n10536 ));
    InMux I__6082 (
            .O(N__32715),
            .I(N__32712));
    LocalMux I__6081 (
            .O(N__32712),
            .I(N__32708));
    InMux I__6080 (
            .O(N__32711),
            .I(N__32705));
    Span4Mux_v I__6079 (
            .O(N__32708),
            .I(N__32702));
    LocalMux I__6078 (
            .O(N__32705),
            .I(acadc_skipcnt_13));
    Odrv4 I__6077 (
            .O(N__32702),
            .I(acadc_skipcnt_13));
    InMux I__6076 (
            .O(N__32697),
            .I(n19622));
    InMux I__6075 (
            .O(N__32694),
            .I(N__32690));
    InMux I__6074 (
            .O(N__32693),
            .I(N__32687));
    LocalMux I__6073 (
            .O(N__32690),
            .I(N__32684));
    LocalMux I__6072 (
            .O(N__32687),
            .I(acadc_skipcnt_14));
    Odrv4 I__6071 (
            .O(N__32684),
            .I(acadc_skipcnt_14));
    InMux I__6070 (
            .O(N__32679),
            .I(n19623));
    InMux I__6069 (
            .O(N__32676),
            .I(n19624));
    InMux I__6068 (
            .O(N__32673),
            .I(N__32669));
    InMux I__6067 (
            .O(N__32672),
            .I(N__32666));
    LocalMux I__6066 (
            .O(N__32669),
            .I(N__32663));
    LocalMux I__6065 (
            .O(N__32666),
            .I(acadc_skipcnt_15));
    Odrv12 I__6064 (
            .O(N__32663),
            .I(acadc_skipcnt_15));
    CEMux I__6063 (
            .O(N__32658),
            .I(N__32653));
    CEMux I__6062 (
            .O(N__32657),
            .I(N__32650));
    CEMux I__6061 (
            .O(N__32656),
            .I(N__32647));
    LocalMux I__6060 (
            .O(N__32653),
            .I(N__32643));
    LocalMux I__6059 (
            .O(N__32650),
            .I(N__32638));
    LocalMux I__6058 (
            .O(N__32647),
            .I(N__32638));
    InMux I__6057 (
            .O(N__32646),
            .I(N__32635));
    Span4Mux_v I__6056 (
            .O(N__32643),
            .I(N__32630));
    Span4Mux_v I__6055 (
            .O(N__32638),
            .I(N__32630));
    LocalMux I__6054 (
            .O(N__32635),
            .I(N__32627));
    Odrv4 I__6053 (
            .O(N__32630),
            .I(n11654));
    Odrv4 I__6052 (
            .O(N__32627),
            .I(n11654));
    SRMux I__6051 (
            .O(N__32622),
            .I(N__32619));
    LocalMux I__6050 (
            .O(N__32619),
            .I(N__32615));
    SRMux I__6049 (
            .O(N__32618),
            .I(N__32612));
    Span4Mux_v I__6048 (
            .O(N__32615),
            .I(N__32609));
    LocalMux I__6047 (
            .O(N__32612),
            .I(N__32606));
    Span4Mux_h I__6046 (
            .O(N__32609),
            .I(N__32601));
    Span4Mux_v I__6045 (
            .O(N__32606),
            .I(N__32601));
    Odrv4 I__6044 (
            .O(N__32601),
            .I(n14671));
    CEMux I__6043 (
            .O(N__32598),
            .I(N__32595));
    LocalMux I__6042 (
            .O(N__32595),
            .I(N__32592));
    Odrv4 I__6041 (
            .O(N__32592),
            .I(\ADC_VDC.n17 ));
    SRMux I__6040 (
            .O(N__32589),
            .I(N__32586));
    LocalMux I__6039 (
            .O(N__32586),
            .I(N__32583));
    Span4Mux_h I__6038 (
            .O(N__32583),
            .I(N__32580));
    Odrv4 I__6037 (
            .O(N__32580),
            .I(\ADC_VDC.n4 ));
    InMux I__6036 (
            .O(N__32577),
            .I(N__32574));
    LocalMux I__6035 (
            .O(N__32574),
            .I(\ADC_VDC.n7_adj_1398 ));
    CascadeMux I__6034 (
            .O(N__32571),
            .I(\ADC_VDC.n7_adj_1398_cascade_ ));
    InMux I__6033 (
            .O(N__32568),
            .I(N__32564));
    InMux I__6032 (
            .O(N__32567),
            .I(N__32561));
    LocalMux I__6031 (
            .O(N__32564),
            .I(\ADC_VDC.n77 ));
    LocalMux I__6030 (
            .O(N__32561),
            .I(\ADC_VDC.n77 ));
    CascadeMux I__6029 (
            .O(N__32556),
            .I(N__32552));
    InMux I__6028 (
            .O(N__32555),
            .I(N__32549));
    InMux I__6027 (
            .O(N__32552),
            .I(N__32546));
    LocalMux I__6026 (
            .O(N__32549),
            .I(acadc_skipcnt_4));
    LocalMux I__6025 (
            .O(N__32546),
            .I(acadc_skipcnt_4));
    InMux I__6024 (
            .O(N__32541),
            .I(n19613));
    InMux I__6023 (
            .O(N__32538),
            .I(N__32534));
    InMux I__6022 (
            .O(N__32537),
            .I(N__32531));
    LocalMux I__6021 (
            .O(N__32534),
            .I(N__32528));
    LocalMux I__6020 (
            .O(N__32531),
            .I(acadc_skipcnt_5));
    Odrv4 I__6019 (
            .O(N__32528),
            .I(acadc_skipcnt_5));
    InMux I__6018 (
            .O(N__32523),
            .I(n19614));
    InMux I__6017 (
            .O(N__32520),
            .I(n19615));
    InMux I__6016 (
            .O(N__32517),
            .I(n19616));
    InMux I__6015 (
            .O(N__32514),
            .I(N__32510));
    InMux I__6014 (
            .O(N__32513),
            .I(N__32507));
    LocalMux I__6013 (
            .O(N__32510),
            .I(N__32504));
    LocalMux I__6012 (
            .O(N__32507),
            .I(acadc_skipcnt_8));
    Odrv4 I__6011 (
            .O(N__32504),
            .I(acadc_skipcnt_8));
    InMux I__6010 (
            .O(N__32499),
            .I(n19617));
    InMux I__6009 (
            .O(N__32496),
            .I(N__32492));
    InMux I__6008 (
            .O(N__32495),
            .I(N__32489));
    LocalMux I__6007 (
            .O(N__32492),
            .I(N__32486));
    LocalMux I__6006 (
            .O(N__32489),
            .I(acadc_skipcnt_9));
    Odrv4 I__6005 (
            .O(N__32486),
            .I(acadc_skipcnt_9));
    InMux I__6004 (
            .O(N__32481),
            .I(bfn_12_20_0_));
    InMux I__6003 (
            .O(N__32478),
            .I(N__32475));
    LocalMux I__6002 (
            .O(N__32475),
            .I(N__32471));
    InMux I__6001 (
            .O(N__32474),
            .I(N__32468));
    Span4Mux_h I__6000 (
            .O(N__32471),
            .I(N__32465));
    LocalMux I__5999 (
            .O(N__32468),
            .I(acadc_skipcnt_10));
    Odrv4 I__5998 (
            .O(N__32465),
            .I(acadc_skipcnt_10));
    InMux I__5997 (
            .O(N__32460),
            .I(n19619));
    InMux I__5996 (
            .O(N__32457),
            .I(N__32453));
    InMux I__5995 (
            .O(N__32456),
            .I(N__32450));
    LocalMux I__5994 (
            .O(N__32453),
            .I(N__32447));
    LocalMux I__5993 (
            .O(N__32450),
            .I(acadc_skipcnt_11));
    Odrv4 I__5992 (
            .O(N__32447),
            .I(acadc_skipcnt_11));
    InMux I__5991 (
            .O(N__32442),
            .I(n19620));
    InMux I__5990 (
            .O(N__32439),
            .I(N__32436));
    LocalMux I__5989 (
            .O(N__32436),
            .I(N__32432));
    InMux I__5988 (
            .O(N__32435),
            .I(N__32429));
    Span4Mux_h I__5987 (
            .O(N__32432),
            .I(N__32426));
    LocalMux I__5986 (
            .O(N__32429),
            .I(acadc_skipcnt_12));
    Odrv4 I__5985 (
            .O(N__32426),
            .I(acadc_skipcnt_12));
    InMux I__5984 (
            .O(N__32421),
            .I(n19621));
    InMux I__5983 (
            .O(N__32418),
            .I(N__32414));
    InMux I__5982 (
            .O(N__32417),
            .I(N__32411));
    LocalMux I__5981 (
            .O(N__32414),
            .I(acadc_skipcnt_1));
    LocalMux I__5980 (
            .O(N__32411),
            .I(acadc_skipcnt_1));
    InMux I__5979 (
            .O(N__32406),
            .I(bfn_12_19_0_));
    InMux I__5978 (
            .O(N__32403),
            .I(n19611));
    InMux I__5977 (
            .O(N__32400),
            .I(N__32396));
    InMux I__5976 (
            .O(N__32399),
            .I(N__32393));
    LocalMux I__5975 (
            .O(N__32396),
            .I(N__32390));
    LocalMux I__5974 (
            .O(N__32393),
            .I(acadc_skipcnt_3));
    Odrv4 I__5973 (
            .O(N__32390),
            .I(acadc_skipcnt_3));
    InMux I__5972 (
            .O(N__32385),
            .I(n19612));
    InMux I__5971 (
            .O(N__32382),
            .I(N__32379));
    LocalMux I__5970 (
            .O(N__32379),
            .I(n23_adj_1501));
    InMux I__5969 (
            .O(N__32376),
            .I(N__32373));
    LocalMux I__5968 (
            .O(N__32373),
            .I(n24_adj_1642));
    InMux I__5967 (
            .O(N__32370),
            .I(N__32367));
    LocalMux I__5966 (
            .O(N__32367),
            .I(N__32364));
    Span4Mux_h I__5965 (
            .O(N__32364),
            .I(N__32361));
    Span4Mux_v I__5964 (
            .O(N__32361),
            .I(N__32356));
    InMux I__5963 (
            .O(N__32360),
            .I(N__32351));
    InMux I__5962 (
            .O(N__32359),
            .I(N__32351));
    Odrv4 I__5961 (
            .O(N__32356),
            .I(acadc_skipCount_15));
    LocalMux I__5960 (
            .O(N__32351),
            .I(acadc_skipCount_15));
    SRMux I__5959 (
            .O(N__32346),
            .I(N__32343));
    LocalMux I__5958 (
            .O(N__32343),
            .I(N__32340));
    Span4Mux_v I__5957 (
            .O(N__32340),
            .I(N__32337));
    Span4Mux_v I__5956 (
            .O(N__32337),
            .I(N__32334));
    Odrv4 I__5955 (
            .O(N__32334),
            .I(n21037));
    InMux I__5954 (
            .O(N__32331),
            .I(N__32328));
    LocalMux I__5953 (
            .O(N__32328),
            .I(\SIG_DDS.tmp_buf_6 ));
    InMux I__5952 (
            .O(N__32325),
            .I(N__32322));
    LocalMux I__5951 (
            .O(N__32322),
            .I(N__32318));
    InMux I__5950 (
            .O(N__32321),
            .I(N__32314));
    Span4Mux_v I__5949 (
            .O(N__32318),
            .I(N__32311));
    InMux I__5948 (
            .O(N__32317),
            .I(N__32308));
    LocalMux I__5947 (
            .O(N__32314),
            .I(buf_dds0_7));
    Odrv4 I__5946 (
            .O(N__32311),
            .I(buf_dds0_7));
    LocalMux I__5945 (
            .O(N__32308),
            .I(buf_dds0_7));
    InMux I__5944 (
            .O(N__32301),
            .I(N__32298));
    LocalMux I__5943 (
            .O(N__32298),
            .I(\SIG_DDS.tmp_buf_7 ));
    InMux I__5942 (
            .O(N__32295),
            .I(N__32291));
    InMux I__5941 (
            .O(N__32294),
            .I(N__32287));
    LocalMux I__5940 (
            .O(N__32291),
            .I(N__32284));
    InMux I__5939 (
            .O(N__32290),
            .I(N__32281));
    LocalMux I__5938 (
            .O(N__32287),
            .I(acadc_skipCount_12));
    Odrv4 I__5937 (
            .O(N__32284),
            .I(acadc_skipCount_12));
    LocalMux I__5936 (
            .O(N__32281),
            .I(acadc_skipCount_12));
    CascadeMux I__5935 (
            .O(N__32274),
            .I(N__32269));
    CascadeMux I__5934 (
            .O(N__32273),
            .I(N__32266));
    InMux I__5933 (
            .O(N__32272),
            .I(N__32263));
    InMux I__5932 (
            .O(N__32269),
            .I(N__32260));
    InMux I__5931 (
            .O(N__32266),
            .I(N__32257));
    LocalMux I__5930 (
            .O(N__32263),
            .I(N__32252));
    LocalMux I__5929 (
            .O(N__32260),
            .I(N__32252));
    LocalMux I__5928 (
            .O(N__32257),
            .I(acadc_skipCount_10));
    Odrv4 I__5927 (
            .O(N__32252),
            .I(acadc_skipCount_10));
    InMux I__5926 (
            .O(N__32247),
            .I(N__32244));
    LocalMux I__5925 (
            .O(N__32244),
            .I(N__32240));
    InMux I__5924 (
            .O(N__32243),
            .I(N__32236));
    Span4Mux_h I__5923 (
            .O(N__32240),
            .I(N__32233));
    InMux I__5922 (
            .O(N__32239),
            .I(N__32230));
    LocalMux I__5921 (
            .O(N__32236),
            .I(acadc_skipCount_13));
    Odrv4 I__5920 (
            .O(N__32233),
            .I(acadc_skipCount_13));
    LocalMux I__5919 (
            .O(N__32230),
            .I(acadc_skipCount_13));
    InMux I__5918 (
            .O(N__32223),
            .I(N__32220));
    LocalMux I__5917 (
            .O(N__32220),
            .I(n20));
    InMux I__5916 (
            .O(N__32217),
            .I(N__32214));
    LocalMux I__5915 (
            .O(N__32214),
            .I(N__32208));
    InMux I__5914 (
            .O(N__32213),
            .I(N__32201));
    InMux I__5913 (
            .O(N__32212),
            .I(N__32201));
    InMux I__5912 (
            .O(N__32211),
            .I(N__32198));
    Span4Mux_h I__5911 (
            .O(N__32208),
            .I(N__32195));
    InMux I__5910 (
            .O(N__32207),
            .I(N__32190));
    InMux I__5909 (
            .O(N__32206),
            .I(N__32190));
    LocalMux I__5908 (
            .O(N__32201),
            .I(N__32187));
    LocalMux I__5907 (
            .O(N__32198),
            .I(acadc_dtrig_v));
    Odrv4 I__5906 (
            .O(N__32195),
            .I(acadc_dtrig_v));
    LocalMux I__5905 (
            .O(N__32190),
            .I(acadc_dtrig_v));
    Odrv4 I__5904 (
            .O(N__32187),
            .I(acadc_dtrig_v));
    InMux I__5903 (
            .O(N__32178),
            .I(N__32170));
    InMux I__5902 (
            .O(N__32177),
            .I(N__32165));
    InMux I__5901 (
            .O(N__32176),
            .I(N__32165));
    InMux I__5900 (
            .O(N__32175),
            .I(N__32158));
    InMux I__5899 (
            .O(N__32174),
            .I(N__32158));
    InMux I__5898 (
            .O(N__32173),
            .I(N__32158));
    LocalMux I__5897 (
            .O(N__32170),
            .I(acadc_dtrig_i));
    LocalMux I__5896 (
            .O(N__32165),
            .I(acadc_dtrig_i));
    LocalMux I__5895 (
            .O(N__32158),
            .I(acadc_dtrig_i));
    InMux I__5894 (
            .O(N__32151),
            .I(N__32148));
    LocalMux I__5893 (
            .O(N__32148),
            .I(n4_adj_1546));
    InMux I__5892 (
            .O(N__32145),
            .I(N__32141));
    InMux I__5891 (
            .O(N__32144),
            .I(N__32138));
    LocalMux I__5890 (
            .O(N__32141),
            .I(N__32135));
    LocalMux I__5889 (
            .O(N__32138),
            .I(N__32131));
    Span4Mux_h I__5888 (
            .O(N__32135),
            .I(N__32128));
    InMux I__5887 (
            .O(N__32134),
            .I(N__32125));
    Span4Mux_h I__5886 (
            .O(N__32131),
            .I(N__32122));
    Span4Mux_v I__5885 (
            .O(N__32128),
            .I(N__32119));
    LocalMux I__5884 (
            .O(N__32125),
            .I(buf_dds0_1));
    Odrv4 I__5883 (
            .O(N__32122),
            .I(buf_dds0_1));
    Odrv4 I__5882 (
            .O(N__32119),
            .I(buf_dds0_1));
    InMux I__5881 (
            .O(N__32112),
            .I(N__32109));
    LocalMux I__5880 (
            .O(N__32109),
            .I(\SIG_DDS.tmp_buf_0 ));
    InMux I__5879 (
            .O(N__32106),
            .I(N__32103));
    LocalMux I__5878 (
            .O(N__32103),
            .I(\SIG_DDS.tmp_buf_1 ));
    InMux I__5877 (
            .O(N__32100),
            .I(N__32097));
    LocalMux I__5876 (
            .O(N__32097),
            .I(\SIG_DDS.tmp_buf_2 ));
    InMux I__5875 (
            .O(N__32094),
            .I(N__32091));
    LocalMux I__5874 (
            .O(N__32091),
            .I(\SIG_DDS.tmp_buf_14 ));
    CascadeMux I__5873 (
            .O(N__32088),
            .I(N__32085));
    InMux I__5872 (
            .O(N__32085),
            .I(N__32082));
    LocalMux I__5871 (
            .O(N__32082),
            .I(N__32079));
    Span4Mux_h I__5870 (
            .O(N__32079),
            .I(N__32075));
    InMux I__5869 (
            .O(N__32078),
            .I(N__32071));
    Span4Mux_v I__5868 (
            .O(N__32075),
            .I(N__32068));
    InMux I__5867 (
            .O(N__32074),
            .I(N__32065));
    LocalMux I__5866 (
            .O(N__32071),
            .I(buf_dds0_15));
    Odrv4 I__5865 (
            .O(N__32068),
            .I(buf_dds0_15));
    LocalMux I__5864 (
            .O(N__32065),
            .I(buf_dds0_15));
    InMux I__5863 (
            .O(N__32058),
            .I(N__32055));
    LocalMux I__5862 (
            .O(N__32055),
            .I(\SIG_DDS.tmp_buf_3 ));
    CascadeMux I__5861 (
            .O(N__32052),
            .I(N__32049));
    InMux I__5860 (
            .O(N__32049),
            .I(N__32046));
    LocalMux I__5859 (
            .O(N__32046),
            .I(\SIG_DDS.tmp_buf_4 ));
    CascadeMux I__5858 (
            .O(N__32043),
            .I(N__32040));
    InMux I__5857 (
            .O(N__32040),
            .I(N__32037));
    LocalMux I__5856 (
            .O(N__32037),
            .I(N__32032));
    InMux I__5855 (
            .O(N__32036),
            .I(N__32029));
    InMux I__5854 (
            .O(N__32035),
            .I(N__32026));
    Span12Mux_h I__5853 (
            .O(N__32032),
            .I(N__32023));
    LocalMux I__5852 (
            .O(N__32029),
            .I(N__32020));
    LocalMux I__5851 (
            .O(N__32026),
            .I(buf_dds0_8));
    Odrv12 I__5850 (
            .O(N__32023),
            .I(buf_dds0_8));
    Odrv4 I__5849 (
            .O(N__32020),
            .I(buf_dds0_8));
    CascadeMux I__5848 (
            .O(N__32013),
            .I(N__32010));
    InMux I__5847 (
            .O(N__32010),
            .I(N__32007));
    LocalMux I__5846 (
            .O(N__32007),
            .I(N__32004));
    Odrv4 I__5845 (
            .O(N__32004),
            .I(\SIG_DDS.tmp_buf_8 ));
    CascadeMux I__5844 (
            .O(N__32001),
            .I(N__31998));
    InMux I__5843 (
            .O(N__31998),
            .I(N__31995));
    LocalMux I__5842 (
            .O(N__31995),
            .I(N__31990));
    InMux I__5841 (
            .O(N__31994),
            .I(N__31987));
    CascadeMux I__5840 (
            .O(N__31993),
            .I(N__31984));
    Span12Mux_v I__5839 (
            .O(N__31990),
            .I(N__31981));
    LocalMux I__5838 (
            .O(N__31987),
            .I(N__31978));
    InMux I__5837 (
            .O(N__31984),
            .I(N__31975));
    Odrv12 I__5836 (
            .O(N__31981),
            .I(cmd_rdadctmp_19));
    Odrv4 I__5835 (
            .O(N__31978),
            .I(cmd_rdadctmp_19));
    LocalMux I__5834 (
            .O(N__31975),
            .I(cmd_rdadctmp_19));
    CascadeMux I__5833 (
            .O(N__31968),
            .I(N__31965));
    InMux I__5832 (
            .O(N__31965),
            .I(N__31960));
    CascadeMux I__5831 (
            .O(N__31964),
            .I(N__31957));
    InMux I__5830 (
            .O(N__31963),
            .I(N__31954));
    LocalMux I__5829 (
            .O(N__31960),
            .I(N__31951));
    InMux I__5828 (
            .O(N__31957),
            .I(N__31948));
    LocalMux I__5827 (
            .O(N__31954),
            .I(N__31943));
    Span4Mux_h I__5826 (
            .O(N__31951),
            .I(N__31943));
    LocalMux I__5825 (
            .O(N__31948),
            .I(cmd_rdadctmp_25));
    Odrv4 I__5824 (
            .O(N__31943),
            .I(cmd_rdadctmp_25));
    InMux I__5823 (
            .O(N__31938),
            .I(N__31934));
    InMux I__5822 (
            .O(N__31937),
            .I(N__31930));
    LocalMux I__5821 (
            .O(N__31934),
            .I(N__31927));
    CascadeMux I__5820 (
            .O(N__31933),
            .I(N__31924));
    LocalMux I__5819 (
            .O(N__31930),
            .I(N__31921));
    Span12Mux_h I__5818 (
            .O(N__31927),
            .I(N__31918));
    InMux I__5817 (
            .O(N__31924),
            .I(N__31915));
    Span4Mux_h I__5816 (
            .O(N__31921),
            .I(N__31912));
    Span12Mux_v I__5815 (
            .O(N__31918),
            .I(N__31909));
    LocalMux I__5814 (
            .O(N__31915),
            .I(buf_adcdata_iac_22));
    Odrv4 I__5813 (
            .O(N__31912),
            .I(buf_adcdata_iac_22));
    Odrv12 I__5812 (
            .O(N__31909),
            .I(buf_adcdata_iac_22));
    IoInMux I__5811 (
            .O(N__31902),
            .I(N__31899));
    LocalMux I__5810 (
            .O(N__31899),
            .I(N__31896));
    Span4Mux_s2_h I__5809 (
            .O(N__31896),
            .I(N__31892));
    InMux I__5808 (
            .O(N__31895),
            .I(N__31889));
    Sp12to4 I__5807 (
            .O(N__31892),
            .I(N__31886));
    LocalMux I__5806 (
            .O(N__31889),
            .I(N__31882));
    Span12Mux_v I__5805 (
            .O(N__31886),
            .I(N__31879));
    InMux I__5804 (
            .O(N__31885),
            .I(N__31876));
    Span4Mux_h I__5803 (
            .O(N__31882),
            .I(N__31873));
    Odrv12 I__5802 (
            .O(N__31879),
            .I(VAC_FLT0));
    LocalMux I__5801 (
            .O(N__31876),
            .I(VAC_FLT0));
    Odrv4 I__5800 (
            .O(N__31873),
            .I(VAC_FLT0));
    IoInMux I__5799 (
            .O(N__31866),
            .I(N__31863));
    LocalMux I__5798 (
            .O(N__31863),
            .I(N__31860));
    Span4Mux_s0_h I__5797 (
            .O(N__31860),
            .I(N__31856));
    CascadeMux I__5796 (
            .O(N__31859),
            .I(N__31853));
    Sp12to4 I__5795 (
            .O(N__31856),
            .I(N__31850));
    InMux I__5794 (
            .O(N__31853),
            .I(N__31846));
    Span12Mux_v I__5793 (
            .O(N__31850),
            .I(N__31843));
    CascadeMux I__5792 (
            .O(N__31849),
            .I(N__31840));
    LocalMux I__5791 (
            .O(N__31846),
            .I(N__31837));
    Span12Mux_h I__5790 (
            .O(N__31843),
            .I(N__31834));
    InMux I__5789 (
            .O(N__31840),
            .I(N__31831));
    Span4Mux_v I__5788 (
            .O(N__31837),
            .I(N__31828));
    Odrv12 I__5787 (
            .O(N__31834),
            .I(VDC_RNG0));
    LocalMux I__5786 (
            .O(N__31831),
            .I(VDC_RNG0));
    Odrv4 I__5785 (
            .O(N__31828),
            .I(VDC_RNG0));
    CascadeMux I__5784 (
            .O(N__31821),
            .I(N__31818));
    InMux I__5783 (
            .O(N__31818),
            .I(N__31815));
    LocalMux I__5782 (
            .O(N__31815),
            .I(N__31812));
    Span4Mux_v I__5781 (
            .O(N__31812),
            .I(N__31809));
    Odrv4 I__5780 (
            .O(N__31809),
            .I(\SIG_DDS.n10 ));
    InMux I__5779 (
            .O(N__31806),
            .I(N__31803));
    LocalMux I__5778 (
            .O(N__31803),
            .I(N__31799));
    InMux I__5777 (
            .O(N__31802),
            .I(N__31795));
    Span4Mux_h I__5776 (
            .O(N__31799),
            .I(N__31792));
    InMux I__5775 (
            .O(N__31798),
            .I(N__31789));
    LocalMux I__5774 (
            .O(N__31795),
            .I(buf_dds1_10));
    Odrv4 I__5773 (
            .O(N__31792),
            .I(buf_dds1_10));
    LocalMux I__5772 (
            .O(N__31789),
            .I(buf_dds1_10));
    IoInMux I__5771 (
            .O(N__31782),
            .I(N__31779));
    LocalMux I__5770 (
            .O(N__31779),
            .I(N__31776));
    Span4Mux_s1_v I__5769 (
            .O(N__31776),
            .I(N__31772));
    InMux I__5768 (
            .O(N__31775),
            .I(N__31769));
    Sp12to4 I__5767 (
            .O(N__31772),
            .I(N__31766));
    LocalMux I__5766 (
            .O(N__31769),
            .I(N__31762));
    Span12Mux_h I__5765 (
            .O(N__31766),
            .I(N__31759));
    InMux I__5764 (
            .O(N__31765),
            .I(N__31756));
    Span4Mux_v I__5763 (
            .O(N__31762),
            .I(N__31753));
    Odrv12 I__5762 (
            .O(N__31759),
            .I(SELIRNG0));
    LocalMux I__5761 (
            .O(N__31756),
            .I(SELIRNG0));
    Odrv4 I__5760 (
            .O(N__31753),
            .I(SELIRNG0));
    InMux I__5759 (
            .O(N__31746),
            .I(N__31743));
    LocalMux I__5758 (
            .O(N__31743),
            .I(N__31740));
    Span4Mux_v I__5757 (
            .O(N__31740),
            .I(N__31737));
    Span4Mux_h I__5756 (
            .O(N__31737),
            .I(N__31734));
    Span4Mux_h I__5755 (
            .O(N__31734),
            .I(N__31731));
    Odrv4 I__5754 (
            .O(N__31731),
            .I(buf_data_iac_3));
    InMux I__5753 (
            .O(N__31728),
            .I(N__31725));
    LocalMux I__5752 (
            .O(N__31725),
            .I(n22_adj_1637));
    InMux I__5751 (
            .O(N__31722),
            .I(N__31718));
    InMux I__5750 (
            .O(N__31721),
            .I(N__31715));
    LocalMux I__5749 (
            .O(N__31718),
            .I(N__31712));
    LocalMux I__5748 (
            .O(N__31715),
            .I(N__31706));
    Span4Mux_v I__5747 (
            .O(N__31712),
            .I(N__31706));
    CascadeMux I__5746 (
            .O(N__31711),
            .I(N__31703));
    Span4Mux_h I__5745 (
            .O(N__31706),
            .I(N__31700));
    InMux I__5744 (
            .O(N__31703),
            .I(N__31697));
    Odrv4 I__5743 (
            .O(N__31700),
            .I(cmd_rdadctmp_17_adj_1433));
    LocalMux I__5742 (
            .O(N__31697),
            .I(cmd_rdadctmp_17_adj_1433));
    InMux I__5741 (
            .O(N__31692),
            .I(N__31678));
    InMux I__5740 (
            .O(N__31691),
            .I(N__31678));
    InMux I__5739 (
            .O(N__31690),
            .I(N__31673));
    InMux I__5738 (
            .O(N__31689),
            .I(N__31673));
    InMux I__5737 (
            .O(N__31688),
            .I(N__31661));
    InMux I__5736 (
            .O(N__31687),
            .I(N__31661));
    InMux I__5735 (
            .O(N__31686),
            .I(N__31661));
    InMux I__5734 (
            .O(N__31685),
            .I(N__31648));
    InMux I__5733 (
            .O(N__31684),
            .I(N__31648));
    InMux I__5732 (
            .O(N__31683),
            .I(N__31648));
    LocalMux I__5731 (
            .O(N__31678),
            .I(N__31645));
    LocalMux I__5730 (
            .O(N__31673),
            .I(N__31642));
    InMux I__5729 (
            .O(N__31672),
            .I(N__31637));
    InMux I__5728 (
            .O(N__31671),
            .I(N__31637));
    InMux I__5727 (
            .O(N__31670),
            .I(N__31630));
    InMux I__5726 (
            .O(N__31669),
            .I(N__31630));
    InMux I__5725 (
            .O(N__31668),
            .I(N__31630));
    LocalMux I__5724 (
            .O(N__31661),
            .I(N__31625));
    InMux I__5723 (
            .O(N__31660),
            .I(N__31620));
    InMux I__5722 (
            .O(N__31659),
            .I(N__31620));
    InMux I__5721 (
            .O(N__31658),
            .I(N__31610));
    InMux I__5720 (
            .O(N__31657),
            .I(N__31610));
    InMux I__5719 (
            .O(N__31656),
            .I(N__31610));
    InMux I__5718 (
            .O(N__31655),
            .I(N__31610));
    LocalMux I__5717 (
            .O(N__31648),
            .I(N__31607));
    Span4Mux_v I__5716 (
            .O(N__31645),
            .I(N__31598));
    Span4Mux_h I__5715 (
            .O(N__31642),
            .I(N__31598));
    LocalMux I__5714 (
            .O(N__31637),
            .I(N__31598));
    LocalMux I__5713 (
            .O(N__31630),
            .I(N__31598));
    InMux I__5712 (
            .O(N__31629),
            .I(N__31593));
    InMux I__5711 (
            .O(N__31628),
            .I(N__31593));
    Span4Mux_v I__5710 (
            .O(N__31625),
            .I(N__31587));
    LocalMux I__5709 (
            .O(N__31620),
            .I(N__31587));
    InMux I__5708 (
            .O(N__31619),
            .I(N__31584));
    LocalMux I__5707 (
            .O(N__31610),
            .I(N__31581));
    Span4Mux_v I__5706 (
            .O(N__31607),
            .I(N__31574));
    Span4Mux_h I__5705 (
            .O(N__31598),
            .I(N__31574));
    LocalMux I__5704 (
            .O(N__31593),
            .I(N__31574));
    InMux I__5703 (
            .O(N__31592),
            .I(N__31571));
    Span4Mux_h I__5702 (
            .O(N__31587),
            .I(N__31566));
    LocalMux I__5701 (
            .O(N__31584),
            .I(N__31566));
    Span12Mux_v I__5700 (
            .O(N__31581),
            .I(N__31556));
    Span4Mux_v I__5699 (
            .O(N__31574),
            .I(N__31553));
    LocalMux I__5698 (
            .O(N__31571),
            .I(N__31550));
    Span4Mux_h I__5697 (
            .O(N__31566),
            .I(N__31547));
    InMux I__5696 (
            .O(N__31565),
            .I(N__31542));
    InMux I__5695 (
            .O(N__31564),
            .I(N__31542));
    InMux I__5694 (
            .O(N__31563),
            .I(N__31537));
    InMux I__5693 (
            .O(N__31562),
            .I(N__31537));
    InMux I__5692 (
            .O(N__31561),
            .I(N__31530));
    InMux I__5691 (
            .O(N__31560),
            .I(N__31530));
    InMux I__5690 (
            .O(N__31559),
            .I(N__31530));
    Odrv12 I__5689 (
            .O(N__31556),
            .I(n12653));
    Odrv4 I__5688 (
            .O(N__31553),
            .I(n12653));
    Odrv12 I__5687 (
            .O(N__31550),
            .I(n12653));
    Odrv4 I__5686 (
            .O(N__31547),
            .I(n12653));
    LocalMux I__5685 (
            .O(N__31542),
            .I(n12653));
    LocalMux I__5684 (
            .O(N__31537),
            .I(n12653));
    LocalMux I__5683 (
            .O(N__31530),
            .I(n12653));
    InMux I__5682 (
            .O(N__31515),
            .I(N__31511));
    InMux I__5681 (
            .O(N__31514),
            .I(N__31508));
    LocalMux I__5680 (
            .O(N__31511),
            .I(N__31505));
    LocalMux I__5679 (
            .O(N__31508),
            .I(N__31502));
    Span4Mux_v I__5678 (
            .O(N__31505),
            .I(N__31499));
    Span4Mux_h I__5677 (
            .O(N__31502),
            .I(N__31495));
    Span4Mux_h I__5676 (
            .O(N__31499),
            .I(N__31492));
    InMux I__5675 (
            .O(N__31498),
            .I(N__31489));
    Odrv4 I__5674 (
            .O(N__31495),
            .I(cmd_rdadctmp_19_adj_1431));
    Odrv4 I__5673 (
            .O(N__31492),
            .I(cmd_rdadctmp_19_adj_1431));
    LocalMux I__5672 (
            .O(N__31489),
            .I(cmd_rdadctmp_19_adj_1431));
    InMux I__5671 (
            .O(N__31482),
            .I(N__31478));
    InMux I__5670 (
            .O(N__31481),
            .I(N__31475));
    LocalMux I__5669 (
            .O(N__31478),
            .I(secclk_cnt_21));
    LocalMux I__5668 (
            .O(N__31475),
            .I(secclk_cnt_21));
    InMux I__5667 (
            .O(N__31470),
            .I(N__31466));
    InMux I__5666 (
            .O(N__31469),
            .I(N__31463));
    LocalMux I__5665 (
            .O(N__31466),
            .I(secclk_cnt_19));
    LocalMux I__5664 (
            .O(N__31463),
            .I(secclk_cnt_19));
    CascadeMux I__5663 (
            .O(N__31458),
            .I(N__31454));
    InMux I__5662 (
            .O(N__31457),
            .I(N__31451));
    InMux I__5661 (
            .O(N__31454),
            .I(N__31448));
    LocalMux I__5660 (
            .O(N__31451),
            .I(secclk_cnt_12));
    LocalMux I__5659 (
            .O(N__31448),
            .I(secclk_cnt_12));
    InMux I__5658 (
            .O(N__31443),
            .I(N__31439));
    InMux I__5657 (
            .O(N__31442),
            .I(N__31436));
    LocalMux I__5656 (
            .O(N__31439),
            .I(secclk_cnt_22));
    LocalMux I__5655 (
            .O(N__31436),
            .I(secclk_cnt_22));
    InMux I__5654 (
            .O(N__31431),
            .I(N__31428));
    LocalMux I__5653 (
            .O(N__31428),
            .I(N__31425));
    Odrv4 I__5652 (
            .O(N__31425),
            .I(n14_adj_1599));
    InMux I__5651 (
            .O(N__31422),
            .I(N__31419));
    LocalMux I__5650 (
            .O(N__31419),
            .I(N__31415));
    InMux I__5649 (
            .O(N__31418),
            .I(N__31412));
    Sp12to4 I__5648 (
            .O(N__31415),
            .I(N__31407));
    LocalMux I__5647 (
            .O(N__31412),
            .I(N__31407));
    Odrv12 I__5646 (
            .O(N__31407),
            .I(\comm_spi.n14610 ));
    InMux I__5645 (
            .O(N__31404),
            .I(N__31400));
    CascadeMux I__5644 (
            .O(N__31403),
            .I(N__31397));
    LocalMux I__5643 (
            .O(N__31400),
            .I(N__31394));
    InMux I__5642 (
            .O(N__31397),
            .I(N__31391));
    Odrv12 I__5641 (
            .O(N__31394),
            .I(buf_readRTD_14));
    LocalMux I__5640 (
            .O(N__31391),
            .I(buf_readRTD_14));
    InMux I__5639 (
            .O(N__31386),
            .I(N__31382));
    CascadeMux I__5638 (
            .O(N__31385),
            .I(N__31379));
    LocalMux I__5637 (
            .O(N__31382),
            .I(N__31375));
    InMux I__5636 (
            .O(N__31379),
            .I(N__31372));
    InMux I__5635 (
            .O(N__31378),
            .I(N__31368));
    Span4Mux_h I__5634 (
            .O(N__31375),
            .I(N__31365));
    LocalMux I__5633 (
            .O(N__31372),
            .I(N__31362));
    InMux I__5632 (
            .O(N__31371),
            .I(N__31359));
    LocalMux I__5631 (
            .O(N__31368),
            .I(N__31356));
    Span4Mux_v I__5630 (
            .O(N__31365),
            .I(N__31353));
    Span4Mux_v I__5629 (
            .O(N__31362),
            .I(N__31349));
    LocalMux I__5628 (
            .O(N__31359),
            .I(N__31346));
    Span12Mux_s11_h I__5627 (
            .O(N__31356),
            .I(N__31343));
    Span4Mux_v I__5626 (
            .O(N__31353),
            .I(N__31340));
    InMux I__5625 (
            .O(N__31352),
            .I(N__31337));
    Span4Mux_h I__5624 (
            .O(N__31349),
            .I(N__31332));
    Span4Mux_h I__5623 (
            .O(N__31346),
            .I(N__31332));
    Odrv12 I__5622 (
            .O(N__31343),
            .I(buf_cfgRTD_6));
    Odrv4 I__5621 (
            .O(N__31340),
            .I(buf_cfgRTD_6));
    LocalMux I__5620 (
            .O(N__31337),
            .I(buf_cfgRTD_6));
    Odrv4 I__5619 (
            .O(N__31332),
            .I(buf_cfgRTD_6));
    InMux I__5618 (
            .O(N__31323),
            .I(N__31320));
    LocalMux I__5617 (
            .O(N__31320),
            .I(N__31316));
    CascadeMux I__5616 (
            .O(N__31319),
            .I(N__31313));
    Span4Mux_h I__5615 (
            .O(N__31316),
            .I(N__31310));
    InMux I__5614 (
            .O(N__31313),
            .I(N__31307));
    Odrv4 I__5613 (
            .O(N__31310),
            .I(buf_readRTD_15));
    LocalMux I__5612 (
            .O(N__31307),
            .I(buf_readRTD_15));
    CascadeMux I__5611 (
            .O(N__31302),
            .I(N__31297));
    InMux I__5610 (
            .O(N__31301),
            .I(N__31294));
    CascadeMux I__5609 (
            .O(N__31300),
            .I(N__31291));
    InMux I__5608 (
            .O(N__31297),
            .I(N__31288));
    LocalMux I__5607 (
            .O(N__31294),
            .I(N__31284));
    InMux I__5606 (
            .O(N__31291),
            .I(N__31281));
    LocalMux I__5605 (
            .O(N__31288),
            .I(N__31277));
    InMux I__5604 (
            .O(N__31287),
            .I(N__31274));
    Sp12to4 I__5603 (
            .O(N__31284),
            .I(N__31269));
    LocalMux I__5602 (
            .O(N__31281),
            .I(N__31269));
    CascadeMux I__5601 (
            .O(N__31280),
            .I(N__31266));
    Span4Mux_v I__5600 (
            .O(N__31277),
            .I(N__31263));
    LocalMux I__5599 (
            .O(N__31274),
            .I(N__31260));
    Span12Mux_v I__5598 (
            .O(N__31269),
            .I(N__31257));
    InMux I__5597 (
            .O(N__31266),
            .I(N__31254));
    Span4Mux_h I__5596 (
            .O(N__31263),
            .I(N__31249));
    Span4Mux_h I__5595 (
            .O(N__31260),
            .I(N__31249));
    Odrv12 I__5594 (
            .O(N__31257),
            .I(buf_cfgRTD_7));
    LocalMux I__5593 (
            .O(N__31254),
            .I(buf_cfgRTD_7));
    Odrv4 I__5592 (
            .O(N__31249),
            .I(buf_cfgRTD_7));
    CascadeMux I__5591 (
            .O(N__31242),
            .I(N__31239));
    InMux I__5590 (
            .O(N__31239),
            .I(N__31236));
    LocalMux I__5589 (
            .O(N__31236),
            .I(N__31233));
    Span4Mux_h I__5588 (
            .O(N__31233),
            .I(N__31230));
    Odrv4 I__5587 (
            .O(N__31230),
            .I(n20_adj_1528));
    InMux I__5586 (
            .O(N__31227),
            .I(N__31223));
    InMux I__5585 (
            .O(N__31226),
            .I(N__31220));
    LocalMux I__5584 (
            .O(N__31223),
            .I(secclk_cnt_16));
    LocalMux I__5583 (
            .O(N__31220),
            .I(secclk_cnt_16));
    InMux I__5582 (
            .O(N__31215),
            .I(N__31211));
    InMux I__5581 (
            .O(N__31214),
            .I(N__31208));
    LocalMux I__5580 (
            .O(N__31211),
            .I(secclk_cnt_2));
    LocalMux I__5579 (
            .O(N__31208),
            .I(secclk_cnt_2));
    CascadeMux I__5578 (
            .O(N__31203),
            .I(N__31200));
    InMux I__5577 (
            .O(N__31200),
            .I(N__31196));
    InMux I__5576 (
            .O(N__31199),
            .I(N__31193));
    LocalMux I__5575 (
            .O(N__31196),
            .I(secclk_cnt_7));
    LocalMux I__5574 (
            .O(N__31193),
            .I(secclk_cnt_7));
    InMux I__5573 (
            .O(N__31188),
            .I(N__31184));
    InMux I__5572 (
            .O(N__31187),
            .I(N__31181));
    LocalMux I__5571 (
            .O(N__31184),
            .I(secclk_cnt_13));
    LocalMux I__5570 (
            .O(N__31181),
            .I(secclk_cnt_13));
    InMux I__5569 (
            .O(N__31176),
            .I(N__31173));
    LocalMux I__5568 (
            .O(N__31173),
            .I(n27_adj_1597));
    CascadeMux I__5567 (
            .O(N__31170),
            .I(n26_adj_1575_cascade_));
    InMux I__5566 (
            .O(N__31167),
            .I(N__31164));
    LocalMux I__5565 (
            .O(N__31164),
            .I(n25_adj_1574));
    CascadeMux I__5564 (
            .O(N__31161),
            .I(n19856_cascade_));
    InMux I__5563 (
            .O(N__31158),
            .I(N__31154));
    InMux I__5562 (
            .O(N__31157),
            .I(N__31151));
    LocalMux I__5561 (
            .O(N__31154),
            .I(secclk_cnt_20));
    LocalMux I__5560 (
            .O(N__31151),
            .I(secclk_cnt_20));
    SRMux I__5559 (
            .O(N__31146),
            .I(N__31142));
    SRMux I__5558 (
            .O(N__31145),
            .I(N__31139));
    LocalMux I__5557 (
            .O(N__31142),
            .I(N__31134));
    LocalMux I__5556 (
            .O(N__31139),
            .I(N__31131));
    SRMux I__5555 (
            .O(N__31138),
            .I(N__31128));
    InMux I__5554 (
            .O(N__31137),
            .I(N__31125));
    Span4Mux_v I__5553 (
            .O(N__31134),
            .I(N__31122));
    Span4Mux_h I__5552 (
            .O(N__31131),
            .I(N__31117));
    LocalMux I__5551 (
            .O(N__31128),
            .I(N__31117));
    LocalMux I__5550 (
            .O(N__31125),
            .I(N__31114));
    Odrv4 I__5549 (
            .O(N__31122),
            .I(n14715));
    Odrv4 I__5548 (
            .O(N__31117),
            .I(n14715));
    Odrv12 I__5547 (
            .O(N__31114),
            .I(n14715));
    InMux I__5546 (
            .O(N__31107),
            .I(N__31103));
    InMux I__5545 (
            .O(N__31106),
            .I(N__31100));
    LocalMux I__5544 (
            .O(N__31103),
            .I(secclk_cnt_0));
    LocalMux I__5543 (
            .O(N__31100),
            .I(secclk_cnt_0));
    InMux I__5542 (
            .O(N__31095),
            .I(N__31091));
    InMux I__5541 (
            .O(N__31094),
            .I(N__31088));
    LocalMux I__5540 (
            .O(N__31091),
            .I(secclk_cnt_18));
    LocalMux I__5539 (
            .O(N__31088),
            .I(secclk_cnt_18));
    CascadeMux I__5538 (
            .O(N__31083),
            .I(N__31079));
    InMux I__5537 (
            .O(N__31082),
            .I(N__31076));
    InMux I__5536 (
            .O(N__31079),
            .I(N__31073));
    LocalMux I__5535 (
            .O(N__31076),
            .I(secclk_cnt_11));
    LocalMux I__5534 (
            .O(N__31073),
            .I(secclk_cnt_11));
    InMux I__5533 (
            .O(N__31068),
            .I(N__31064));
    InMux I__5532 (
            .O(N__31067),
            .I(N__31061));
    LocalMux I__5531 (
            .O(N__31064),
            .I(secclk_cnt_4));
    LocalMux I__5530 (
            .O(N__31061),
            .I(secclk_cnt_4));
    InMux I__5529 (
            .O(N__31056),
            .I(N__31053));
    LocalMux I__5528 (
            .O(N__31053),
            .I(n28_adj_1505));
    InMux I__5527 (
            .O(N__31050),
            .I(N__31047));
    LocalMux I__5526 (
            .O(N__31047),
            .I(N__31044));
    Span4Mux_h I__5525 (
            .O(N__31044),
            .I(N__31041));
    Span4Mux_h I__5524 (
            .O(N__31041),
            .I(N__31036));
    InMux I__5523 (
            .O(N__31040),
            .I(N__31033));
    InMux I__5522 (
            .O(N__31039),
            .I(N__31030));
    Span4Mux_h I__5521 (
            .O(N__31036),
            .I(N__31027));
    LocalMux I__5520 (
            .O(N__31033),
            .I(N__31024));
    LocalMux I__5519 (
            .O(N__31030),
            .I(buf_adcdata_iac_3));
    Odrv4 I__5518 (
            .O(N__31027),
            .I(buf_adcdata_iac_3));
    Odrv4 I__5517 (
            .O(N__31024),
            .I(buf_adcdata_iac_3));
    InMux I__5516 (
            .O(N__31017),
            .I(N__31014));
    LocalMux I__5515 (
            .O(N__31014),
            .I(N__31011));
    Odrv4 I__5514 (
            .O(N__31011),
            .I(n19_adj_1636));
    InMux I__5513 (
            .O(N__31008),
            .I(N__31004));
    InMux I__5512 (
            .O(N__31007),
            .I(N__31001));
    LocalMux I__5511 (
            .O(N__31004),
            .I(secclk_cnt_17));
    LocalMux I__5510 (
            .O(N__31001),
            .I(secclk_cnt_17));
    InMux I__5509 (
            .O(N__30996),
            .I(N__30992));
    InMux I__5508 (
            .O(N__30995),
            .I(N__30989));
    LocalMux I__5507 (
            .O(N__30992),
            .I(secclk_cnt_9));
    LocalMux I__5506 (
            .O(N__30989),
            .I(secclk_cnt_9));
    InMux I__5505 (
            .O(N__30984),
            .I(N__30981));
    LocalMux I__5504 (
            .O(N__30981),
            .I(n10_adj_1601));
    InMux I__5503 (
            .O(N__30978),
            .I(N__30975));
    LocalMux I__5502 (
            .O(N__30975),
            .I(N__30971));
    InMux I__5501 (
            .O(N__30974),
            .I(N__30968));
    Odrv12 I__5500 (
            .O(N__30971),
            .I(dds0_mclkcnt_6));
    LocalMux I__5499 (
            .O(N__30968),
            .I(dds0_mclkcnt_6));
    InMux I__5498 (
            .O(N__30963),
            .I(N__30960));
    LocalMux I__5497 (
            .O(N__30960),
            .I(N__30957));
    Odrv12 I__5496 (
            .O(N__30957),
            .I(n20799));
    InMux I__5495 (
            .O(N__30954),
            .I(N__30950));
    InMux I__5494 (
            .O(N__30953),
            .I(N__30947));
    LocalMux I__5493 (
            .O(N__30950),
            .I(secclk_cnt_6));
    LocalMux I__5492 (
            .O(N__30947),
            .I(secclk_cnt_6));
    InMux I__5491 (
            .O(N__30942),
            .I(N__30938));
    InMux I__5490 (
            .O(N__30941),
            .I(N__30935));
    LocalMux I__5489 (
            .O(N__30938),
            .I(secclk_cnt_14));
    LocalMux I__5488 (
            .O(N__30935),
            .I(secclk_cnt_14));
    CascadeMux I__5487 (
            .O(N__30930),
            .I(N__30926));
    InMux I__5486 (
            .O(N__30929),
            .I(N__30923));
    InMux I__5485 (
            .O(N__30926),
            .I(N__30920));
    LocalMux I__5484 (
            .O(N__30923),
            .I(secclk_cnt_10));
    LocalMux I__5483 (
            .O(N__30920),
            .I(secclk_cnt_10));
    InMux I__5482 (
            .O(N__30915),
            .I(N__30911));
    InMux I__5481 (
            .O(N__30914),
            .I(N__30908));
    LocalMux I__5480 (
            .O(N__30911),
            .I(secclk_cnt_3));
    LocalMux I__5479 (
            .O(N__30908),
            .I(secclk_cnt_3));
    InMux I__5478 (
            .O(N__30903),
            .I(N__30899));
    InMux I__5477 (
            .O(N__30902),
            .I(N__30896));
    LocalMux I__5476 (
            .O(N__30899),
            .I(secclk_cnt_15));
    LocalMux I__5475 (
            .O(N__30896),
            .I(secclk_cnt_15));
    InMux I__5474 (
            .O(N__30891),
            .I(N__30887));
    InMux I__5473 (
            .O(N__30890),
            .I(N__30884));
    LocalMux I__5472 (
            .O(N__30887),
            .I(secclk_cnt_8));
    LocalMux I__5471 (
            .O(N__30884),
            .I(secclk_cnt_8));
    CascadeMux I__5470 (
            .O(N__30879),
            .I(N__30875));
    InMux I__5469 (
            .O(N__30878),
            .I(N__30872));
    InMux I__5468 (
            .O(N__30875),
            .I(N__30869));
    LocalMux I__5467 (
            .O(N__30872),
            .I(secclk_cnt_1));
    LocalMux I__5466 (
            .O(N__30869),
            .I(secclk_cnt_1));
    InMux I__5465 (
            .O(N__30864),
            .I(N__30860));
    InMux I__5464 (
            .O(N__30863),
            .I(N__30857));
    LocalMux I__5463 (
            .O(N__30860),
            .I(secclk_cnt_5));
    LocalMux I__5462 (
            .O(N__30857),
            .I(secclk_cnt_5));
    InMux I__5461 (
            .O(N__30852),
            .I(N__30848));
    InMux I__5460 (
            .O(N__30851),
            .I(N__30845));
    LocalMux I__5459 (
            .O(N__30848),
            .I(dds0_mclkcnt_5));
    LocalMux I__5458 (
            .O(N__30845),
            .I(dds0_mclkcnt_5));
    CascadeMux I__5457 (
            .O(N__30840),
            .I(N__30836));
    InMux I__5456 (
            .O(N__30839),
            .I(N__30833));
    InMux I__5455 (
            .O(N__30836),
            .I(N__30830));
    LocalMux I__5454 (
            .O(N__30833),
            .I(dds0_mclkcnt_1));
    LocalMux I__5453 (
            .O(N__30830),
            .I(dds0_mclkcnt_1));
    InMux I__5452 (
            .O(N__30825),
            .I(N__30821));
    InMux I__5451 (
            .O(N__30824),
            .I(N__30818));
    LocalMux I__5450 (
            .O(N__30821),
            .I(dds0_mclkcnt_4));
    LocalMux I__5449 (
            .O(N__30818),
            .I(dds0_mclkcnt_4));
    InMux I__5448 (
            .O(N__30813),
            .I(N__30809));
    InMux I__5447 (
            .O(N__30812),
            .I(N__30806));
    LocalMux I__5446 (
            .O(N__30809),
            .I(dds0_mclkcnt_2));
    LocalMux I__5445 (
            .O(N__30806),
            .I(dds0_mclkcnt_2));
    InMux I__5444 (
            .O(N__30801),
            .I(N__30797));
    InMux I__5443 (
            .O(N__30800),
            .I(N__30794));
    LocalMux I__5442 (
            .O(N__30797),
            .I(dds0_mclkcnt_0));
    LocalMux I__5441 (
            .O(N__30794),
            .I(dds0_mclkcnt_0));
    CascadeMux I__5440 (
            .O(N__30789),
            .I(n12_adj_1480_cascade_));
    InMux I__5439 (
            .O(N__30786),
            .I(N__30782));
    InMux I__5438 (
            .O(N__30785),
            .I(N__30779));
    LocalMux I__5437 (
            .O(N__30782),
            .I(dds0_mclkcnt_7));
    LocalMux I__5436 (
            .O(N__30779),
            .I(dds0_mclkcnt_7));
    CascadeMux I__5435 (
            .O(N__30774),
            .I(n20799_cascade_));
    InMux I__5434 (
            .O(N__30771),
            .I(N__30768));
    LocalMux I__5433 (
            .O(N__30768),
            .I(n10));
    InMux I__5432 (
            .O(N__30765),
            .I(N__30762));
    LocalMux I__5431 (
            .O(N__30762),
            .I(N__30758));
    InMux I__5430 (
            .O(N__30761),
            .I(N__30755));
    Odrv4 I__5429 (
            .O(N__30758),
            .I(\comm_spi.n14611 ));
    LocalMux I__5428 (
            .O(N__30755),
            .I(\comm_spi.n14611 ));
    InMux I__5427 (
            .O(N__30750),
            .I(N__30746));
    CEMux I__5426 (
            .O(N__30749),
            .I(N__30743));
    LocalMux I__5425 (
            .O(N__30746),
            .I(N__30740));
    LocalMux I__5424 (
            .O(N__30743),
            .I(N__30737));
    Span12Mux_h I__5423 (
            .O(N__30740),
            .I(N__30734));
    Odrv4 I__5422 (
            .O(N__30737),
            .I(\ADC_VAC.n12594 ));
    Odrv12 I__5421 (
            .O(N__30734),
            .I(\ADC_VAC.n12594 ));
    InMux I__5420 (
            .O(N__30729),
            .I(N__30725));
    InMux I__5419 (
            .O(N__30728),
            .I(N__30722));
    LocalMux I__5418 (
            .O(N__30725),
            .I(N__30717));
    LocalMux I__5417 (
            .O(N__30722),
            .I(N__30714));
    InMux I__5416 (
            .O(N__30721),
            .I(N__30710));
    CascadeMux I__5415 (
            .O(N__30720),
            .I(N__30703));
    Span4Mux_v I__5414 (
            .O(N__30717),
            .I(N__30697));
    Sp12to4 I__5413 (
            .O(N__30714),
            .I(N__30694));
    InMux I__5412 (
            .O(N__30713),
            .I(N__30691));
    LocalMux I__5411 (
            .O(N__30710),
            .I(N__30688));
    InMux I__5410 (
            .O(N__30709),
            .I(N__30685));
    InMux I__5409 (
            .O(N__30708),
            .I(N__30682));
    InMux I__5408 (
            .O(N__30707),
            .I(N__30679));
    InMux I__5407 (
            .O(N__30706),
            .I(N__30676));
    InMux I__5406 (
            .O(N__30703),
            .I(N__30673));
    InMux I__5405 (
            .O(N__30702),
            .I(N__30666));
    InMux I__5404 (
            .O(N__30701),
            .I(N__30666));
    InMux I__5403 (
            .O(N__30700),
            .I(N__30666));
    Sp12to4 I__5402 (
            .O(N__30697),
            .I(N__30661));
    Span12Mux_v I__5401 (
            .O(N__30694),
            .I(N__30661));
    LocalMux I__5400 (
            .O(N__30691),
            .I(N__30654));
    Span4Mux_v I__5399 (
            .O(N__30688),
            .I(N__30654));
    LocalMux I__5398 (
            .O(N__30685),
            .I(N__30654));
    LocalMux I__5397 (
            .O(N__30682),
            .I(DTRIG_N_918_adj_1451));
    LocalMux I__5396 (
            .O(N__30679),
            .I(DTRIG_N_918_adj_1451));
    LocalMux I__5395 (
            .O(N__30676),
            .I(DTRIG_N_918_adj_1451));
    LocalMux I__5394 (
            .O(N__30673),
            .I(DTRIG_N_918_adj_1451));
    LocalMux I__5393 (
            .O(N__30666),
            .I(DTRIG_N_918_adj_1451));
    Odrv12 I__5392 (
            .O(N__30661),
            .I(DTRIG_N_918_adj_1451));
    Odrv4 I__5391 (
            .O(N__30654),
            .I(DTRIG_N_918_adj_1451));
    SRMux I__5390 (
            .O(N__30639),
            .I(N__30636));
    LocalMux I__5389 (
            .O(N__30636),
            .I(N__30633));
    Span4Mux_v I__5388 (
            .O(N__30633),
            .I(N__30630));
    Span4Mux_h I__5387 (
            .O(N__30630),
            .I(N__30627));
    Span4Mux_v I__5386 (
            .O(N__30627),
            .I(N__30624));
    Odrv4 I__5385 (
            .O(N__30624),
            .I(\ADC_VAC.n14844 ));
    InMux I__5384 (
            .O(N__30621),
            .I(n19741));
    InMux I__5383 (
            .O(N__30618),
            .I(n19742));
    InMux I__5382 (
            .O(N__30615),
            .I(n19743));
    InMux I__5381 (
            .O(N__30612),
            .I(n19744));
    InMux I__5380 (
            .O(N__30609),
            .I(n19745));
    InMux I__5379 (
            .O(N__30606),
            .I(N__30602));
    InMux I__5378 (
            .O(N__30605),
            .I(N__30599));
    LocalMux I__5377 (
            .O(N__30602),
            .I(clk_cnt_0));
    LocalMux I__5376 (
            .O(N__30599),
            .I(clk_cnt_0));
    InMux I__5375 (
            .O(N__30594),
            .I(N__30590));
    InMux I__5374 (
            .O(N__30593),
            .I(N__30587));
    LocalMux I__5373 (
            .O(N__30590),
            .I(clk_cnt_4));
    LocalMux I__5372 (
            .O(N__30587),
            .I(clk_cnt_4));
    InMux I__5371 (
            .O(N__30582),
            .I(N__30578));
    InMux I__5370 (
            .O(N__30581),
            .I(N__30575));
    LocalMux I__5369 (
            .O(N__30578),
            .I(clk_cnt_2));
    LocalMux I__5368 (
            .O(N__30575),
            .I(clk_cnt_2));
    InMux I__5367 (
            .O(N__30570),
            .I(N__30566));
    InMux I__5366 (
            .O(N__30569),
            .I(N__30563));
    LocalMux I__5365 (
            .O(N__30566),
            .I(clk_cnt_1));
    LocalMux I__5364 (
            .O(N__30563),
            .I(clk_cnt_1));
    CascadeMux I__5363 (
            .O(N__30558),
            .I(n6_cascade_));
    InMux I__5362 (
            .O(N__30555),
            .I(N__30551));
    InMux I__5361 (
            .O(N__30554),
            .I(N__30548));
    LocalMux I__5360 (
            .O(N__30551),
            .I(clk_cnt_3));
    LocalMux I__5359 (
            .O(N__30548),
            .I(clk_cnt_3));
    SRMux I__5358 (
            .O(N__30543),
            .I(N__30540));
    LocalMux I__5357 (
            .O(N__30540),
            .I(N__30537));
    Sp12to4 I__5356 (
            .O(N__30537),
            .I(N__30534));
    Odrv12 I__5355 (
            .O(N__30534),
            .I(n14714));
    CascadeMux I__5354 (
            .O(N__30531),
            .I(n14714_cascade_));
    ClkMux I__5353 (
            .O(N__30528),
            .I(N__30522));
    ClkMux I__5352 (
            .O(N__30527),
            .I(N__30519));
    ClkMux I__5351 (
            .O(N__30526),
            .I(N__30514));
    ClkMux I__5350 (
            .O(N__30525),
            .I(N__30510));
    LocalMux I__5349 (
            .O(N__30522),
            .I(N__30501));
    LocalMux I__5348 (
            .O(N__30519),
            .I(N__30501));
    ClkMux I__5347 (
            .O(N__30518),
            .I(N__30498));
    ClkMux I__5346 (
            .O(N__30517),
            .I(N__30495));
    LocalMux I__5345 (
            .O(N__30514),
            .I(N__30489));
    ClkMux I__5344 (
            .O(N__30513),
            .I(N__30486));
    LocalMux I__5343 (
            .O(N__30510),
            .I(N__30483));
    ClkMux I__5342 (
            .O(N__30509),
            .I(N__30480));
    ClkMux I__5341 (
            .O(N__30508),
            .I(N__30477));
    ClkMux I__5340 (
            .O(N__30507),
            .I(N__30473));
    ClkMux I__5339 (
            .O(N__30506),
            .I(N__30469));
    Span4Mux_v I__5338 (
            .O(N__30501),
            .I(N__30460));
    LocalMux I__5337 (
            .O(N__30498),
            .I(N__30460));
    LocalMux I__5336 (
            .O(N__30495),
            .I(N__30460));
    ClkMux I__5335 (
            .O(N__30494),
            .I(N__30456));
    ClkMux I__5334 (
            .O(N__30493),
            .I(N__30453));
    ClkMux I__5333 (
            .O(N__30492),
            .I(N__30450));
    Span4Mux_v I__5332 (
            .O(N__30489),
            .I(N__30446));
    LocalMux I__5331 (
            .O(N__30486),
            .I(N__30443));
    Span4Mux_h I__5330 (
            .O(N__30483),
            .I(N__30438));
    LocalMux I__5329 (
            .O(N__30480),
            .I(N__30438));
    LocalMux I__5328 (
            .O(N__30477),
            .I(N__30435));
    ClkMux I__5327 (
            .O(N__30476),
            .I(N__30432));
    LocalMux I__5326 (
            .O(N__30473),
            .I(N__30429));
    ClkMux I__5325 (
            .O(N__30472),
            .I(N__30426));
    LocalMux I__5324 (
            .O(N__30469),
            .I(N__30423));
    ClkMux I__5323 (
            .O(N__30468),
            .I(N__30420));
    ClkMux I__5322 (
            .O(N__30467),
            .I(N__30417));
    Span4Mux_v I__5321 (
            .O(N__30460),
            .I(N__30413));
    ClkMux I__5320 (
            .O(N__30459),
            .I(N__30410));
    LocalMux I__5319 (
            .O(N__30456),
            .I(N__30403));
    LocalMux I__5318 (
            .O(N__30453),
            .I(N__30403));
    LocalMux I__5317 (
            .O(N__30450),
            .I(N__30403));
    ClkMux I__5316 (
            .O(N__30449),
            .I(N__30400));
    Span4Mux_h I__5315 (
            .O(N__30446),
            .I(N__30395));
    Span4Mux_v I__5314 (
            .O(N__30443),
            .I(N__30395));
    Span4Mux_v I__5313 (
            .O(N__30438),
            .I(N__30392));
    Span4Mux_h I__5312 (
            .O(N__30435),
            .I(N__30387));
    LocalMux I__5311 (
            .O(N__30432),
            .I(N__30387));
    Span4Mux_v I__5310 (
            .O(N__30429),
            .I(N__30382));
    LocalMux I__5309 (
            .O(N__30426),
            .I(N__30382));
    Span4Mux_v I__5308 (
            .O(N__30423),
            .I(N__30375));
    LocalMux I__5307 (
            .O(N__30420),
            .I(N__30375));
    LocalMux I__5306 (
            .O(N__30417),
            .I(N__30375));
    ClkMux I__5305 (
            .O(N__30416),
            .I(N__30372));
    Span4Mux_h I__5304 (
            .O(N__30413),
            .I(N__30369));
    LocalMux I__5303 (
            .O(N__30410),
            .I(N__30362));
    Sp12to4 I__5302 (
            .O(N__30403),
            .I(N__30362));
    LocalMux I__5301 (
            .O(N__30400),
            .I(N__30362));
    Span4Mux_h I__5300 (
            .O(N__30395),
            .I(N__30359));
    Span4Mux_h I__5299 (
            .O(N__30392),
            .I(N__30354));
    Span4Mux_h I__5298 (
            .O(N__30387),
            .I(N__30354));
    Span4Mux_h I__5297 (
            .O(N__30382),
            .I(N__30347));
    Span4Mux_v I__5296 (
            .O(N__30375),
            .I(N__30347));
    LocalMux I__5295 (
            .O(N__30372),
            .I(N__30347));
    Sp12to4 I__5294 (
            .O(N__30369),
            .I(N__30341));
    Span12Mux_v I__5293 (
            .O(N__30362),
            .I(N__30341));
    Span4Mux_v I__5292 (
            .O(N__30359),
            .I(N__30336));
    Span4Mux_h I__5291 (
            .O(N__30354),
            .I(N__30336));
    Span4Mux_h I__5290 (
            .O(N__30347),
            .I(N__30333));
    InMux I__5289 (
            .O(N__30346),
            .I(N__30330));
    Odrv12 I__5288 (
            .O(N__30341),
            .I(clk_RTD));
    Odrv4 I__5287 (
            .O(N__30336),
            .I(clk_RTD));
    Odrv4 I__5286 (
            .O(N__30333),
            .I(clk_RTD));
    LocalMux I__5285 (
            .O(N__30330),
            .I(clk_RTD));
    InMux I__5284 (
            .O(N__30321),
            .I(N__30317));
    InMux I__5283 (
            .O(N__30320),
            .I(N__30314));
    LocalMux I__5282 (
            .O(N__30317),
            .I(dds0_mclkcnt_3));
    LocalMux I__5281 (
            .O(N__30314),
            .I(dds0_mclkcnt_3));
    InMux I__5280 (
            .O(N__30309),
            .I(N__30303));
    InMux I__5279 (
            .O(N__30308),
            .I(N__30299));
    InMux I__5278 (
            .O(N__30307),
            .I(N__30290));
    InMux I__5277 (
            .O(N__30306),
            .I(N__30290));
    LocalMux I__5276 (
            .O(N__30303),
            .I(N__30287));
    CascadeMux I__5275 (
            .O(N__30302),
            .I(N__30282));
    LocalMux I__5274 (
            .O(N__30299),
            .I(N__30278));
    CascadeMux I__5273 (
            .O(N__30298),
            .I(N__30275));
    InMux I__5272 (
            .O(N__30297),
            .I(N__30267));
    InMux I__5271 (
            .O(N__30296),
            .I(N__30267));
    InMux I__5270 (
            .O(N__30295),
            .I(N__30264));
    LocalMux I__5269 (
            .O(N__30290),
            .I(N__30259));
    Span4Mux_v I__5268 (
            .O(N__30287),
            .I(N__30259));
    InMux I__5267 (
            .O(N__30286),
            .I(N__30250));
    InMux I__5266 (
            .O(N__30285),
            .I(N__30250));
    InMux I__5265 (
            .O(N__30282),
            .I(N__30250));
    InMux I__5264 (
            .O(N__30281),
            .I(N__30250));
    Span4Mux_h I__5263 (
            .O(N__30278),
            .I(N__30247));
    InMux I__5262 (
            .O(N__30275),
            .I(N__30244));
    InMux I__5261 (
            .O(N__30274),
            .I(N__30239));
    InMux I__5260 (
            .O(N__30273),
            .I(N__30239));
    InMux I__5259 (
            .O(N__30272),
            .I(N__30236));
    LocalMux I__5258 (
            .O(N__30267),
            .I(N__30233));
    LocalMux I__5257 (
            .O(N__30264),
            .I(N__30226));
    Span4Mux_v I__5256 (
            .O(N__30259),
            .I(N__30226));
    LocalMux I__5255 (
            .O(N__30250),
            .I(N__30226));
    Odrv4 I__5254 (
            .O(N__30247),
            .I(eis_end_N_724));
    LocalMux I__5253 (
            .O(N__30244),
            .I(eis_end_N_724));
    LocalMux I__5252 (
            .O(N__30239),
            .I(eis_end_N_724));
    LocalMux I__5251 (
            .O(N__30236),
            .I(eis_end_N_724));
    Odrv12 I__5250 (
            .O(N__30233),
            .I(eis_end_N_724));
    Odrv4 I__5249 (
            .O(N__30226),
            .I(eis_end_N_724));
    CascadeMux I__5248 (
            .O(N__30213),
            .I(\ADC_VDC.n10119_cascade_ ));
    CEMux I__5247 (
            .O(N__30210),
            .I(N__30207));
    LocalMux I__5246 (
            .O(N__30207),
            .I(\ADC_VDC.n12807 ));
    InMux I__5245 (
            .O(N__30204),
            .I(bfn_12_4_0_));
    InMux I__5244 (
            .O(N__30201),
            .I(n19739));
    InMux I__5243 (
            .O(N__30198),
            .I(n19740));
    InMux I__5242 (
            .O(N__30195),
            .I(N__30192));
    LocalMux I__5241 (
            .O(N__30192),
            .I(N__30188));
    InMux I__5240 (
            .O(N__30191),
            .I(N__30185));
    Odrv4 I__5239 (
            .O(N__30188),
            .I(n20915));
    LocalMux I__5238 (
            .O(N__30185),
            .I(n20915));
    InMux I__5237 (
            .O(N__30180),
            .I(N__30177));
    LocalMux I__5236 (
            .O(N__30177),
            .I(N__30174));
    Odrv4 I__5235 (
            .O(N__30174),
            .I(n20985));
    InMux I__5234 (
            .O(N__30171),
            .I(N__30167));
    InMux I__5233 (
            .O(N__30170),
            .I(N__30164));
    LocalMux I__5232 (
            .O(N__30167),
            .I(n16571));
    LocalMux I__5231 (
            .O(N__30164),
            .I(n16571));
    CascadeMux I__5230 (
            .O(N__30159),
            .I(n13_cascade_));
    InMux I__5229 (
            .O(N__30156),
            .I(N__30153));
    LocalMux I__5228 (
            .O(N__30153),
            .I(n21337));
    InMux I__5227 (
            .O(N__30150),
            .I(N__30147));
    LocalMux I__5226 (
            .O(N__30147),
            .I(N__30144));
    Odrv4 I__5225 (
            .O(N__30144),
            .I(n17507));
    CascadeMux I__5224 (
            .O(N__30141),
            .I(N__30136));
    InMux I__5223 (
            .O(N__30140),
            .I(N__30128));
    InMux I__5222 (
            .O(N__30139),
            .I(N__30128));
    InMux I__5221 (
            .O(N__30136),
            .I(N__30128));
    CascadeMux I__5220 (
            .O(N__30135),
            .I(N__30123));
    LocalMux I__5219 (
            .O(N__30128),
            .I(N__30119));
    InMux I__5218 (
            .O(N__30127),
            .I(N__30111));
    InMux I__5217 (
            .O(N__30126),
            .I(N__30108));
    InMux I__5216 (
            .O(N__30123),
            .I(N__30103));
    InMux I__5215 (
            .O(N__30122),
            .I(N__30103));
    Span4Mux_h I__5214 (
            .O(N__30119),
            .I(N__30100));
    InMux I__5213 (
            .O(N__30118),
            .I(N__30089));
    InMux I__5212 (
            .O(N__30117),
            .I(N__30089));
    InMux I__5211 (
            .O(N__30116),
            .I(N__30089));
    InMux I__5210 (
            .O(N__30115),
            .I(N__30089));
    InMux I__5209 (
            .O(N__30114),
            .I(N__30089));
    LocalMux I__5208 (
            .O(N__30111),
            .I(eis_state_0));
    LocalMux I__5207 (
            .O(N__30108),
            .I(eis_state_0));
    LocalMux I__5206 (
            .O(N__30103),
            .I(eis_state_0));
    Odrv4 I__5205 (
            .O(N__30100),
            .I(eis_state_0));
    LocalMux I__5204 (
            .O(N__30089),
            .I(eis_state_0));
    CascadeMux I__5203 (
            .O(N__30078),
            .I(n11_adj_1621_cascade_));
    CEMux I__5202 (
            .O(N__30075),
            .I(N__30071));
    CEMux I__5201 (
            .O(N__30074),
            .I(N__30068));
    LocalMux I__5200 (
            .O(N__30071),
            .I(N__30065));
    LocalMux I__5199 (
            .O(N__30068),
            .I(N__30062));
    Span4Mux_h I__5198 (
            .O(N__30065),
            .I(N__30059));
    Sp12to4 I__5197 (
            .O(N__30062),
            .I(N__30056));
    Odrv4 I__5196 (
            .O(N__30059),
            .I(n11744));
    Odrv12 I__5195 (
            .O(N__30056),
            .I(n11744));
    InMux I__5194 (
            .O(N__30051),
            .I(N__30045));
    InMux I__5193 (
            .O(N__30050),
            .I(N__30045));
    LocalMux I__5192 (
            .O(N__30045),
            .I(eis_end));
    InMux I__5191 (
            .O(N__30042),
            .I(N__30039));
    LocalMux I__5190 (
            .O(N__30039),
            .I(n26_adj_1530));
    InMux I__5189 (
            .O(N__30036),
            .I(N__30033));
    LocalMux I__5188 (
            .O(N__30033),
            .I(n21234));
    CascadeMux I__5187 (
            .O(N__30030),
            .I(N__30027));
    InMux I__5186 (
            .O(N__30027),
            .I(N__30024));
    LocalMux I__5185 (
            .O(N__30024),
            .I(n21));
    CascadeMux I__5184 (
            .O(N__30021),
            .I(n30_adj_1604_cascade_));
    InMux I__5183 (
            .O(N__30018),
            .I(N__30014));
    InMux I__5182 (
            .O(N__30017),
            .I(N__30011));
    LocalMux I__5181 (
            .O(N__30014),
            .I(n31));
    LocalMux I__5180 (
            .O(N__30011),
            .I(n31));
    CascadeMux I__5179 (
            .O(N__30006),
            .I(N__30003));
    InMux I__5178 (
            .O(N__30003),
            .I(N__29997));
    InMux I__5177 (
            .O(N__30002),
            .I(N__29990));
    InMux I__5176 (
            .O(N__30001),
            .I(N__29987));
    InMux I__5175 (
            .O(N__30000),
            .I(N__29984));
    LocalMux I__5174 (
            .O(N__29997),
            .I(N__29981));
    CascadeMux I__5173 (
            .O(N__29996),
            .I(N__29978));
    CascadeMux I__5172 (
            .O(N__29995),
            .I(N__29975));
    InMux I__5171 (
            .O(N__29994),
            .I(N__29968));
    InMux I__5170 (
            .O(N__29993),
            .I(N__29968));
    LocalMux I__5169 (
            .O(N__29990),
            .I(N__29960));
    LocalMux I__5168 (
            .O(N__29987),
            .I(N__29960));
    LocalMux I__5167 (
            .O(N__29984),
            .I(N__29960));
    Span4Mux_h I__5166 (
            .O(N__29981),
            .I(N__29956));
    InMux I__5165 (
            .O(N__29978),
            .I(N__29953));
    InMux I__5164 (
            .O(N__29975),
            .I(N__29948));
    InMux I__5163 (
            .O(N__29974),
            .I(N__29948));
    InMux I__5162 (
            .O(N__29973),
            .I(N__29945));
    LocalMux I__5161 (
            .O(N__29968),
            .I(N__29942));
    InMux I__5160 (
            .O(N__29967),
            .I(N__29939));
    Span4Mux_v I__5159 (
            .O(N__29960),
            .I(N__29936));
    InMux I__5158 (
            .O(N__29959),
            .I(N__29933));
    Odrv4 I__5157 (
            .O(N__29956),
            .I(DTRIG_N_918));
    LocalMux I__5156 (
            .O(N__29953),
            .I(DTRIG_N_918));
    LocalMux I__5155 (
            .O(N__29948),
            .I(DTRIG_N_918));
    LocalMux I__5154 (
            .O(N__29945),
            .I(DTRIG_N_918));
    Odrv4 I__5153 (
            .O(N__29942),
            .I(DTRIG_N_918));
    LocalMux I__5152 (
            .O(N__29939),
            .I(DTRIG_N_918));
    Odrv4 I__5151 (
            .O(N__29936),
            .I(DTRIG_N_918));
    LocalMux I__5150 (
            .O(N__29933),
            .I(DTRIG_N_918));
    CascadeMux I__5149 (
            .O(N__29916),
            .I(N__29913));
    InMux I__5148 (
            .O(N__29913),
            .I(N__29906));
    InMux I__5147 (
            .O(N__29912),
            .I(N__29903));
    InMux I__5146 (
            .O(N__29911),
            .I(N__29896));
    InMux I__5145 (
            .O(N__29910),
            .I(N__29891));
    InMux I__5144 (
            .O(N__29909),
            .I(N__29891));
    LocalMux I__5143 (
            .O(N__29906),
            .I(N__29887));
    LocalMux I__5142 (
            .O(N__29903),
            .I(N__29884));
    InMux I__5141 (
            .O(N__29902),
            .I(N__29879));
    InMux I__5140 (
            .O(N__29901),
            .I(N__29874));
    InMux I__5139 (
            .O(N__29900),
            .I(N__29874));
    InMux I__5138 (
            .O(N__29899),
            .I(N__29871));
    LocalMux I__5137 (
            .O(N__29896),
            .I(N__29866));
    LocalMux I__5136 (
            .O(N__29891),
            .I(N__29866));
    InMux I__5135 (
            .O(N__29890),
            .I(N__29863));
    Span4Mux_v I__5134 (
            .O(N__29887),
            .I(N__29858));
    Span4Mux_h I__5133 (
            .O(N__29884),
            .I(N__29858));
    InMux I__5132 (
            .O(N__29883),
            .I(N__29853));
    InMux I__5131 (
            .O(N__29882),
            .I(N__29853));
    LocalMux I__5130 (
            .O(N__29879),
            .I(N__29850));
    LocalMux I__5129 (
            .O(N__29874),
            .I(N__29843));
    LocalMux I__5128 (
            .O(N__29871),
            .I(N__29843));
    Span4Mux_v I__5127 (
            .O(N__29866),
            .I(N__29843));
    LocalMux I__5126 (
            .O(N__29863),
            .I(adc_state_1));
    Odrv4 I__5125 (
            .O(N__29858),
            .I(adc_state_1));
    LocalMux I__5124 (
            .O(N__29853),
            .I(adc_state_1));
    Odrv4 I__5123 (
            .O(N__29850),
            .I(adc_state_1));
    Odrv4 I__5122 (
            .O(N__29843),
            .I(adc_state_1));
    CascadeMux I__5121 (
            .O(N__29832),
            .I(n14_adj_1509_cascade_));
    InMux I__5120 (
            .O(N__29829),
            .I(N__29826));
    LocalMux I__5119 (
            .O(N__29826),
            .I(n26_adj_1508));
    InMux I__5118 (
            .O(N__29823),
            .I(N__29820));
    LocalMux I__5117 (
            .O(N__29820),
            .I(n18_adj_1609));
    CascadeMux I__5116 (
            .O(N__29817),
            .I(N__29814));
    InMux I__5115 (
            .O(N__29814),
            .I(N__29811));
    LocalMux I__5114 (
            .O(N__29811),
            .I(\SIG_DDS.tmp_buf_9 ));
    CascadeMux I__5113 (
            .O(N__29808),
            .I(N__29805));
    InMux I__5112 (
            .O(N__29805),
            .I(N__29802));
    LocalMux I__5111 (
            .O(N__29802),
            .I(\SIG_DDS.tmp_buf_5 ));
    InMux I__5110 (
            .O(N__29799),
            .I(N__29793));
    InMux I__5109 (
            .O(N__29798),
            .I(N__29793));
    LocalMux I__5108 (
            .O(N__29793),
            .I(n16554));
    CascadeMux I__5107 (
            .O(N__29790),
            .I(iac_raw_buf_N_736_cascade_));
    InMux I__5106 (
            .O(N__29787),
            .I(N__29784));
    LocalMux I__5105 (
            .O(N__29784),
            .I(n17_adj_1622));
    CascadeMux I__5104 (
            .O(N__29781),
            .I(n20826_cascade_));
    CascadeMux I__5103 (
            .O(N__29778),
            .I(N__29775));
    CascadeBuf I__5102 (
            .O(N__29775),
            .I(N__29772));
    CascadeMux I__5101 (
            .O(N__29772),
            .I(N__29769));
    CascadeBuf I__5100 (
            .O(N__29769),
            .I(N__29766));
    CascadeMux I__5099 (
            .O(N__29766),
            .I(N__29763));
    CascadeBuf I__5098 (
            .O(N__29763),
            .I(N__29760));
    CascadeMux I__5097 (
            .O(N__29760),
            .I(N__29757));
    CascadeBuf I__5096 (
            .O(N__29757),
            .I(N__29754));
    CascadeMux I__5095 (
            .O(N__29754),
            .I(N__29751));
    CascadeBuf I__5094 (
            .O(N__29751),
            .I(N__29748));
    CascadeMux I__5093 (
            .O(N__29748),
            .I(N__29745));
    CascadeBuf I__5092 (
            .O(N__29745),
            .I(N__29742));
    CascadeMux I__5091 (
            .O(N__29742),
            .I(N__29739));
    CascadeBuf I__5090 (
            .O(N__29739),
            .I(N__29736));
    CascadeMux I__5089 (
            .O(N__29736),
            .I(N__29732));
    CascadeMux I__5088 (
            .O(N__29735),
            .I(N__29729));
    CascadeBuf I__5087 (
            .O(N__29732),
            .I(N__29726));
    CascadeBuf I__5086 (
            .O(N__29729),
            .I(N__29723));
    CascadeMux I__5085 (
            .O(N__29726),
            .I(N__29720));
    CascadeMux I__5084 (
            .O(N__29723),
            .I(N__29717));
    CascadeBuf I__5083 (
            .O(N__29720),
            .I(N__29714));
    InMux I__5082 (
            .O(N__29717),
            .I(N__29711));
    CascadeMux I__5081 (
            .O(N__29714),
            .I(N__29708));
    LocalMux I__5080 (
            .O(N__29711),
            .I(N__29705));
    InMux I__5079 (
            .O(N__29708),
            .I(N__29702));
    Sp12to4 I__5078 (
            .O(N__29705),
            .I(N__29698));
    LocalMux I__5077 (
            .O(N__29702),
            .I(N__29695));
    InMux I__5076 (
            .O(N__29701),
            .I(N__29692));
    Span12Mux_h I__5075 (
            .O(N__29698),
            .I(N__29687));
    Span12Mux_h I__5074 (
            .O(N__29695),
            .I(N__29687));
    LocalMux I__5073 (
            .O(N__29692),
            .I(data_count_7));
    Odrv12 I__5072 (
            .O(N__29687),
            .I(data_count_7));
    InMux I__5071 (
            .O(N__29682),
            .I(n19592));
    CascadeMux I__5070 (
            .O(N__29679),
            .I(N__29676));
    CascadeBuf I__5069 (
            .O(N__29676),
            .I(N__29673));
    CascadeMux I__5068 (
            .O(N__29673),
            .I(N__29670));
    CascadeBuf I__5067 (
            .O(N__29670),
            .I(N__29667));
    CascadeMux I__5066 (
            .O(N__29667),
            .I(N__29664));
    CascadeBuf I__5065 (
            .O(N__29664),
            .I(N__29661));
    CascadeMux I__5064 (
            .O(N__29661),
            .I(N__29658));
    CascadeBuf I__5063 (
            .O(N__29658),
            .I(N__29655));
    CascadeMux I__5062 (
            .O(N__29655),
            .I(N__29652));
    CascadeBuf I__5061 (
            .O(N__29652),
            .I(N__29649));
    CascadeMux I__5060 (
            .O(N__29649),
            .I(N__29646));
    CascadeBuf I__5059 (
            .O(N__29646),
            .I(N__29643));
    CascadeMux I__5058 (
            .O(N__29643),
            .I(N__29640));
    CascadeBuf I__5057 (
            .O(N__29640),
            .I(N__29637));
    CascadeMux I__5056 (
            .O(N__29637),
            .I(N__29634));
    CascadeBuf I__5055 (
            .O(N__29634),
            .I(N__29630));
    CascadeMux I__5054 (
            .O(N__29633),
            .I(N__29627));
    CascadeMux I__5053 (
            .O(N__29630),
            .I(N__29624));
    CascadeBuf I__5052 (
            .O(N__29627),
            .I(N__29621));
    CascadeBuf I__5051 (
            .O(N__29624),
            .I(N__29618));
    CascadeMux I__5050 (
            .O(N__29621),
            .I(N__29615));
    CascadeMux I__5049 (
            .O(N__29618),
            .I(N__29612));
    InMux I__5048 (
            .O(N__29615),
            .I(N__29609));
    InMux I__5047 (
            .O(N__29612),
            .I(N__29606));
    LocalMux I__5046 (
            .O(N__29609),
            .I(N__29603));
    LocalMux I__5045 (
            .O(N__29606),
            .I(N__29600));
    Span4Mux_h I__5044 (
            .O(N__29603),
            .I(N__29597));
    Span4Mux_v I__5043 (
            .O(N__29600),
            .I(N__29594));
    Span4Mux_h I__5042 (
            .O(N__29597),
            .I(N__29590));
    Sp12to4 I__5041 (
            .O(N__29594),
            .I(N__29587));
    InMux I__5040 (
            .O(N__29593),
            .I(N__29584));
    Sp12to4 I__5039 (
            .O(N__29590),
            .I(N__29579));
    Span12Mux_h I__5038 (
            .O(N__29587),
            .I(N__29579));
    LocalMux I__5037 (
            .O(N__29584),
            .I(data_count_8));
    Odrv12 I__5036 (
            .O(N__29579),
            .I(data_count_8));
    InMux I__5035 (
            .O(N__29574),
            .I(bfn_11_14_0_));
    InMux I__5034 (
            .O(N__29571),
            .I(n19594));
    CascadeMux I__5033 (
            .O(N__29568),
            .I(N__29565));
    CascadeBuf I__5032 (
            .O(N__29565),
            .I(N__29562));
    CascadeMux I__5031 (
            .O(N__29562),
            .I(N__29559));
    CascadeBuf I__5030 (
            .O(N__29559),
            .I(N__29556));
    CascadeMux I__5029 (
            .O(N__29556),
            .I(N__29553));
    CascadeBuf I__5028 (
            .O(N__29553),
            .I(N__29550));
    CascadeMux I__5027 (
            .O(N__29550),
            .I(N__29547));
    CascadeBuf I__5026 (
            .O(N__29547),
            .I(N__29544));
    CascadeMux I__5025 (
            .O(N__29544),
            .I(N__29541));
    CascadeBuf I__5024 (
            .O(N__29541),
            .I(N__29538));
    CascadeMux I__5023 (
            .O(N__29538),
            .I(N__29535));
    CascadeBuf I__5022 (
            .O(N__29535),
            .I(N__29532));
    CascadeMux I__5021 (
            .O(N__29532),
            .I(N__29529));
    CascadeBuf I__5020 (
            .O(N__29529),
            .I(N__29526));
    CascadeMux I__5019 (
            .O(N__29526),
            .I(N__29523));
    CascadeBuf I__5018 (
            .O(N__29523),
            .I(N__29519));
    CascadeMux I__5017 (
            .O(N__29522),
            .I(N__29516));
    CascadeMux I__5016 (
            .O(N__29519),
            .I(N__29513));
    CascadeBuf I__5015 (
            .O(N__29516),
            .I(N__29510));
    CascadeBuf I__5014 (
            .O(N__29513),
            .I(N__29507));
    CascadeMux I__5013 (
            .O(N__29510),
            .I(N__29504));
    CascadeMux I__5012 (
            .O(N__29507),
            .I(N__29501));
    InMux I__5011 (
            .O(N__29504),
            .I(N__29498));
    InMux I__5010 (
            .O(N__29501),
            .I(N__29495));
    LocalMux I__5009 (
            .O(N__29498),
            .I(N__29492));
    LocalMux I__5008 (
            .O(N__29495),
            .I(N__29489));
    Span4Mux_v I__5007 (
            .O(N__29492),
            .I(N__29486));
    Span4Mux_v I__5006 (
            .O(N__29489),
            .I(N__29483));
    Sp12to4 I__5005 (
            .O(N__29486),
            .I(N__29479));
    Sp12to4 I__5004 (
            .O(N__29483),
            .I(N__29476));
    InMux I__5003 (
            .O(N__29482),
            .I(N__29473));
    Span12Mux_h I__5002 (
            .O(N__29479),
            .I(N__29468));
    Span12Mux_h I__5001 (
            .O(N__29476),
            .I(N__29468));
    LocalMux I__5000 (
            .O(N__29473),
            .I(data_count_9));
    Odrv12 I__4999 (
            .O(N__29468),
            .I(data_count_9));
    CascadeMux I__4998 (
            .O(N__29463),
            .I(N__29460));
    InMux I__4997 (
            .O(N__29460),
            .I(N__29457));
    LocalMux I__4996 (
            .O(N__29457),
            .I(\SIG_DDS.tmp_buf_10 ));
    CascadeMux I__4995 (
            .O(N__29454),
            .I(N__29450));
    InMux I__4994 (
            .O(N__29453),
            .I(N__29446));
    InMux I__4993 (
            .O(N__29450),
            .I(N__29441));
    InMux I__4992 (
            .O(N__29449),
            .I(N__29441));
    LocalMux I__4991 (
            .O(N__29446),
            .I(buf_dds0_5));
    LocalMux I__4990 (
            .O(N__29441),
            .I(buf_dds0_5));
    CascadeMux I__4989 (
            .O(N__29436),
            .I(N__29433));
    InMux I__4988 (
            .O(N__29433),
            .I(N__29430));
    LocalMux I__4987 (
            .O(N__29430),
            .I(N__29425));
    InMux I__4986 (
            .O(N__29429),
            .I(N__29420));
    InMux I__4985 (
            .O(N__29428),
            .I(N__29420));
    Odrv12 I__4984 (
            .O(N__29425),
            .I(buf_dds0_14));
    LocalMux I__4983 (
            .O(N__29420),
            .I(buf_dds0_14));
    InMux I__4982 (
            .O(N__29415),
            .I(N__29412));
    LocalMux I__4981 (
            .O(N__29412),
            .I(\SIG_DDS.tmp_buf_13 ));
    CascadeMux I__4980 (
            .O(N__29409),
            .I(N__29406));
    InMux I__4979 (
            .O(N__29406),
            .I(N__29403));
    LocalMux I__4978 (
            .O(N__29403),
            .I(\SIG_DDS.tmp_buf_11 ));
    CascadeMux I__4977 (
            .O(N__29400),
            .I(N__29397));
    InMux I__4976 (
            .O(N__29397),
            .I(N__29394));
    LocalMux I__4975 (
            .O(N__29394),
            .I(\SIG_DDS.tmp_buf_12 ));
    InMux I__4974 (
            .O(N__29391),
            .I(N__29388));
    LocalMux I__4973 (
            .O(N__29388),
            .I(\CLK_DDS.tmp_buf_8 ));
    CascadeMux I__4972 (
            .O(N__29385),
            .I(N__29382));
    InMux I__4971 (
            .O(N__29382),
            .I(N__29379));
    LocalMux I__4970 (
            .O(N__29379),
            .I(\CLK_DDS.tmp_buf_9 ));
    CascadeMux I__4969 (
            .O(N__29376),
            .I(N__29373));
    CascadeBuf I__4968 (
            .O(N__29373),
            .I(N__29370));
    CascadeMux I__4967 (
            .O(N__29370),
            .I(N__29367));
    CascadeBuf I__4966 (
            .O(N__29367),
            .I(N__29364));
    CascadeMux I__4965 (
            .O(N__29364),
            .I(N__29361));
    CascadeBuf I__4964 (
            .O(N__29361),
            .I(N__29358));
    CascadeMux I__4963 (
            .O(N__29358),
            .I(N__29355));
    CascadeBuf I__4962 (
            .O(N__29355),
            .I(N__29352));
    CascadeMux I__4961 (
            .O(N__29352),
            .I(N__29349));
    CascadeBuf I__4960 (
            .O(N__29349),
            .I(N__29346));
    CascadeMux I__4959 (
            .O(N__29346),
            .I(N__29343));
    CascadeBuf I__4958 (
            .O(N__29343),
            .I(N__29340));
    CascadeMux I__4957 (
            .O(N__29340),
            .I(N__29337));
    CascadeBuf I__4956 (
            .O(N__29337),
            .I(N__29334));
    CascadeMux I__4955 (
            .O(N__29334),
            .I(N__29331));
    CascadeBuf I__4954 (
            .O(N__29331),
            .I(N__29328));
    CascadeMux I__4953 (
            .O(N__29328),
            .I(N__29324));
    CascadeMux I__4952 (
            .O(N__29327),
            .I(N__29321));
    CascadeBuf I__4951 (
            .O(N__29324),
            .I(N__29318));
    CascadeBuf I__4950 (
            .O(N__29321),
            .I(N__29315));
    CascadeMux I__4949 (
            .O(N__29318),
            .I(N__29312));
    CascadeMux I__4948 (
            .O(N__29315),
            .I(N__29309));
    InMux I__4947 (
            .O(N__29312),
            .I(N__29306));
    InMux I__4946 (
            .O(N__29309),
            .I(N__29303));
    LocalMux I__4945 (
            .O(N__29306),
            .I(N__29300));
    LocalMux I__4944 (
            .O(N__29303),
            .I(N__29297));
    Span4Mux_v I__4943 (
            .O(N__29300),
            .I(N__29294));
    Span4Mux_v I__4942 (
            .O(N__29297),
            .I(N__29290));
    Span4Mux_h I__4941 (
            .O(N__29294),
            .I(N__29287));
    CascadeMux I__4940 (
            .O(N__29293),
            .I(N__29284));
    Span4Mux_v I__4939 (
            .O(N__29290),
            .I(N__29281));
    Span4Mux_h I__4938 (
            .O(N__29287),
            .I(N__29278));
    InMux I__4937 (
            .O(N__29284),
            .I(N__29275));
    Span4Mux_h I__4936 (
            .O(N__29281),
            .I(N__29270));
    Span4Mux_v I__4935 (
            .O(N__29278),
            .I(N__29270));
    LocalMux I__4934 (
            .O(N__29275),
            .I(data_count_0));
    Odrv4 I__4933 (
            .O(N__29270),
            .I(data_count_0));
    CascadeMux I__4932 (
            .O(N__29265),
            .I(N__29262));
    CascadeBuf I__4931 (
            .O(N__29262),
            .I(N__29259));
    CascadeMux I__4930 (
            .O(N__29259),
            .I(N__29256));
    CascadeBuf I__4929 (
            .O(N__29256),
            .I(N__29253));
    CascadeMux I__4928 (
            .O(N__29253),
            .I(N__29250));
    CascadeBuf I__4927 (
            .O(N__29250),
            .I(N__29247));
    CascadeMux I__4926 (
            .O(N__29247),
            .I(N__29244));
    CascadeBuf I__4925 (
            .O(N__29244),
            .I(N__29241));
    CascadeMux I__4924 (
            .O(N__29241),
            .I(N__29238));
    CascadeBuf I__4923 (
            .O(N__29238),
            .I(N__29235));
    CascadeMux I__4922 (
            .O(N__29235),
            .I(N__29232));
    CascadeBuf I__4921 (
            .O(N__29232),
            .I(N__29229));
    CascadeMux I__4920 (
            .O(N__29229),
            .I(N__29226));
    CascadeBuf I__4919 (
            .O(N__29226),
            .I(N__29223));
    CascadeMux I__4918 (
            .O(N__29223),
            .I(N__29220));
    CascadeBuf I__4917 (
            .O(N__29220),
            .I(N__29216));
    CascadeMux I__4916 (
            .O(N__29219),
            .I(N__29213));
    CascadeMux I__4915 (
            .O(N__29216),
            .I(N__29210));
    CascadeBuf I__4914 (
            .O(N__29213),
            .I(N__29207));
    CascadeBuf I__4913 (
            .O(N__29210),
            .I(N__29204));
    CascadeMux I__4912 (
            .O(N__29207),
            .I(N__29201));
    CascadeMux I__4911 (
            .O(N__29204),
            .I(N__29198));
    InMux I__4910 (
            .O(N__29201),
            .I(N__29195));
    InMux I__4909 (
            .O(N__29198),
            .I(N__29192));
    LocalMux I__4908 (
            .O(N__29195),
            .I(N__29189));
    LocalMux I__4907 (
            .O(N__29192),
            .I(N__29186));
    Span4Mux_h I__4906 (
            .O(N__29189),
            .I(N__29183));
    Span4Mux_h I__4905 (
            .O(N__29186),
            .I(N__29180));
    Sp12to4 I__4904 (
            .O(N__29183),
            .I(N__29176));
    Sp12to4 I__4903 (
            .O(N__29180),
            .I(N__29173));
    InMux I__4902 (
            .O(N__29179),
            .I(N__29170));
    Span12Mux_v I__4901 (
            .O(N__29176),
            .I(N__29165));
    Span12Mux_v I__4900 (
            .O(N__29173),
            .I(N__29165));
    LocalMux I__4899 (
            .O(N__29170),
            .I(data_count_1));
    Odrv12 I__4898 (
            .O(N__29165),
            .I(data_count_1));
    InMux I__4897 (
            .O(N__29160),
            .I(n19586));
    CascadeMux I__4896 (
            .O(N__29157),
            .I(N__29154));
    CascadeBuf I__4895 (
            .O(N__29154),
            .I(N__29151));
    CascadeMux I__4894 (
            .O(N__29151),
            .I(N__29148));
    CascadeBuf I__4893 (
            .O(N__29148),
            .I(N__29145));
    CascadeMux I__4892 (
            .O(N__29145),
            .I(N__29142));
    CascadeBuf I__4891 (
            .O(N__29142),
            .I(N__29139));
    CascadeMux I__4890 (
            .O(N__29139),
            .I(N__29136));
    CascadeBuf I__4889 (
            .O(N__29136),
            .I(N__29133));
    CascadeMux I__4888 (
            .O(N__29133),
            .I(N__29130));
    CascadeBuf I__4887 (
            .O(N__29130),
            .I(N__29127));
    CascadeMux I__4886 (
            .O(N__29127),
            .I(N__29124));
    CascadeBuf I__4885 (
            .O(N__29124),
            .I(N__29121));
    CascadeMux I__4884 (
            .O(N__29121),
            .I(N__29118));
    CascadeBuf I__4883 (
            .O(N__29118),
            .I(N__29115));
    CascadeMux I__4882 (
            .O(N__29115),
            .I(N__29112));
    CascadeBuf I__4881 (
            .O(N__29112),
            .I(N__29109));
    CascadeMux I__4880 (
            .O(N__29109),
            .I(N__29105));
    CascadeMux I__4879 (
            .O(N__29108),
            .I(N__29102));
    CascadeBuf I__4878 (
            .O(N__29105),
            .I(N__29099));
    CascadeBuf I__4877 (
            .O(N__29102),
            .I(N__29096));
    CascadeMux I__4876 (
            .O(N__29099),
            .I(N__29093));
    CascadeMux I__4875 (
            .O(N__29096),
            .I(N__29090));
    InMux I__4874 (
            .O(N__29093),
            .I(N__29087));
    InMux I__4873 (
            .O(N__29090),
            .I(N__29084));
    LocalMux I__4872 (
            .O(N__29087),
            .I(N__29081));
    LocalMux I__4871 (
            .O(N__29084),
            .I(N__29078));
    Span4Mux_v I__4870 (
            .O(N__29081),
            .I(N__29075));
    Sp12to4 I__4869 (
            .O(N__29078),
            .I(N__29071));
    Sp12to4 I__4868 (
            .O(N__29075),
            .I(N__29068));
    InMux I__4867 (
            .O(N__29074),
            .I(N__29065));
    Span12Mux_v I__4866 (
            .O(N__29071),
            .I(N__29062));
    Span12Mux_h I__4865 (
            .O(N__29068),
            .I(N__29059));
    LocalMux I__4864 (
            .O(N__29065),
            .I(data_count_2));
    Odrv12 I__4863 (
            .O(N__29062),
            .I(data_count_2));
    Odrv12 I__4862 (
            .O(N__29059),
            .I(data_count_2));
    InMux I__4861 (
            .O(N__29052),
            .I(n19587));
    CascadeMux I__4860 (
            .O(N__29049),
            .I(N__29046));
    CascadeBuf I__4859 (
            .O(N__29046),
            .I(N__29043));
    CascadeMux I__4858 (
            .O(N__29043),
            .I(N__29040));
    CascadeBuf I__4857 (
            .O(N__29040),
            .I(N__29037));
    CascadeMux I__4856 (
            .O(N__29037),
            .I(N__29034));
    CascadeBuf I__4855 (
            .O(N__29034),
            .I(N__29031));
    CascadeMux I__4854 (
            .O(N__29031),
            .I(N__29028));
    CascadeBuf I__4853 (
            .O(N__29028),
            .I(N__29025));
    CascadeMux I__4852 (
            .O(N__29025),
            .I(N__29022));
    CascadeBuf I__4851 (
            .O(N__29022),
            .I(N__29019));
    CascadeMux I__4850 (
            .O(N__29019),
            .I(N__29016));
    CascadeBuf I__4849 (
            .O(N__29016),
            .I(N__29013));
    CascadeMux I__4848 (
            .O(N__29013),
            .I(N__29010));
    CascadeBuf I__4847 (
            .O(N__29010),
            .I(N__29007));
    CascadeMux I__4846 (
            .O(N__29007),
            .I(N__29004));
    CascadeBuf I__4845 (
            .O(N__29004),
            .I(N__29001));
    CascadeMux I__4844 (
            .O(N__29001),
            .I(N__28998));
    CascadeBuf I__4843 (
            .O(N__28998),
            .I(N__28994));
    CascadeMux I__4842 (
            .O(N__28997),
            .I(N__28991));
    CascadeMux I__4841 (
            .O(N__28994),
            .I(N__28988));
    CascadeBuf I__4840 (
            .O(N__28991),
            .I(N__28985));
    InMux I__4839 (
            .O(N__28988),
            .I(N__28982));
    CascadeMux I__4838 (
            .O(N__28985),
            .I(N__28979));
    LocalMux I__4837 (
            .O(N__28982),
            .I(N__28976));
    InMux I__4836 (
            .O(N__28979),
            .I(N__28973));
    Span4Mux_v I__4835 (
            .O(N__28976),
            .I(N__28970));
    LocalMux I__4834 (
            .O(N__28973),
            .I(N__28966));
    Sp12to4 I__4833 (
            .O(N__28970),
            .I(N__28963));
    InMux I__4832 (
            .O(N__28969),
            .I(N__28960));
    Span12Mux_v I__4831 (
            .O(N__28966),
            .I(N__28957));
    Span12Mux_h I__4830 (
            .O(N__28963),
            .I(N__28954));
    LocalMux I__4829 (
            .O(N__28960),
            .I(data_count_3));
    Odrv12 I__4828 (
            .O(N__28957),
            .I(data_count_3));
    Odrv12 I__4827 (
            .O(N__28954),
            .I(data_count_3));
    InMux I__4826 (
            .O(N__28947),
            .I(n19588));
    CascadeMux I__4825 (
            .O(N__28944),
            .I(N__28941));
    CascadeBuf I__4824 (
            .O(N__28941),
            .I(N__28938));
    CascadeMux I__4823 (
            .O(N__28938),
            .I(N__28935));
    CascadeBuf I__4822 (
            .O(N__28935),
            .I(N__28932));
    CascadeMux I__4821 (
            .O(N__28932),
            .I(N__28929));
    CascadeBuf I__4820 (
            .O(N__28929),
            .I(N__28926));
    CascadeMux I__4819 (
            .O(N__28926),
            .I(N__28923));
    CascadeBuf I__4818 (
            .O(N__28923),
            .I(N__28920));
    CascadeMux I__4817 (
            .O(N__28920),
            .I(N__28917));
    CascadeBuf I__4816 (
            .O(N__28917),
            .I(N__28914));
    CascadeMux I__4815 (
            .O(N__28914),
            .I(N__28911));
    CascadeBuf I__4814 (
            .O(N__28911),
            .I(N__28908));
    CascadeMux I__4813 (
            .O(N__28908),
            .I(N__28905));
    CascadeBuf I__4812 (
            .O(N__28905),
            .I(N__28902));
    CascadeMux I__4811 (
            .O(N__28902),
            .I(N__28899));
    CascadeBuf I__4810 (
            .O(N__28899),
            .I(N__28895));
    CascadeMux I__4809 (
            .O(N__28898),
            .I(N__28892));
    CascadeMux I__4808 (
            .O(N__28895),
            .I(N__28889));
    CascadeBuf I__4807 (
            .O(N__28892),
            .I(N__28886));
    CascadeBuf I__4806 (
            .O(N__28889),
            .I(N__28883));
    CascadeMux I__4805 (
            .O(N__28886),
            .I(N__28880));
    CascadeMux I__4804 (
            .O(N__28883),
            .I(N__28877));
    InMux I__4803 (
            .O(N__28880),
            .I(N__28874));
    InMux I__4802 (
            .O(N__28877),
            .I(N__28871));
    LocalMux I__4801 (
            .O(N__28874),
            .I(N__28868));
    LocalMux I__4800 (
            .O(N__28871),
            .I(N__28865));
    Span4Mux_h I__4799 (
            .O(N__28868),
            .I(N__28862));
    Span4Mux_v I__4798 (
            .O(N__28865),
            .I(N__28859));
    Span4Mux_v I__4797 (
            .O(N__28862),
            .I(N__28855));
    Span4Mux_v I__4796 (
            .O(N__28859),
            .I(N__28852));
    InMux I__4795 (
            .O(N__28858),
            .I(N__28849));
    Span4Mux_h I__4794 (
            .O(N__28855),
            .I(N__28846));
    Sp12to4 I__4793 (
            .O(N__28852),
            .I(N__28843));
    LocalMux I__4792 (
            .O(N__28849),
            .I(data_count_4));
    Odrv4 I__4791 (
            .O(N__28846),
            .I(data_count_4));
    Odrv12 I__4790 (
            .O(N__28843),
            .I(data_count_4));
    InMux I__4789 (
            .O(N__28836),
            .I(n19589));
    CascadeMux I__4788 (
            .O(N__28833),
            .I(N__28830));
    CascadeBuf I__4787 (
            .O(N__28830),
            .I(N__28827));
    CascadeMux I__4786 (
            .O(N__28827),
            .I(N__28824));
    CascadeBuf I__4785 (
            .O(N__28824),
            .I(N__28821));
    CascadeMux I__4784 (
            .O(N__28821),
            .I(N__28818));
    CascadeBuf I__4783 (
            .O(N__28818),
            .I(N__28815));
    CascadeMux I__4782 (
            .O(N__28815),
            .I(N__28812));
    CascadeBuf I__4781 (
            .O(N__28812),
            .I(N__28809));
    CascadeMux I__4780 (
            .O(N__28809),
            .I(N__28806));
    CascadeBuf I__4779 (
            .O(N__28806),
            .I(N__28803));
    CascadeMux I__4778 (
            .O(N__28803),
            .I(N__28800));
    CascadeBuf I__4777 (
            .O(N__28800),
            .I(N__28797));
    CascadeMux I__4776 (
            .O(N__28797),
            .I(N__28794));
    CascadeBuf I__4775 (
            .O(N__28794),
            .I(N__28791));
    CascadeMux I__4774 (
            .O(N__28791),
            .I(N__28787));
    CascadeMux I__4773 (
            .O(N__28790),
            .I(N__28784));
    CascadeBuf I__4772 (
            .O(N__28787),
            .I(N__28781));
    CascadeBuf I__4771 (
            .O(N__28784),
            .I(N__28778));
    CascadeMux I__4770 (
            .O(N__28781),
            .I(N__28775));
    CascadeMux I__4769 (
            .O(N__28778),
            .I(N__28772));
    CascadeBuf I__4768 (
            .O(N__28775),
            .I(N__28769));
    InMux I__4767 (
            .O(N__28772),
            .I(N__28766));
    CascadeMux I__4766 (
            .O(N__28769),
            .I(N__28763));
    LocalMux I__4765 (
            .O(N__28766),
            .I(N__28760));
    InMux I__4764 (
            .O(N__28763),
            .I(N__28757));
    Span4Mux_h I__4763 (
            .O(N__28760),
            .I(N__28754));
    LocalMux I__4762 (
            .O(N__28757),
            .I(N__28750));
    Span4Mux_v I__4761 (
            .O(N__28754),
            .I(N__28747));
    InMux I__4760 (
            .O(N__28753),
            .I(N__28744));
    Sp12to4 I__4759 (
            .O(N__28750),
            .I(N__28741));
    Span4Mux_h I__4758 (
            .O(N__28747),
            .I(N__28738));
    LocalMux I__4757 (
            .O(N__28744),
            .I(N__28733));
    Span12Mux_v I__4756 (
            .O(N__28741),
            .I(N__28733));
    Odrv4 I__4755 (
            .O(N__28738),
            .I(data_count_5));
    Odrv12 I__4754 (
            .O(N__28733),
            .I(data_count_5));
    InMux I__4753 (
            .O(N__28728),
            .I(n19590));
    CascadeMux I__4752 (
            .O(N__28725),
            .I(N__28722));
    CascadeBuf I__4751 (
            .O(N__28722),
            .I(N__28719));
    CascadeMux I__4750 (
            .O(N__28719),
            .I(N__28716));
    CascadeBuf I__4749 (
            .O(N__28716),
            .I(N__28713));
    CascadeMux I__4748 (
            .O(N__28713),
            .I(N__28710));
    CascadeBuf I__4747 (
            .O(N__28710),
            .I(N__28707));
    CascadeMux I__4746 (
            .O(N__28707),
            .I(N__28704));
    CascadeBuf I__4745 (
            .O(N__28704),
            .I(N__28701));
    CascadeMux I__4744 (
            .O(N__28701),
            .I(N__28698));
    CascadeBuf I__4743 (
            .O(N__28698),
            .I(N__28695));
    CascadeMux I__4742 (
            .O(N__28695),
            .I(N__28692));
    CascadeBuf I__4741 (
            .O(N__28692),
            .I(N__28689));
    CascadeMux I__4740 (
            .O(N__28689),
            .I(N__28686));
    CascadeBuf I__4739 (
            .O(N__28686),
            .I(N__28682));
    CascadeMux I__4738 (
            .O(N__28685),
            .I(N__28679));
    CascadeMux I__4737 (
            .O(N__28682),
            .I(N__28676));
    CascadeBuf I__4736 (
            .O(N__28679),
            .I(N__28673));
    CascadeBuf I__4735 (
            .O(N__28676),
            .I(N__28670));
    CascadeMux I__4734 (
            .O(N__28673),
            .I(N__28667));
    CascadeMux I__4733 (
            .O(N__28670),
            .I(N__28664));
    InMux I__4732 (
            .O(N__28667),
            .I(N__28661));
    CascadeBuf I__4731 (
            .O(N__28664),
            .I(N__28658));
    LocalMux I__4730 (
            .O(N__28661),
            .I(N__28655));
    CascadeMux I__4729 (
            .O(N__28658),
            .I(N__28652));
    Span4Mux_v I__4728 (
            .O(N__28655),
            .I(N__28649));
    InMux I__4727 (
            .O(N__28652),
            .I(N__28646));
    Span4Mux_v I__4726 (
            .O(N__28649),
            .I(N__28642));
    LocalMux I__4725 (
            .O(N__28646),
            .I(N__28639));
    InMux I__4724 (
            .O(N__28645),
            .I(N__28636));
    Span4Mux_h I__4723 (
            .O(N__28642),
            .I(N__28633));
    Span12Mux_v I__4722 (
            .O(N__28639),
            .I(N__28630));
    LocalMux I__4721 (
            .O(N__28636),
            .I(data_count_6));
    Odrv4 I__4720 (
            .O(N__28633),
            .I(data_count_6));
    Odrv12 I__4719 (
            .O(N__28630),
            .I(data_count_6));
    InMux I__4718 (
            .O(N__28623),
            .I(n19591));
    InMux I__4717 (
            .O(N__28620),
            .I(n19770));
    InMux I__4716 (
            .O(N__28617),
            .I(n19771));
    CascadeMux I__4715 (
            .O(N__28614),
            .I(N__28611));
    InMux I__4714 (
            .O(N__28611),
            .I(N__28608));
    LocalMux I__4713 (
            .O(N__28608),
            .I(N__28603));
    InMux I__4712 (
            .O(N__28607),
            .I(N__28600));
    InMux I__4711 (
            .O(N__28606),
            .I(N__28597));
    Span4Mux_h I__4710 (
            .O(N__28603),
            .I(N__28594));
    LocalMux I__4709 (
            .O(N__28600),
            .I(N__28591));
    LocalMux I__4708 (
            .O(N__28597),
            .I(buf_dds1_14));
    Odrv4 I__4707 (
            .O(N__28594),
            .I(buf_dds1_14));
    Odrv4 I__4706 (
            .O(N__28591),
            .I(buf_dds1_14));
    InMux I__4705 (
            .O(N__28584),
            .I(N__28581));
    LocalMux I__4704 (
            .O(N__28581),
            .I(\CLK_DDS.tmp_buf_13 ));
    CascadeMux I__4703 (
            .O(N__28578),
            .I(N__28575));
    InMux I__4702 (
            .O(N__28575),
            .I(N__28572));
    LocalMux I__4701 (
            .O(N__28572),
            .I(\CLK_DDS.tmp_buf_14 ));
    InMux I__4700 (
            .O(N__28569),
            .I(N__28566));
    LocalMux I__4699 (
            .O(N__28566),
            .I(\CLK_DDS.tmp_buf_0 ));
    CascadeMux I__4698 (
            .O(N__28563),
            .I(N__28560));
    InMux I__4697 (
            .O(N__28560),
            .I(N__28557));
    LocalMux I__4696 (
            .O(N__28557),
            .I(\CLK_DDS.tmp_buf_1 ));
    CascadeMux I__4695 (
            .O(N__28554),
            .I(N__28551));
    InMux I__4694 (
            .O(N__28551),
            .I(N__28548));
    LocalMux I__4693 (
            .O(N__28548),
            .I(\CLK_DDS.tmp_buf_2 ));
    CascadeMux I__4692 (
            .O(N__28545),
            .I(N__28542));
    InMux I__4691 (
            .O(N__28542),
            .I(N__28539));
    LocalMux I__4690 (
            .O(N__28539),
            .I(\CLK_DDS.tmp_buf_3 ));
    CascadeMux I__4689 (
            .O(N__28536),
            .I(N__28533));
    InMux I__4688 (
            .O(N__28533),
            .I(N__28530));
    LocalMux I__4687 (
            .O(N__28530),
            .I(\CLK_DDS.tmp_buf_4 ));
    CascadeMux I__4686 (
            .O(N__28527),
            .I(N__28524));
    InMux I__4685 (
            .O(N__28524),
            .I(N__28521));
    LocalMux I__4684 (
            .O(N__28521),
            .I(\CLK_DDS.tmp_buf_5 ));
    InMux I__4683 (
            .O(N__28518),
            .I(N__28515));
    LocalMux I__4682 (
            .O(N__28515),
            .I(\CLK_DDS.tmp_buf_6 ));
    InMux I__4681 (
            .O(N__28512),
            .I(n19761));
    InMux I__4680 (
            .O(N__28509),
            .I(n19762));
    InMux I__4679 (
            .O(N__28506),
            .I(n19763));
    InMux I__4678 (
            .O(N__28503),
            .I(n19764));
    InMux I__4677 (
            .O(N__28500),
            .I(bfn_11_11_0_));
    InMux I__4676 (
            .O(N__28497),
            .I(n19766));
    InMux I__4675 (
            .O(N__28494),
            .I(n19767));
    InMux I__4674 (
            .O(N__28491),
            .I(n19768));
    InMux I__4673 (
            .O(N__28488),
            .I(n19769));
    InMux I__4672 (
            .O(N__28485),
            .I(n19752));
    InMux I__4671 (
            .O(N__28482),
            .I(n19753));
    InMux I__4670 (
            .O(N__28479),
            .I(n19754));
    InMux I__4669 (
            .O(N__28476),
            .I(n19755));
    InMux I__4668 (
            .O(N__28473),
            .I(n19756));
    InMux I__4667 (
            .O(N__28470),
            .I(bfn_11_10_0_));
    InMux I__4666 (
            .O(N__28467),
            .I(n19758));
    InMux I__4665 (
            .O(N__28464),
            .I(n19759));
    InMux I__4664 (
            .O(N__28461),
            .I(n19760));
    InMux I__4663 (
            .O(N__28458),
            .I(N__28448));
    InMux I__4662 (
            .O(N__28457),
            .I(N__28448));
    InMux I__4661 (
            .O(N__28456),
            .I(N__28448));
    InMux I__4660 (
            .O(N__28455),
            .I(N__28445));
    LocalMux I__4659 (
            .O(N__28448),
            .I(\comm_spi.bit_cnt_1 ));
    LocalMux I__4658 (
            .O(N__28445),
            .I(\comm_spi.bit_cnt_1 ));
    CascadeMux I__4657 (
            .O(N__28440),
            .I(N__28435));
    InMux I__4656 (
            .O(N__28439),
            .I(N__28430));
    InMux I__4655 (
            .O(N__28438),
            .I(N__28430));
    InMux I__4654 (
            .O(N__28435),
            .I(N__28427));
    LocalMux I__4653 (
            .O(N__28430),
            .I(\comm_spi.bit_cnt_2 ));
    LocalMux I__4652 (
            .O(N__28427),
            .I(\comm_spi.bit_cnt_2 ));
    CascadeMux I__4651 (
            .O(N__28422),
            .I(N__28419));
    InMux I__4650 (
            .O(N__28419),
            .I(N__28406));
    InMux I__4649 (
            .O(N__28418),
            .I(N__28406));
    InMux I__4648 (
            .O(N__28417),
            .I(N__28406));
    InMux I__4647 (
            .O(N__28416),
            .I(N__28406));
    InMux I__4646 (
            .O(N__28415),
            .I(N__28403));
    LocalMux I__4645 (
            .O(N__28406),
            .I(\comm_spi.bit_cnt_0 ));
    LocalMux I__4644 (
            .O(N__28403),
            .I(\comm_spi.bit_cnt_0 ));
    CascadeMux I__4643 (
            .O(N__28398),
            .I(N__28394));
    CascadeMux I__4642 (
            .O(N__28397),
            .I(N__28391));
    InMux I__4641 (
            .O(N__28394),
            .I(N__28388));
    InMux I__4640 (
            .O(N__28391),
            .I(N__28384));
    LocalMux I__4639 (
            .O(N__28388),
            .I(N__28381));
    InMux I__4638 (
            .O(N__28387),
            .I(N__28378));
    LocalMux I__4637 (
            .O(N__28384),
            .I(cmd_rdadctmp_11));
    Odrv12 I__4636 (
            .O(N__28381),
            .I(cmd_rdadctmp_11));
    LocalMux I__4635 (
            .O(N__28378),
            .I(cmd_rdadctmp_11));
    InMux I__4634 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__4633 (
            .O(N__28368),
            .I(N__28365));
    Span4Mux_v I__4632 (
            .O(N__28365),
            .I(N__28362));
    Sp12to4 I__4631 (
            .O(N__28362),
            .I(N__28357));
    InMux I__4630 (
            .O(N__28361),
            .I(N__28352));
    InMux I__4629 (
            .O(N__28360),
            .I(N__28352));
    Odrv12 I__4628 (
            .O(N__28357),
            .I(buf_adcdata_vac_3));
    LocalMux I__4627 (
            .O(N__28352),
            .I(buf_adcdata_vac_3));
    InMux I__4626 (
            .O(N__28347),
            .I(N__28343));
    CascadeMux I__4625 (
            .O(N__28346),
            .I(N__28340));
    LocalMux I__4624 (
            .O(N__28343),
            .I(N__28337));
    InMux I__4623 (
            .O(N__28340),
            .I(N__28334));
    Span4Mux_v I__4622 (
            .O(N__28337),
            .I(N__28328));
    LocalMux I__4621 (
            .O(N__28334),
            .I(N__28328));
    CascadeMux I__4620 (
            .O(N__28333),
            .I(N__28325));
    Span4Mux_h I__4619 (
            .O(N__28328),
            .I(N__28322));
    InMux I__4618 (
            .O(N__28325),
            .I(N__28319));
    Odrv4 I__4617 (
            .O(N__28322),
            .I(cmd_rdadctmp_10_adj_1440));
    LocalMux I__4616 (
            .O(N__28319),
            .I(cmd_rdadctmp_10_adj_1440));
    CascadeMux I__4615 (
            .O(N__28314),
            .I(N__28310));
    CascadeMux I__4614 (
            .O(N__28313),
            .I(N__28307));
    InMux I__4613 (
            .O(N__28310),
            .I(N__28299));
    InMux I__4612 (
            .O(N__28307),
            .I(N__28299));
    InMux I__4611 (
            .O(N__28306),
            .I(N__28299));
    LocalMux I__4610 (
            .O(N__28299),
            .I(cmd_rdadctmp_11_adj_1439));
    CascadeMux I__4609 (
            .O(N__28296),
            .I(N__28293));
    InMux I__4608 (
            .O(N__28293),
            .I(N__28289));
    CascadeMux I__4607 (
            .O(N__28292),
            .I(N__28286));
    LocalMux I__4606 (
            .O(N__28289),
            .I(N__28283));
    InMux I__4605 (
            .O(N__28286),
            .I(N__28279));
    Span4Mux_h I__4604 (
            .O(N__28283),
            .I(N__28276));
    InMux I__4603 (
            .O(N__28282),
            .I(N__28273));
    LocalMux I__4602 (
            .O(N__28279),
            .I(N__28270));
    Span4Mux_h I__4601 (
            .O(N__28276),
            .I(N__28267));
    LocalMux I__4600 (
            .O(N__28273),
            .I(cmd_rdadctmp_12_adj_1438));
    Odrv12 I__4599 (
            .O(N__28270),
            .I(cmd_rdadctmp_12_adj_1438));
    Odrv4 I__4598 (
            .O(N__28267),
            .I(cmd_rdadctmp_12_adj_1438));
    InMux I__4597 (
            .O(N__28260),
            .I(N__28257));
    LocalMux I__4596 (
            .O(N__28257),
            .I(n22_adj_1640));
    InMux I__4595 (
            .O(N__28254),
            .I(N__28251));
    LocalMux I__4594 (
            .O(N__28251),
            .I(N__28248));
    Sp12to4 I__4593 (
            .O(N__28248),
            .I(N__28245));
    Span12Mux_h I__4592 (
            .O(N__28245),
            .I(N__28242));
    Odrv12 I__4591 (
            .O(N__28242),
            .I(buf_data_iac_2));
    InMux I__4590 (
            .O(N__28239),
            .I(bfn_11_9_0_));
    InMux I__4589 (
            .O(N__28236),
            .I(n19750));
    InMux I__4588 (
            .O(N__28233),
            .I(n19751));
    InMux I__4587 (
            .O(N__28230),
            .I(N__28227));
    LocalMux I__4586 (
            .O(N__28227),
            .I(N__28223));
    CascadeMux I__4585 (
            .O(N__28226),
            .I(N__28220));
    Span4Mux_h I__4584 (
            .O(N__28223),
            .I(N__28217));
    InMux I__4583 (
            .O(N__28220),
            .I(N__28214));
    Odrv4 I__4582 (
            .O(N__28217),
            .I(buf_adcdata_vdc_2));
    LocalMux I__4581 (
            .O(N__28214),
            .I(buf_adcdata_vdc_2));
    CascadeMux I__4580 (
            .O(N__28209),
            .I(n19_adj_1639_cascade_));
    InMux I__4579 (
            .O(N__28206),
            .I(N__28203));
    LocalMux I__4578 (
            .O(N__28203),
            .I(N__28200));
    Span4Mux_h I__4577 (
            .O(N__28200),
            .I(N__28197));
    Odrv4 I__4576 (
            .O(N__28197),
            .I(buf_data_iac_5));
    InMux I__4575 (
            .O(N__28194),
            .I(N__28191));
    LocalMux I__4574 (
            .O(N__28191),
            .I(N__28188));
    Span4Mux_v I__4573 (
            .O(N__28188),
            .I(N__28185));
    Span4Mux_h I__4572 (
            .O(N__28185),
            .I(N__28182));
    Odrv4 I__4571 (
            .O(N__28182),
            .I(n22_adj_1630));
    InMux I__4570 (
            .O(N__28179),
            .I(N__28176));
    LocalMux I__4569 (
            .O(N__28176),
            .I(N__28173));
    Span4Mux_v I__4568 (
            .O(N__28173),
            .I(N__28168));
    InMux I__4567 (
            .O(N__28172),
            .I(N__28163));
    InMux I__4566 (
            .O(N__28171),
            .I(N__28163));
    Sp12to4 I__4565 (
            .O(N__28168),
            .I(N__28160));
    LocalMux I__4564 (
            .O(N__28163),
            .I(buf_adcdata_iac_2));
    Odrv12 I__4563 (
            .O(N__28160),
            .I(buf_adcdata_iac_2));
    InMux I__4562 (
            .O(N__28155),
            .I(N__28148));
    InMux I__4561 (
            .O(N__28154),
            .I(N__28148));
    InMux I__4560 (
            .O(N__28153),
            .I(N__28145));
    LocalMux I__4559 (
            .O(N__28148),
            .I(cmd_rdadctmp_9));
    LocalMux I__4558 (
            .O(N__28145),
            .I(cmd_rdadctmp_9));
    CascadeMux I__4557 (
            .O(N__28140),
            .I(N__28135));
    InMux I__4556 (
            .O(N__28139),
            .I(N__28128));
    InMux I__4555 (
            .O(N__28138),
            .I(N__28128));
    InMux I__4554 (
            .O(N__28135),
            .I(N__28128));
    LocalMux I__4553 (
            .O(N__28128),
            .I(cmd_rdadctmp_10));
    InMux I__4552 (
            .O(N__28125),
            .I(N__28119));
    CascadeMux I__4551 (
            .O(N__28124),
            .I(N__28109));
    CascadeMux I__4550 (
            .O(N__28123),
            .I(N__28105));
    CascadeMux I__4549 (
            .O(N__28122),
            .I(N__28100));
    LocalMux I__4548 (
            .O(N__28119),
            .I(N__28094));
    CascadeMux I__4547 (
            .O(N__28118),
            .I(N__28088));
    InMux I__4546 (
            .O(N__28117),
            .I(N__28083));
    InMux I__4545 (
            .O(N__28116),
            .I(N__28083));
    InMux I__4544 (
            .O(N__28115),
            .I(N__28076));
    InMux I__4543 (
            .O(N__28114),
            .I(N__28076));
    InMux I__4542 (
            .O(N__28113),
            .I(N__28076));
    InMux I__4541 (
            .O(N__28112),
            .I(N__28073));
    InMux I__4540 (
            .O(N__28109),
            .I(N__28070));
    CascadeMux I__4539 (
            .O(N__28108),
            .I(N__28067));
    InMux I__4538 (
            .O(N__28105),
            .I(N__28056));
    InMux I__4537 (
            .O(N__28104),
            .I(N__28056));
    InMux I__4536 (
            .O(N__28103),
            .I(N__28056));
    InMux I__4535 (
            .O(N__28100),
            .I(N__28051));
    InMux I__4534 (
            .O(N__28099),
            .I(N__28051));
    InMux I__4533 (
            .O(N__28098),
            .I(N__28048));
    InMux I__4532 (
            .O(N__28097),
            .I(N__28042));
    Span4Mux_h I__4531 (
            .O(N__28094),
            .I(N__28039));
    InMux I__4530 (
            .O(N__28093),
            .I(N__28036));
    InMux I__4529 (
            .O(N__28092),
            .I(N__28031));
    InMux I__4528 (
            .O(N__28091),
            .I(N__28028));
    InMux I__4527 (
            .O(N__28088),
            .I(N__28025));
    LocalMux I__4526 (
            .O(N__28083),
            .I(N__28020));
    LocalMux I__4525 (
            .O(N__28076),
            .I(N__28020));
    LocalMux I__4524 (
            .O(N__28073),
            .I(N__28017));
    LocalMux I__4523 (
            .O(N__28070),
            .I(N__28014));
    InMux I__4522 (
            .O(N__28067),
            .I(N__28009));
    InMux I__4521 (
            .O(N__28066),
            .I(N__28009));
    CascadeMux I__4520 (
            .O(N__28065),
            .I(N__28006));
    InMux I__4519 (
            .O(N__28064),
            .I(N__28002));
    InMux I__4518 (
            .O(N__28063),
            .I(N__27999));
    LocalMux I__4517 (
            .O(N__28056),
            .I(N__27996));
    LocalMux I__4516 (
            .O(N__28051),
            .I(N__27991));
    LocalMux I__4515 (
            .O(N__28048),
            .I(N__27991));
    InMux I__4514 (
            .O(N__28047),
            .I(N__27984));
    InMux I__4513 (
            .O(N__28046),
            .I(N__27984));
    InMux I__4512 (
            .O(N__28045),
            .I(N__27984));
    LocalMux I__4511 (
            .O(N__28042),
            .I(N__27979));
    Span4Mux_v I__4510 (
            .O(N__28039),
            .I(N__27979));
    LocalMux I__4509 (
            .O(N__28036),
            .I(N__27976));
    InMux I__4508 (
            .O(N__28035),
            .I(N__27970));
    InMux I__4507 (
            .O(N__28034),
            .I(N__27970));
    LocalMux I__4506 (
            .O(N__28031),
            .I(N__27959));
    LocalMux I__4505 (
            .O(N__28028),
            .I(N__27959));
    LocalMux I__4504 (
            .O(N__28025),
            .I(N__27959));
    Span4Mux_v I__4503 (
            .O(N__28020),
            .I(N__27959));
    Span4Mux_v I__4502 (
            .O(N__28017),
            .I(N__27959));
    Sp12to4 I__4501 (
            .O(N__28014),
            .I(N__27954));
    LocalMux I__4500 (
            .O(N__28009),
            .I(N__27954));
    InMux I__4499 (
            .O(N__28006),
            .I(N__27949));
    InMux I__4498 (
            .O(N__28005),
            .I(N__27949));
    LocalMux I__4497 (
            .O(N__28002),
            .I(N__27946));
    LocalMux I__4496 (
            .O(N__27999),
            .I(N__27943));
    Span4Mux_v I__4495 (
            .O(N__27996),
            .I(N__27938));
    Span4Mux_h I__4494 (
            .O(N__27991),
            .I(N__27938));
    LocalMux I__4493 (
            .O(N__27984),
            .I(N__27931));
    Span4Mux_h I__4492 (
            .O(N__27979),
            .I(N__27931));
    Span4Mux_h I__4491 (
            .O(N__27976),
            .I(N__27931));
    InMux I__4490 (
            .O(N__27975),
            .I(N__27928));
    LocalMux I__4489 (
            .O(N__27970),
            .I(N__27923));
    Span4Mux_v I__4488 (
            .O(N__27959),
            .I(N__27923));
    Span12Mux_v I__4487 (
            .O(N__27954),
            .I(N__27920));
    LocalMux I__4486 (
            .O(N__27949),
            .I(N__27911));
    Span4Mux_h I__4485 (
            .O(N__27946),
            .I(N__27911));
    Span4Mux_v I__4484 (
            .O(N__27943),
            .I(N__27911));
    Span4Mux_v I__4483 (
            .O(N__27938),
            .I(N__27911));
    Span4Mux_v I__4482 (
            .O(N__27931),
            .I(N__27908));
    LocalMux I__4481 (
            .O(N__27928),
            .I(n12498));
    Odrv4 I__4480 (
            .O(N__27923),
            .I(n12498));
    Odrv12 I__4479 (
            .O(N__27920),
            .I(n12498));
    Odrv4 I__4478 (
            .O(N__27911),
            .I(n12498));
    Odrv4 I__4477 (
            .O(N__27908),
            .I(n12498));
    InMux I__4476 (
            .O(N__27897),
            .I(N__27894));
    LocalMux I__4475 (
            .O(N__27894),
            .I(N__27891));
    Span4Mux_h I__4474 (
            .O(N__27891),
            .I(N__27888));
    Span4Mux_h I__4473 (
            .O(N__27888),
            .I(N__27883));
    InMux I__4472 (
            .O(N__27887),
            .I(N__27878));
    InMux I__4471 (
            .O(N__27886),
            .I(N__27878));
    Span4Mux_h I__4470 (
            .O(N__27883),
            .I(N__27875));
    LocalMux I__4469 (
            .O(N__27878),
            .I(buf_adcdata_vac_2));
    Odrv4 I__4468 (
            .O(N__27875),
            .I(buf_adcdata_vac_2));
    InMux I__4467 (
            .O(N__27870),
            .I(N__27867));
    LocalMux I__4466 (
            .O(N__27867),
            .I(N__27863));
    CascadeMux I__4465 (
            .O(N__27866),
            .I(N__27860));
    Span4Mux_v I__4464 (
            .O(N__27863),
            .I(N__27857));
    InMux I__4463 (
            .O(N__27860),
            .I(N__27854));
    Odrv4 I__4462 (
            .O(N__27857),
            .I(buf_adcdata_vdc_3));
    LocalMux I__4461 (
            .O(N__27854),
            .I(buf_adcdata_vdc_3));
    InMux I__4460 (
            .O(N__27849),
            .I(N__27846));
    LocalMux I__4459 (
            .O(N__27846),
            .I(\ADC_VDC.n21952 ));
    InMux I__4458 (
            .O(N__27843),
            .I(bfn_11_5_0_));
    InMux I__4457 (
            .O(N__27840),
            .I(n19746));
    InMux I__4456 (
            .O(N__27837),
            .I(n19747));
    InMux I__4455 (
            .O(N__27834),
            .I(n19748));
    InMux I__4454 (
            .O(N__27831),
            .I(n19749));
    CascadeMux I__4453 (
            .O(N__27828),
            .I(N__27825));
    InMux I__4452 (
            .O(N__27825),
            .I(N__27817));
    InMux I__4451 (
            .O(N__27824),
            .I(N__27817));
    InMux I__4450 (
            .O(N__27823),
            .I(N__27814));
    InMux I__4449 (
            .O(N__27822),
            .I(N__27811));
    LocalMux I__4448 (
            .O(N__27817),
            .I(N__27803));
    LocalMux I__4447 (
            .O(N__27814),
            .I(N__27803));
    LocalMux I__4446 (
            .O(N__27811),
            .I(N__27803));
    InMux I__4445 (
            .O(N__27810),
            .I(N__27800));
    Span4Mux_v I__4444 (
            .O(N__27803),
            .I(N__27795));
    LocalMux I__4443 (
            .O(N__27800),
            .I(N__27795));
    Span4Mux_v I__4442 (
            .O(N__27795),
            .I(N__27792));
    Span4Mux_v I__4441 (
            .O(N__27792),
            .I(N__27789));
    Sp12to4 I__4440 (
            .O(N__27789),
            .I(N__27786));
    Span12Mux_h I__4439 (
            .O(N__27786),
            .I(N__27783));
    Odrv12 I__4438 (
            .O(N__27783),
            .I(ICE_SPI_SCLK));
    InMux I__4437 (
            .O(N__27780),
            .I(N__27777));
    LocalMux I__4436 (
            .O(N__27777),
            .I(\comm_spi.n14596 ));
    SRMux I__4435 (
            .O(N__27774),
            .I(N__27771));
    LocalMux I__4434 (
            .O(N__27771),
            .I(N__27768));
    Odrv4 I__4433 (
            .O(N__27768),
            .I(\comm_spi.iclk_N_762 ));
    InMux I__4432 (
            .O(N__27765),
            .I(N__27762));
    LocalMux I__4431 (
            .O(N__27762),
            .I(n22255));
    SRMux I__4430 (
            .O(N__27759),
            .I(N__27753));
    SRMux I__4429 (
            .O(N__27758),
            .I(N__27750));
    SRMux I__4428 (
            .O(N__27757),
            .I(N__27745));
    SRMux I__4427 (
            .O(N__27756),
            .I(N__27742));
    LocalMux I__4426 (
            .O(N__27753),
            .I(N__27737));
    LocalMux I__4425 (
            .O(N__27750),
            .I(N__27737));
    SRMux I__4424 (
            .O(N__27749),
            .I(N__27734));
    SRMux I__4423 (
            .O(N__27748),
            .I(N__27731));
    LocalMux I__4422 (
            .O(N__27745),
            .I(N__27726));
    LocalMux I__4421 (
            .O(N__27742),
            .I(N__27723));
    Span4Mux_v I__4420 (
            .O(N__27737),
            .I(N__27716));
    LocalMux I__4419 (
            .O(N__27734),
            .I(N__27716));
    LocalMux I__4418 (
            .O(N__27731),
            .I(N__27716));
    SRMux I__4417 (
            .O(N__27730),
            .I(N__27713));
    SRMux I__4416 (
            .O(N__27729),
            .I(N__27710));
    Span4Mux_v I__4415 (
            .O(N__27726),
            .I(N__27703));
    Span4Mux_h I__4414 (
            .O(N__27723),
            .I(N__27700));
    Span4Mux_v I__4413 (
            .O(N__27716),
            .I(N__27693));
    LocalMux I__4412 (
            .O(N__27713),
            .I(N__27693));
    LocalMux I__4411 (
            .O(N__27710),
            .I(N__27693));
    SRMux I__4410 (
            .O(N__27709),
            .I(N__27690));
    SRMux I__4409 (
            .O(N__27708),
            .I(N__27687));
    SRMux I__4408 (
            .O(N__27707),
            .I(N__27684));
    SRMux I__4407 (
            .O(N__27706),
            .I(N__27681));
    Span4Mux_v I__4406 (
            .O(N__27703),
            .I(N__27678));
    Span4Mux_v I__4405 (
            .O(N__27700),
            .I(N__27675));
    Span4Mux_v I__4404 (
            .O(N__27693),
            .I(N__27668));
    LocalMux I__4403 (
            .O(N__27690),
            .I(N__27668));
    LocalMux I__4402 (
            .O(N__27687),
            .I(N__27668));
    LocalMux I__4401 (
            .O(N__27684),
            .I(N__27663));
    LocalMux I__4400 (
            .O(N__27681),
            .I(N__27663));
    Span4Mux_v I__4399 (
            .O(N__27678),
            .I(N__27660));
    Span4Mux_v I__4398 (
            .O(N__27675),
            .I(N__27657));
    Span4Mux_v I__4397 (
            .O(N__27668),
            .I(N__27652));
    Span4Mux_v I__4396 (
            .O(N__27663),
            .I(N__27652));
    Span4Mux_h I__4395 (
            .O(N__27660),
            .I(N__27649));
    Span4Mux_h I__4394 (
            .O(N__27657),
            .I(N__27646));
    Sp12to4 I__4393 (
            .O(N__27652),
            .I(N__27643));
    Odrv4 I__4392 (
            .O(N__27649),
            .I(iac_raw_buf_N_734));
    Odrv4 I__4391 (
            .O(N__27646),
            .I(iac_raw_buf_N_734));
    Odrv12 I__4390 (
            .O(N__27643),
            .I(iac_raw_buf_N_734));
    IoInMux I__4389 (
            .O(N__27636),
            .I(N__27633));
    LocalMux I__4388 (
            .O(N__27633),
            .I(N__27630));
    Span4Mux_s1_v I__4387 (
            .O(N__27630),
            .I(N__27626));
    InMux I__4386 (
            .O(N__27629),
            .I(N__27622));
    Sp12to4 I__4385 (
            .O(N__27626),
            .I(N__27619));
    CascadeMux I__4384 (
            .O(N__27625),
            .I(N__27616));
    LocalMux I__4383 (
            .O(N__27622),
            .I(N__27613));
    Span12Mux_h I__4382 (
            .O(N__27619),
            .I(N__27610));
    InMux I__4381 (
            .O(N__27616),
            .I(N__27607));
    Span4Mux_h I__4380 (
            .O(N__27613),
            .I(N__27604));
    Odrv12 I__4379 (
            .O(N__27610),
            .I(IAC_OSR0));
    LocalMux I__4378 (
            .O(N__27607),
            .I(IAC_OSR0));
    Odrv4 I__4377 (
            .O(N__27604),
            .I(IAC_OSR0));
    CascadeMux I__4376 (
            .O(N__27597),
            .I(n12367_cascade_));
    CascadeMux I__4375 (
            .O(N__27594),
            .I(n16563_cascade_));
    CascadeMux I__4374 (
            .O(N__27591),
            .I(N__27587));
    CascadeMux I__4373 (
            .O(N__27590),
            .I(N__27583));
    InMux I__4372 (
            .O(N__27587),
            .I(N__27580));
    InMux I__4371 (
            .O(N__27586),
            .I(N__27577));
    InMux I__4370 (
            .O(N__27583),
            .I(N__27574));
    LocalMux I__4369 (
            .O(N__27580),
            .I(N__27571));
    LocalMux I__4368 (
            .O(N__27577),
            .I(N__27568));
    LocalMux I__4367 (
            .O(N__27574),
            .I(N__27565));
    Odrv4 I__4366 (
            .O(N__27571),
            .I(cmd_rdadctmp_27));
    Odrv4 I__4365 (
            .O(N__27568),
            .I(cmd_rdadctmp_27));
    Odrv4 I__4364 (
            .O(N__27565),
            .I(cmd_rdadctmp_27));
    CascadeMux I__4363 (
            .O(N__27558),
            .I(N__27555));
    InMux I__4362 (
            .O(N__27555),
            .I(N__27552));
    LocalMux I__4361 (
            .O(N__27552),
            .I(N__27547));
    InMux I__4360 (
            .O(N__27551),
            .I(N__27544));
    InMux I__4359 (
            .O(N__27550),
            .I(N__27541));
    Odrv4 I__4358 (
            .O(N__27547),
            .I(cmd_rdadctmp_28));
    LocalMux I__4357 (
            .O(N__27544),
            .I(cmd_rdadctmp_28));
    LocalMux I__4356 (
            .O(N__27541),
            .I(cmd_rdadctmp_28));
    InMux I__4355 (
            .O(N__27534),
            .I(N__27531));
    LocalMux I__4354 (
            .O(N__27531),
            .I(N__27528));
    Span4Mux_v I__4353 (
            .O(N__27528),
            .I(N__27525));
    Span4Mux_h I__4352 (
            .O(N__27525),
            .I(N__27522));
    Odrv4 I__4351 (
            .O(N__27522),
            .I(n19_adj_1527));
    CascadeMux I__4350 (
            .O(N__27519),
            .I(n22279_cascade_));
    InMux I__4349 (
            .O(N__27516),
            .I(N__27513));
    LocalMux I__4348 (
            .O(N__27513),
            .I(n17_adj_1526));
    InMux I__4347 (
            .O(N__27510),
            .I(N__27507));
    LocalMux I__4346 (
            .O(N__27507),
            .I(N__27504));
    Odrv12 I__4345 (
            .O(N__27504),
            .I(n23_adj_1529));
    CascadeMux I__4344 (
            .O(N__27501),
            .I(n22363_cascade_));
    InMux I__4343 (
            .O(N__27498),
            .I(N__27495));
    LocalMux I__4342 (
            .O(N__27495),
            .I(N__27492));
    Odrv4 I__4341 (
            .O(N__27492),
            .I(n21285));
    InMux I__4340 (
            .O(N__27489),
            .I(N__27486));
    LocalMux I__4339 (
            .O(N__27486),
            .I(n22282));
    CascadeMux I__4338 (
            .O(N__27483),
            .I(n22366_cascade_));
    InMux I__4337 (
            .O(N__27480),
            .I(N__27476));
    InMux I__4336 (
            .O(N__27479),
            .I(N__27472));
    LocalMux I__4335 (
            .O(N__27476),
            .I(N__27469));
    InMux I__4334 (
            .O(N__27475),
            .I(N__27466));
    LocalMux I__4333 (
            .O(N__27472),
            .I(buf_dds1_15));
    Odrv4 I__4332 (
            .O(N__27469),
            .I(buf_dds1_15));
    LocalMux I__4331 (
            .O(N__27466),
            .I(buf_dds1_15));
    InMux I__4330 (
            .O(N__27459),
            .I(N__27456));
    LocalMux I__4329 (
            .O(N__27456),
            .I(n16_adj_1525));
    InMux I__4328 (
            .O(N__27453),
            .I(N__27450));
    LocalMux I__4327 (
            .O(N__27450),
            .I(N__27445));
    InMux I__4326 (
            .O(N__27449),
            .I(N__27442));
    CascadeMux I__4325 (
            .O(N__27448),
            .I(N__27435));
    Span4Mux_v I__4324 (
            .O(N__27445),
            .I(N__27425));
    LocalMux I__4323 (
            .O(N__27442),
            .I(N__27425));
    InMux I__4322 (
            .O(N__27441),
            .I(N__27422));
    InMux I__4321 (
            .O(N__27440),
            .I(N__27419));
    InMux I__4320 (
            .O(N__27439),
            .I(N__27416));
    InMux I__4319 (
            .O(N__27438),
            .I(N__27413));
    InMux I__4318 (
            .O(N__27435),
            .I(N__27410));
    InMux I__4317 (
            .O(N__27434),
            .I(N__27405));
    InMux I__4316 (
            .O(N__27433),
            .I(N__27405));
    InMux I__4315 (
            .O(N__27432),
            .I(N__27398));
    InMux I__4314 (
            .O(N__27431),
            .I(N__27398));
    InMux I__4313 (
            .O(N__27430),
            .I(N__27398));
    Span4Mux_h I__4312 (
            .O(N__27425),
            .I(N__27395));
    LocalMux I__4311 (
            .O(N__27422),
            .I(N__27392));
    LocalMux I__4310 (
            .O(N__27419),
            .I(adc_state_1_adj_1417));
    LocalMux I__4309 (
            .O(N__27416),
            .I(adc_state_1_adj_1417));
    LocalMux I__4308 (
            .O(N__27413),
            .I(adc_state_1_adj_1417));
    LocalMux I__4307 (
            .O(N__27410),
            .I(adc_state_1_adj_1417));
    LocalMux I__4306 (
            .O(N__27405),
            .I(adc_state_1_adj_1417));
    LocalMux I__4305 (
            .O(N__27398),
            .I(adc_state_1_adj_1417));
    Odrv4 I__4304 (
            .O(N__27395),
            .I(adc_state_1_adj_1417));
    Odrv12 I__4303 (
            .O(N__27392),
            .I(adc_state_1_adj_1417));
    CascadeMux I__4302 (
            .O(N__27375),
            .I(N__27370));
    CascadeMux I__4301 (
            .O(N__27374),
            .I(N__27367));
    InMux I__4300 (
            .O(N__27373),
            .I(N__27364));
    InMux I__4299 (
            .O(N__27370),
            .I(N__27361));
    InMux I__4298 (
            .O(N__27367),
            .I(N__27358));
    LocalMux I__4297 (
            .O(N__27364),
            .I(N__27355));
    LocalMux I__4296 (
            .O(N__27361),
            .I(cmd_rdadctmp_24));
    LocalMux I__4295 (
            .O(N__27358),
            .I(cmd_rdadctmp_24));
    Odrv4 I__4294 (
            .O(N__27355),
            .I(cmd_rdadctmp_24));
    InMux I__4293 (
            .O(N__27348),
            .I(N__27345));
    LocalMux I__4292 (
            .O(N__27345),
            .I(N__27340));
    InMux I__4291 (
            .O(N__27344),
            .I(N__27337));
    InMux I__4290 (
            .O(N__27343),
            .I(N__27334));
    Span12Mux_v I__4289 (
            .O(N__27340),
            .I(N__27331));
    LocalMux I__4288 (
            .O(N__27337),
            .I(N__27328));
    LocalMux I__4287 (
            .O(N__27334),
            .I(buf_adcdata_iac_16));
    Odrv12 I__4286 (
            .O(N__27331),
            .I(buf_adcdata_iac_16));
    Odrv4 I__4285 (
            .O(N__27328),
            .I(buf_adcdata_iac_16));
    InMux I__4284 (
            .O(N__27321),
            .I(N__27317));
    CascadeMux I__4283 (
            .O(N__27320),
            .I(N__27314));
    LocalMux I__4282 (
            .O(N__27317),
            .I(N__27310));
    InMux I__4281 (
            .O(N__27314),
            .I(N__27305));
    InMux I__4280 (
            .O(N__27313),
            .I(N__27305));
    Odrv12 I__4279 (
            .O(N__27310),
            .I(cmd_rdadctmp_26));
    LocalMux I__4278 (
            .O(N__27305),
            .I(cmd_rdadctmp_26));
    InMux I__4277 (
            .O(N__27300),
            .I(N__27291));
    InMux I__4276 (
            .O(N__27299),
            .I(N__27284));
    InMux I__4275 (
            .O(N__27298),
            .I(N__27284));
    InMux I__4274 (
            .O(N__27297),
            .I(N__27284));
    InMux I__4273 (
            .O(N__27296),
            .I(N__27281));
    InMux I__4272 (
            .O(N__27295),
            .I(N__27276));
    InMux I__4271 (
            .O(N__27294),
            .I(N__27276));
    LocalMux I__4270 (
            .O(N__27291),
            .I(N__27273));
    LocalMux I__4269 (
            .O(N__27284),
            .I(N__27268));
    LocalMux I__4268 (
            .O(N__27281),
            .I(N__27268));
    LocalMux I__4267 (
            .O(N__27276),
            .I(N__27265));
    Span4Mux_h I__4266 (
            .O(N__27273),
            .I(N__27259));
    Span4Mux_v I__4265 (
            .O(N__27268),
            .I(N__27259));
    Span4Mux_h I__4264 (
            .O(N__27265),
            .I(N__27256));
    InMux I__4263 (
            .O(N__27264),
            .I(N__27253));
    Odrv4 I__4262 (
            .O(N__27259),
            .I(n12395));
    Odrv4 I__4261 (
            .O(N__27256),
            .I(n12395));
    LocalMux I__4260 (
            .O(N__27253),
            .I(n12395));
    CascadeMux I__4259 (
            .O(N__27246),
            .I(N__27243));
    InMux I__4258 (
            .O(N__27243),
            .I(N__27240));
    LocalMux I__4257 (
            .O(N__27240),
            .I(\CLK_DDS.tmp_buf_11 ));
    CascadeMux I__4256 (
            .O(N__27237),
            .I(N__27234));
    InMux I__4255 (
            .O(N__27234),
            .I(N__27231));
    LocalMux I__4254 (
            .O(N__27231),
            .I(\CLK_DDS.tmp_buf_12 ));
    CascadeMux I__4253 (
            .O(N__27228),
            .I(N__27224));
    CascadeMux I__4252 (
            .O(N__27227),
            .I(N__27221));
    InMux I__4251 (
            .O(N__27224),
            .I(N__27218));
    InMux I__4250 (
            .O(N__27221),
            .I(N__27215));
    LocalMux I__4249 (
            .O(N__27218),
            .I(tmp_buf_15_adj_1455));
    LocalMux I__4248 (
            .O(N__27215),
            .I(tmp_buf_15_adj_1455));
    CascadeMux I__4247 (
            .O(N__27210),
            .I(N__27207));
    InMux I__4246 (
            .O(N__27207),
            .I(N__27204));
    LocalMux I__4245 (
            .O(N__27204),
            .I(\CLK_DDS.tmp_buf_7 ));
    InMux I__4244 (
            .O(N__27201),
            .I(N__27196));
    InMux I__4243 (
            .O(N__27200),
            .I(N__27193));
    InMux I__4242 (
            .O(N__27199),
            .I(N__27190));
    LocalMux I__4241 (
            .O(N__27196),
            .I(N__27187));
    LocalMux I__4240 (
            .O(N__27193),
            .I(buf_dds1_8));
    LocalMux I__4239 (
            .O(N__27190),
            .I(buf_dds1_8));
    Odrv4 I__4238 (
            .O(N__27187),
            .I(buf_dds1_8));
    InMux I__4237 (
            .O(N__27180),
            .I(N__27177));
    LocalMux I__4236 (
            .O(N__27177),
            .I(N__27172));
    InMux I__4235 (
            .O(N__27176),
            .I(N__27169));
    InMux I__4234 (
            .O(N__27175),
            .I(N__27166));
    Span4Mux_h I__4233 (
            .O(N__27172),
            .I(N__27163));
    LocalMux I__4232 (
            .O(N__27169),
            .I(buf_dds1_13));
    LocalMux I__4231 (
            .O(N__27166),
            .I(buf_dds1_13));
    Odrv4 I__4230 (
            .O(N__27163),
            .I(buf_dds1_13));
    CascadeMux I__4229 (
            .O(N__27156),
            .I(n11347_cascade_));
    CEMux I__4228 (
            .O(N__27153),
            .I(N__27150));
    LocalMux I__4227 (
            .O(N__27150),
            .I(n11919));
    InMux I__4226 (
            .O(N__27147),
            .I(N__27144));
    LocalMux I__4225 (
            .O(N__27144),
            .I(buf_control_7));
    CascadeMux I__4224 (
            .O(N__27141),
            .I(N__27138));
    InMux I__4223 (
            .O(N__27138),
            .I(N__27135));
    LocalMux I__4222 (
            .O(N__27135),
            .I(\CLK_DDS.tmp_buf_10 ));
    IoInMux I__4221 (
            .O(N__27132),
            .I(N__27129));
    LocalMux I__4220 (
            .O(N__27129),
            .I(N__27126));
    IoSpan4Mux I__4219 (
            .O(N__27126),
            .I(N__27123));
    IoSpan4Mux I__4218 (
            .O(N__27123),
            .I(N__27120));
    Sp12to4 I__4217 (
            .O(N__27120),
            .I(N__27116));
    CascadeMux I__4216 (
            .O(N__27119),
            .I(N__27113));
    Span12Mux_s7_v I__4215 (
            .O(N__27116),
            .I(N__27110));
    InMux I__4214 (
            .O(N__27113),
            .I(N__27107));
    Odrv12 I__4213 (
            .O(N__27110),
            .I(DDS_SCK1));
    LocalMux I__4212 (
            .O(N__27107),
            .I(DDS_SCK1));
    InMux I__4211 (
            .O(N__27102),
            .I(N__27098));
    CascadeMux I__4210 (
            .O(N__27101),
            .I(N__27095));
    LocalMux I__4209 (
            .O(N__27098),
            .I(N__27092));
    InMux I__4208 (
            .O(N__27095),
            .I(N__27089));
    Odrv4 I__4207 (
            .O(N__27092),
            .I(buf_adcdata_vdc_18));
    LocalMux I__4206 (
            .O(N__27089),
            .I(buf_adcdata_vdc_18));
    InMux I__4205 (
            .O(N__27084),
            .I(N__27081));
    LocalMux I__4204 (
            .O(N__27081),
            .I(N__27077));
    InMux I__4203 (
            .O(N__27080),
            .I(N__27073));
    Span12Mux_h I__4202 (
            .O(N__27077),
            .I(N__27070));
    InMux I__4201 (
            .O(N__27076),
            .I(N__27067));
    LocalMux I__4200 (
            .O(N__27073),
            .I(buf_adcdata_vac_18));
    Odrv12 I__4199 (
            .O(N__27070),
            .I(buf_adcdata_vac_18));
    LocalMux I__4198 (
            .O(N__27067),
            .I(buf_adcdata_vac_18));
    InMux I__4197 (
            .O(N__27060),
            .I(N__27057));
    LocalMux I__4196 (
            .O(N__27057),
            .I(N__27054));
    Span4Mux_h I__4195 (
            .O(N__27054),
            .I(N__27051));
    Span4Mux_v I__4194 (
            .O(N__27051),
            .I(N__27048));
    Odrv4 I__4193 (
            .O(N__27048),
            .I(n21081));
    InMux I__4192 (
            .O(N__27045),
            .I(N__27041));
    InMux I__4191 (
            .O(N__27044),
            .I(N__27038));
    LocalMux I__4190 (
            .O(N__27041),
            .I(cmd_rdadctmp_6));
    LocalMux I__4189 (
            .O(N__27038),
            .I(cmd_rdadctmp_6));
    InMux I__4188 (
            .O(N__27033),
            .I(N__27030));
    LocalMux I__4187 (
            .O(N__27030),
            .I(N__27027));
    Span4Mux_v I__4186 (
            .O(N__27027),
            .I(N__27023));
    InMux I__4185 (
            .O(N__27026),
            .I(N__27020));
    Odrv4 I__4184 (
            .O(N__27023),
            .I(cmd_rdadctmp_4));
    LocalMux I__4183 (
            .O(N__27020),
            .I(cmd_rdadctmp_4));
    InMux I__4182 (
            .O(N__27015),
            .I(N__27009));
    InMux I__4181 (
            .O(N__27014),
            .I(N__27009));
    LocalMux I__4180 (
            .O(N__27009),
            .I(cmd_rdadctmp_5));
    InMux I__4179 (
            .O(N__27006),
            .I(N__27003));
    LocalMux I__4178 (
            .O(N__27003),
            .I(N__27000));
    Span12Mux_h I__4177 (
            .O(N__27000),
            .I(N__26997));
    Span12Mux_v I__4176 (
            .O(N__26997),
            .I(N__26994));
    Odrv12 I__4175 (
            .O(N__26994),
            .I(THERMOSTAT));
    InMux I__4174 (
            .O(N__26991),
            .I(N__26988));
    LocalMux I__4173 (
            .O(N__26988),
            .I(N__26985));
    Span4Mux_h I__4172 (
            .O(N__26985),
            .I(N__26982));
    Span4Mux_h I__4171 (
            .O(N__26982),
            .I(N__26979));
    Span4Mux_h I__4170 (
            .O(N__26979),
            .I(N__26976));
    Odrv4 I__4169 (
            .O(N__26976),
            .I(buf_data_iac_0));
    InMux I__4168 (
            .O(N__26973),
            .I(N__26970));
    LocalMux I__4167 (
            .O(N__26970),
            .I(N__26967));
    Span4Mux_h I__4166 (
            .O(N__26967),
            .I(N__26963));
    CascadeMux I__4165 (
            .O(N__26966),
            .I(N__26960));
    Span4Mux_h I__4164 (
            .O(N__26963),
            .I(N__26956));
    InMux I__4163 (
            .O(N__26960),
            .I(N__26953));
    InMux I__4162 (
            .O(N__26959),
            .I(N__26950));
    Span4Mux_h I__4161 (
            .O(N__26956),
            .I(N__26947));
    LocalMux I__4160 (
            .O(N__26953),
            .I(buf_adcdata_iac_0));
    LocalMux I__4159 (
            .O(N__26950),
            .I(buf_adcdata_iac_0));
    Odrv4 I__4158 (
            .O(N__26947),
            .I(buf_adcdata_iac_0));
    CascadeMux I__4157 (
            .O(N__26940),
            .I(N__26937));
    InMux I__4156 (
            .O(N__26937),
            .I(N__26934));
    LocalMux I__4155 (
            .O(N__26934),
            .I(N__26931));
    Span4Mux_h I__4154 (
            .O(N__26931),
            .I(N__26927));
    CascadeMux I__4153 (
            .O(N__26930),
            .I(N__26924));
    Span4Mux_v I__4152 (
            .O(N__26927),
            .I(N__26920));
    InMux I__4151 (
            .O(N__26924),
            .I(N__26917));
    InMux I__4150 (
            .O(N__26923),
            .I(N__26914));
    Odrv4 I__4149 (
            .O(N__26920),
            .I(cmd_rdadctmp_8_adj_1442));
    LocalMux I__4148 (
            .O(N__26917),
            .I(cmd_rdadctmp_8_adj_1442));
    LocalMux I__4147 (
            .O(N__26914),
            .I(cmd_rdadctmp_8_adj_1442));
    InMux I__4146 (
            .O(N__26907),
            .I(N__26904));
    LocalMux I__4145 (
            .O(N__26904),
            .I(N__26901));
    Span4Mux_v I__4144 (
            .O(N__26901),
            .I(N__26898));
    Span4Mux_h I__4143 (
            .O(N__26898),
            .I(N__26895));
    Span4Mux_h I__4142 (
            .O(N__26895),
            .I(N__26890));
    InMux I__4141 (
            .O(N__26894),
            .I(N__26885));
    InMux I__4140 (
            .O(N__26893),
            .I(N__26885));
    Odrv4 I__4139 (
            .O(N__26890),
            .I(buf_adcdata_vac_0));
    LocalMux I__4138 (
            .O(N__26885),
            .I(buf_adcdata_vac_0));
    CascadeMux I__4137 (
            .O(N__26880),
            .I(N__26876));
    InMux I__4136 (
            .O(N__26879),
            .I(N__26871));
    InMux I__4135 (
            .O(N__26876),
            .I(N__26871));
    LocalMux I__4134 (
            .O(N__26871),
            .I(N__26868));
    Span4Mux_h I__4133 (
            .O(N__26868),
            .I(N__26864));
    InMux I__4132 (
            .O(N__26867),
            .I(N__26861));
    Odrv4 I__4131 (
            .O(N__26864),
            .I(cmd_rdadctmp_8));
    LocalMux I__4130 (
            .O(N__26861),
            .I(cmd_rdadctmp_8));
    InMux I__4129 (
            .O(N__26856),
            .I(N__26853));
    LocalMux I__4128 (
            .O(N__26853),
            .I(N__26826));
    InMux I__4127 (
            .O(N__26852),
            .I(N__26821));
    InMux I__4126 (
            .O(N__26851),
            .I(N__26821));
    InMux I__4125 (
            .O(N__26850),
            .I(N__26816));
    InMux I__4124 (
            .O(N__26849),
            .I(N__26798));
    InMux I__4123 (
            .O(N__26848),
            .I(N__26798));
    InMux I__4122 (
            .O(N__26847),
            .I(N__26798));
    InMux I__4121 (
            .O(N__26846),
            .I(N__26798));
    InMux I__4120 (
            .O(N__26845),
            .I(N__26798));
    InMux I__4119 (
            .O(N__26844),
            .I(N__26798));
    InMux I__4118 (
            .O(N__26843),
            .I(N__26798));
    InMux I__4117 (
            .O(N__26842),
            .I(N__26798));
    InMux I__4116 (
            .O(N__26841),
            .I(N__26789));
    InMux I__4115 (
            .O(N__26840),
            .I(N__26789));
    InMux I__4114 (
            .O(N__26839),
            .I(N__26789));
    InMux I__4113 (
            .O(N__26838),
            .I(N__26789));
    CascadeMux I__4112 (
            .O(N__26837),
            .I(N__26786));
    InMux I__4111 (
            .O(N__26836),
            .I(N__26779));
    InMux I__4110 (
            .O(N__26835),
            .I(N__26773));
    InMux I__4109 (
            .O(N__26834),
            .I(N__26773));
    InMux I__4108 (
            .O(N__26833),
            .I(N__26768));
    InMux I__4107 (
            .O(N__26832),
            .I(N__26768));
    InMux I__4106 (
            .O(N__26831),
            .I(N__26757));
    InMux I__4105 (
            .O(N__26830),
            .I(N__26754));
    InMux I__4104 (
            .O(N__26829),
            .I(N__26751));
    Span4Mux_v I__4103 (
            .O(N__26826),
            .I(N__26744));
    LocalMux I__4102 (
            .O(N__26821),
            .I(N__26744));
    InMux I__4101 (
            .O(N__26820),
            .I(N__26739));
    InMux I__4100 (
            .O(N__26819),
            .I(N__26739));
    LocalMux I__4099 (
            .O(N__26816),
            .I(N__26736));
    InMux I__4098 (
            .O(N__26815),
            .I(N__26732));
    LocalMux I__4097 (
            .O(N__26798),
            .I(N__26727));
    LocalMux I__4096 (
            .O(N__26789),
            .I(N__26727));
    InMux I__4095 (
            .O(N__26786),
            .I(N__26717));
    InMux I__4094 (
            .O(N__26785),
            .I(N__26717));
    InMux I__4093 (
            .O(N__26784),
            .I(N__26717));
    InMux I__4092 (
            .O(N__26783),
            .I(N__26714));
    InMux I__4091 (
            .O(N__26782),
            .I(N__26711));
    LocalMux I__4090 (
            .O(N__26779),
            .I(N__26708));
    InMux I__4089 (
            .O(N__26778),
            .I(N__26705));
    LocalMux I__4088 (
            .O(N__26773),
            .I(N__26700));
    LocalMux I__4087 (
            .O(N__26768),
            .I(N__26700));
    InMux I__4086 (
            .O(N__26767),
            .I(N__26693));
    InMux I__4085 (
            .O(N__26766),
            .I(N__26693));
    InMux I__4084 (
            .O(N__26765),
            .I(N__26693));
    InMux I__4083 (
            .O(N__26764),
            .I(N__26686));
    InMux I__4082 (
            .O(N__26763),
            .I(N__26686));
    InMux I__4081 (
            .O(N__26762),
            .I(N__26686));
    InMux I__4080 (
            .O(N__26761),
            .I(N__26681));
    InMux I__4079 (
            .O(N__26760),
            .I(N__26681));
    LocalMux I__4078 (
            .O(N__26757),
            .I(N__26674));
    LocalMux I__4077 (
            .O(N__26754),
            .I(N__26674));
    LocalMux I__4076 (
            .O(N__26751),
            .I(N__26674));
    InMux I__4075 (
            .O(N__26750),
            .I(N__26669));
    InMux I__4074 (
            .O(N__26749),
            .I(N__26669));
    Span4Mux_v I__4073 (
            .O(N__26744),
            .I(N__26662));
    LocalMux I__4072 (
            .O(N__26739),
            .I(N__26662));
    Span4Mux_h I__4071 (
            .O(N__26736),
            .I(N__26662));
    InMux I__4070 (
            .O(N__26735),
            .I(N__26659));
    LocalMux I__4069 (
            .O(N__26732),
            .I(N__26656));
    Span4Mux_v I__4068 (
            .O(N__26727),
            .I(N__26653));
    InMux I__4067 (
            .O(N__26726),
            .I(N__26648));
    InMux I__4066 (
            .O(N__26725),
            .I(N__26648));
    InMux I__4065 (
            .O(N__26724),
            .I(N__26645));
    LocalMux I__4064 (
            .O(N__26717),
            .I(N__26642));
    LocalMux I__4063 (
            .O(N__26714),
            .I(N__26637));
    LocalMux I__4062 (
            .O(N__26711),
            .I(N__26637));
    Span4Mux_v I__4061 (
            .O(N__26708),
            .I(N__26622));
    LocalMux I__4060 (
            .O(N__26705),
            .I(N__26622));
    Span4Mux_v I__4059 (
            .O(N__26700),
            .I(N__26622));
    LocalMux I__4058 (
            .O(N__26693),
            .I(N__26622));
    LocalMux I__4057 (
            .O(N__26686),
            .I(N__26622));
    LocalMux I__4056 (
            .O(N__26681),
            .I(N__26622));
    Span4Mux_v I__4055 (
            .O(N__26674),
            .I(N__26622));
    LocalMux I__4054 (
            .O(N__26669),
            .I(N__26615));
    Span4Mux_h I__4053 (
            .O(N__26662),
            .I(N__26615));
    LocalMux I__4052 (
            .O(N__26659),
            .I(N__26615));
    Odrv12 I__4051 (
            .O(N__26656),
            .I(adc_state_2_adj_1481));
    Odrv4 I__4050 (
            .O(N__26653),
            .I(adc_state_2_adj_1481));
    LocalMux I__4049 (
            .O(N__26648),
            .I(adc_state_2_adj_1481));
    LocalMux I__4048 (
            .O(N__26645),
            .I(adc_state_2_adj_1481));
    Odrv4 I__4047 (
            .O(N__26642),
            .I(adc_state_2_adj_1481));
    Odrv4 I__4046 (
            .O(N__26637),
            .I(adc_state_2_adj_1481));
    Odrv4 I__4045 (
            .O(N__26622),
            .I(adc_state_2_adj_1481));
    Odrv4 I__4044 (
            .O(N__26615),
            .I(adc_state_2_adj_1481));
    InMux I__4043 (
            .O(N__26598),
            .I(N__26586));
    CascadeMux I__4042 (
            .O(N__26597),
            .I(N__26581));
    InMux I__4041 (
            .O(N__26596),
            .I(N__26577));
    InMux I__4040 (
            .O(N__26595),
            .I(N__26572));
    InMux I__4039 (
            .O(N__26594),
            .I(N__26572));
    InMux I__4038 (
            .O(N__26593),
            .I(N__26569));
    InMux I__4037 (
            .O(N__26592),
            .I(N__26566));
    CascadeMux I__4036 (
            .O(N__26591),
            .I(N__26562));
    InMux I__4035 (
            .O(N__26590),
            .I(N__26554));
    InMux I__4034 (
            .O(N__26589),
            .I(N__26554));
    LocalMux I__4033 (
            .O(N__26586),
            .I(N__26551));
    CascadeMux I__4032 (
            .O(N__26585),
            .I(N__26548));
    CascadeMux I__4031 (
            .O(N__26584),
            .I(N__26545));
    InMux I__4030 (
            .O(N__26581),
            .I(N__26536));
    InMux I__4029 (
            .O(N__26580),
            .I(N__26536));
    LocalMux I__4028 (
            .O(N__26577),
            .I(N__26530));
    LocalMux I__4027 (
            .O(N__26572),
            .I(N__26527));
    LocalMux I__4026 (
            .O(N__26569),
            .I(N__26522));
    LocalMux I__4025 (
            .O(N__26566),
            .I(N__26522));
    InMux I__4024 (
            .O(N__26565),
            .I(N__26513));
    InMux I__4023 (
            .O(N__26562),
            .I(N__26513));
    InMux I__4022 (
            .O(N__26561),
            .I(N__26513));
    InMux I__4021 (
            .O(N__26560),
            .I(N__26513));
    InMux I__4020 (
            .O(N__26559),
            .I(N__26510));
    LocalMux I__4019 (
            .O(N__26554),
            .I(N__26505));
    Span4Mux_h I__4018 (
            .O(N__26551),
            .I(N__26505));
    InMux I__4017 (
            .O(N__26548),
            .I(N__26498));
    InMux I__4016 (
            .O(N__26545),
            .I(N__26498));
    InMux I__4015 (
            .O(N__26544),
            .I(N__26498));
    InMux I__4014 (
            .O(N__26543),
            .I(N__26493));
    InMux I__4013 (
            .O(N__26542),
            .I(N__26493));
    InMux I__4012 (
            .O(N__26541),
            .I(N__26490));
    LocalMux I__4011 (
            .O(N__26536),
            .I(N__26487));
    InMux I__4010 (
            .O(N__26535),
            .I(N__26482));
    InMux I__4009 (
            .O(N__26534),
            .I(N__26482));
    InMux I__4008 (
            .O(N__26533),
            .I(N__26479));
    Span4Mux_v I__4007 (
            .O(N__26530),
            .I(N__26470));
    Span4Mux_v I__4006 (
            .O(N__26527),
            .I(N__26470));
    Span4Mux_v I__4005 (
            .O(N__26522),
            .I(N__26470));
    LocalMux I__4004 (
            .O(N__26513),
            .I(N__26470));
    LocalMux I__4003 (
            .O(N__26510),
            .I(N__26463));
    Span4Mux_h I__4002 (
            .O(N__26505),
            .I(N__26463));
    LocalMux I__4001 (
            .O(N__26498),
            .I(N__26463));
    LocalMux I__4000 (
            .O(N__26493),
            .I(\RTD.adc_state_1 ));
    LocalMux I__3999 (
            .O(N__26490),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__3998 (
            .O(N__26487),
            .I(\RTD.adc_state_1 ));
    LocalMux I__3997 (
            .O(N__26482),
            .I(\RTD.adc_state_1 ));
    LocalMux I__3996 (
            .O(N__26479),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__3995 (
            .O(N__26470),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__3994 (
            .O(N__26463),
            .I(\RTD.adc_state_1 ));
    CascadeMux I__3993 (
            .O(N__26448),
            .I(N__26444));
    CascadeMux I__3992 (
            .O(N__26447),
            .I(N__26438));
    InMux I__3991 (
            .O(N__26444),
            .I(N__26428));
    CascadeMux I__3990 (
            .O(N__26443),
            .I(N__26422));
    CascadeMux I__3989 (
            .O(N__26442),
            .I(N__26416));
    CascadeMux I__3988 (
            .O(N__26441),
            .I(N__26412));
    InMux I__3987 (
            .O(N__26438),
            .I(N__26409));
    InMux I__3986 (
            .O(N__26437),
            .I(N__26404));
    InMux I__3985 (
            .O(N__26436),
            .I(N__26404));
    InMux I__3984 (
            .O(N__26435),
            .I(N__26401));
    InMux I__3983 (
            .O(N__26434),
            .I(N__26392));
    InMux I__3982 (
            .O(N__26433),
            .I(N__26392));
    InMux I__3981 (
            .O(N__26432),
            .I(N__26392));
    InMux I__3980 (
            .O(N__26431),
            .I(N__26392));
    LocalMux I__3979 (
            .O(N__26428),
            .I(N__26386));
    CascadeMux I__3978 (
            .O(N__26427),
            .I(N__26382));
    InMux I__3977 (
            .O(N__26426),
            .I(N__26373));
    InMux I__3976 (
            .O(N__26425),
            .I(N__26373));
    InMux I__3975 (
            .O(N__26422),
            .I(N__26373));
    CascadeMux I__3974 (
            .O(N__26421),
            .I(N__26370));
    InMux I__3973 (
            .O(N__26420),
            .I(N__26363));
    InMux I__3972 (
            .O(N__26419),
            .I(N__26363));
    InMux I__3971 (
            .O(N__26416),
            .I(N__26363));
    InMux I__3970 (
            .O(N__26415),
            .I(N__26360));
    InMux I__3969 (
            .O(N__26412),
            .I(N__26357));
    LocalMux I__3968 (
            .O(N__26409),
            .I(N__26350));
    LocalMux I__3967 (
            .O(N__26404),
            .I(N__26350));
    LocalMux I__3966 (
            .O(N__26401),
            .I(N__26350));
    LocalMux I__3965 (
            .O(N__26392),
            .I(N__26347));
    CascadeMux I__3964 (
            .O(N__26391),
            .I(N__26344));
    InMux I__3963 (
            .O(N__26390),
            .I(N__26339));
    InMux I__3962 (
            .O(N__26389),
            .I(N__26339));
    Span4Mux_v I__3961 (
            .O(N__26386),
            .I(N__26336));
    InMux I__3960 (
            .O(N__26385),
            .I(N__26333));
    InMux I__3959 (
            .O(N__26382),
            .I(N__26328));
    InMux I__3958 (
            .O(N__26381),
            .I(N__26328));
    InMux I__3957 (
            .O(N__26380),
            .I(N__26325));
    LocalMux I__3956 (
            .O(N__26373),
            .I(N__26322));
    InMux I__3955 (
            .O(N__26370),
            .I(N__26319));
    LocalMux I__3954 (
            .O(N__26363),
            .I(N__26316));
    LocalMux I__3953 (
            .O(N__26360),
            .I(N__26311));
    LocalMux I__3952 (
            .O(N__26357),
            .I(N__26311));
    Span4Mux_v I__3951 (
            .O(N__26350),
            .I(N__26306));
    Span4Mux_v I__3950 (
            .O(N__26347),
            .I(N__26306));
    InMux I__3949 (
            .O(N__26344),
            .I(N__26303));
    LocalMux I__3948 (
            .O(N__26339),
            .I(N__26298));
    Sp12to4 I__3947 (
            .O(N__26336),
            .I(N__26298));
    LocalMux I__3946 (
            .O(N__26333),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3945 (
            .O(N__26328),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3944 (
            .O(N__26325),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__3943 (
            .O(N__26322),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3942 (
            .O(N__26319),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__3941 (
            .O(N__26316),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__3940 (
            .O(N__26311),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__3939 (
            .O(N__26306),
            .I(\RTD.adc_state_3 ));
    LocalMux I__3938 (
            .O(N__26303),
            .I(\RTD.adc_state_3 ));
    Odrv12 I__3937 (
            .O(N__26298),
            .I(\RTD.adc_state_3 ));
    CascadeMux I__3936 (
            .O(N__26277),
            .I(N__26274));
    InMux I__3935 (
            .O(N__26274),
            .I(N__26254));
    InMux I__3934 (
            .O(N__26273),
            .I(N__26248));
    InMux I__3933 (
            .O(N__26272),
            .I(N__26245));
    InMux I__3932 (
            .O(N__26271),
            .I(N__26242));
    InMux I__3931 (
            .O(N__26270),
            .I(N__26235));
    InMux I__3930 (
            .O(N__26269),
            .I(N__26235));
    InMux I__3929 (
            .O(N__26268),
            .I(N__26235));
    InMux I__3928 (
            .O(N__26267),
            .I(N__26225));
    InMux I__3927 (
            .O(N__26266),
            .I(N__26225));
    InMux I__3926 (
            .O(N__26265),
            .I(N__26225));
    InMux I__3925 (
            .O(N__26264),
            .I(N__26222));
    InMux I__3924 (
            .O(N__26263),
            .I(N__26219));
    InMux I__3923 (
            .O(N__26262),
            .I(N__26214));
    InMux I__3922 (
            .O(N__26261),
            .I(N__26214));
    InMux I__3921 (
            .O(N__26260),
            .I(N__26207));
    InMux I__3920 (
            .O(N__26259),
            .I(N__26207));
    InMux I__3919 (
            .O(N__26258),
            .I(N__26207));
    InMux I__3918 (
            .O(N__26257),
            .I(N__26196));
    LocalMux I__3917 (
            .O(N__26254),
            .I(N__26193));
    InMux I__3916 (
            .O(N__26253),
            .I(N__26190));
    InMux I__3915 (
            .O(N__26252),
            .I(N__26184));
    InMux I__3914 (
            .O(N__26251),
            .I(N__26181));
    LocalMux I__3913 (
            .O(N__26248),
            .I(N__26174));
    LocalMux I__3912 (
            .O(N__26245),
            .I(N__26174));
    LocalMux I__3911 (
            .O(N__26242),
            .I(N__26174));
    LocalMux I__3910 (
            .O(N__26235),
            .I(N__26171));
    InMux I__3909 (
            .O(N__26234),
            .I(N__26164));
    InMux I__3908 (
            .O(N__26233),
            .I(N__26164));
    InMux I__3907 (
            .O(N__26232),
            .I(N__26164));
    LocalMux I__3906 (
            .O(N__26225),
            .I(N__26161));
    LocalMux I__3905 (
            .O(N__26222),
            .I(N__26158));
    LocalMux I__3904 (
            .O(N__26219),
            .I(N__26151));
    LocalMux I__3903 (
            .O(N__26214),
            .I(N__26151));
    LocalMux I__3902 (
            .O(N__26207),
            .I(N__26151));
    InMux I__3901 (
            .O(N__26206),
            .I(N__26134));
    InMux I__3900 (
            .O(N__26205),
            .I(N__26134));
    InMux I__3899 (
            .O(N__26204),
            .I(N__26134));
    InMux I__3898 (
            .O(N__26203),
            .I(N__26134));
    InMux I__3897 (
            .O(N__26202),
            .I(N__26134));
    InMux I__3896 (
            .O(N__26201),
            .I(N__26134));
    InMux I__3895 (
            .O(N__26200),
            .I(N__26134));
    InMux I__3894 (
            .O(N__26199),
            .I(N__26134));
    LocalMux I__3893 (
            .O(N__26196),
            .I(N__26131));
    Span4Mux_h I__3892 (
            .O(N__26193),
            .I(N__26126));
    LocalMux I__3891 (
            .O(N__26190),
            .I(N__26126));
    InMux I__3890 (
            .O(N__26189),
            .I(N__26119));
    InMux I__3889 (
            .O(N__26188),
            .I(N__26119));
    InMux I__3888 (
            .O(N__26187),
            .I(N__26119));
    LocalMux I__3887 (
            .O(N__26184),
            .I(N__26112));
    LocalMux I__3886 (
            .O(N__26181),
            .I(N__26112));
    Span4Mux_v I__3885 (
            .O(N__26174),
            .I(N__26112));
    Span4Mux_v I__3884 (
            .O(N__26171),
            .I(N__26101));
    LocalMux I__3883 (
            .O(N__26164),
            .I(N__26101));
    Span4Mux_v I__3882 (
            .O(N__26161),
            .I(N__26101));
    Span4Mux_h I__3881 (
            .O(N__26158),
            .I(N__26101));
    Span4Mux_v I__3880 (
            .O(N__26151),
            .I(N__26101));
    LocalMux I__3879 (
            .O(N__26134),
            .I(\RTD.adc_state_0 ));
    Odrv12 I__3878 (
            .O(N__26131),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3877 (
            .O(N__26126),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3876 (
            .O(N__26119),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3875 (
            .O(N__26112),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3874 (
            .O(N__26101),
            .I(\RTD.adc_state_0 ));
    SRMux I__3873 (
            .O(N__26088),
            .I(N__26085));
    LocalMux I__3872 (
            .O(N__26085),
            .I(N__26082));
    Sp12to4 I__3871 (
            .O(N__26082),
            .I(N__26079));
    Odrv12 I__3870 (
            .O(N__26079),
            .I(\RTD.n15065 ));
    CascadeMux I__3869 (
            .O(N__26076),
            .I(n13087_cascade_));
    InMux I__3868 (
            .O(N__26073),
            .I(N__26070));
    LocalMux I__3867 (
            .O(N__26070),
            .I(N__26067));
    Span4Mux_h I__3866 (
            .O(N__26067),
            .I(N__26063));
    InMux I__3865 (
            .O(N__26066),
            .I(N__26060));
    Odrv4 I__3864 (
            .O(N__26063),
            .I(cmd_rdadcbuf_26));
    LocalMux I__3863 (
            .O(N__26060),
            .I(cmd_rdadcbuf_26));
    InMux I__3862 (
            .O(N__26055),
            .I(N__26052));
    LocalMux I__3861 (
            .O(N__26052),
            .I(N__26048));
    CascadeMux I__3860 (
            .O(N__26051),
            .I(N__26044));
    Span4Mux_h I__3859 (
            .O(N__26048),
            .I(N__26041));
    InMux I__3858 (
            .O(N__26047),
            .I(N__26038));
    InMux I__3857 (
            .O(N__26044),
            .I(N__26035));
    Odrv4 I__3856 (
            .O(N__26041),
            .I(cmd_rdadctmp_22_adj_1457));
    LocalMux I__3855 (
            .O(N__26038),
            .I(cmd_rdadctmp_22_adj_1457));
    LocalMux I__3854 (
            .O(N__26035),
            .I(cmd_rdadctmp_22_adj_1457));
    CascadeMux I__3853 (
            .O(N__26028),
            .I(N__26025));
    InMux I__3852 (
            .O(N__26025),
            .I(N__26021));
    CascadeMux I__3851 (
            .O(N__26024),
            .I(N__26018));
    LocalMux I__3850 (
            .O(N__26021),
            .I(N__26015));
    InMux I__3849 (
            .O(N__26018),
            .I(N__26012));
    Span4Mux_h I__3848 (
            .O(N__26015),
            .I(N__26009));
    LocalMux I__3847 (
            .O(N__26012),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    Odrv4 I__3846 (
            .O(N__26009),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    CEMux I__3845 (
            .O(N__26004),
            .I(N__26001));
    LocalMux I__3844 (
            .O(N__26001),
            .I(N__25998));
    Span4Mux_h I__3843 (
            .O(N__25998),
            .I(N__25995));
    Odrv4 I__3842 (
            .O(N__25995),
            .I(\ADC_VDC.n12899 ));
    SRMux I__3841 (
            .O(N__25992),
            .I(N__25989));
    LocalMux I__3840 (
            .O(N__25989),
            .I(N__25986));
    Odrv12 I__3839 (
            .O(N__25986),
            .I(\ADC_VDC.n20656 ));
    InMux I__3838 (
            .O(N__25983),
            .I(N__25980));
    LocalMux I__3837 (
            .O(N__25980),
            .I(\comm_spi.n22860 ));
    CascadeMux I__3836 (
            .O(N__25977),
            .I(\comm_spi.n22860_cascade_ ));
    InMux I__3835 (
            .O(N__25974),
            .I(N__25971));
    LocalMux I__3834 (
            .O(N__25971),
            .I(N__25968));
    Odrv4 I__3833 (
            .O(N__25968),
            .I(\comm_spi.n14597 ));
    InMux I__3832 (
            .O(N__25965),
            .I(N__25961));
    CascadeMux I__3831 (
            .O(N__25964),
            .I(N__25958));
    LocalMux I__3830 (
            .O(N__25961),
            .I(N__25955));
    InMux I__3829 (
            .O(N__25958),
            .I(N__25952));
    Odrv4 I__3828 (
            .O(N__25955),
            .I(buf_adcdata_vdc_0));
    LocalMux I__3827 (
            .O(N__25952),
            .I(buf_adcdata_vdc_0));
    CascadeMux I__3826 (
            .O(N__25947),
            .I(n19_adj_1484_cascade_));
    CascadeMux I__3825 (
            .O(N__25944),
            .I(n22_adj_1483_cascade_));
    CascadeMux I__3824 (
            .O(N__25941),
            .I(N__25937));
    CascadeMux I__3823 (
            .O(N__25940),
            .I(N__25933));
    InMux I__3822 (
            .O(N__25937),
            .I(N__25930));
    CascadeMux I__3821 (
            .O(N__25936),
            .I(N__25926));
    InMux I__3820 (
            .O(N__25933),
            .I(N__25923));
    LocalMux I__3819 (
            .O(N__25930),
            .I(N__25919));
    InMux I__3818 (
            .O(N__25929),
            .I(N__25914));
    InMux I__3817 (
            .O(N__25926),
            .I(N__25914));
    LocalMux I__3816 (
            .O(N__25923),
            .I(N__25911));
    CascadeMux I__3815 (
            .O(N__25922),
            .I(N__25908));
    Span4Mux_v I__3814 (
            .O(N__25919),
            .I(N__25905));
    LocalMux I__3813 (
            .O(N__25914),
            .I(N__25902));
    Span4Mux_v I__3812 (
            .O(N__25911),
            .I(N__25899));
    InMux I__3811 (
            .O(N__25908),
            .I(N__25896));
    Span4Mux_h I__3810 (
            .O(N__25905),
            .I(N__25891));
    Span4Mux_v I__3809 (
            .O(N__25902),
            .I(N__25891));
    Sp12to4 I__3808 (
            .O(N__25899),
            .I(N__25884));
    LocalMux I__3807 (
            .O(N__25896),
            .I(N__25884));
    Sp12to4 I__3806 (
            .O(N__25891),
            .I(N__25884));
    Span12Mux_h I__3805 (
            .O(N__25884),
            .I(N__25881));
    Odrv12 I__3804 (
            .O(N__25881),
            .I(IAC_DRDY));
    CEMux I__3803 (
            .O(N__25878),
            .I(N__25874));
    InMux I__3802 (
            .O(N__25877),
            .I(N__25871));
    LocalMux I__3801 (
            .O(N__25874),
            .I(N__25868));
    LocalMux I__3800 (
            .O(N__25871),
            .I(N__25865));
    Span4Mux_h I__3799 (
            .O(N__25868),
            .I(N__25862));
    Span4Mux_h I__3798 (
            .O(N__25865),
            .I(N__25859));
    Odrv4 I__3797 (
            .O(N__25862),
            .I(\ADC_IAC.n12473 ));
    Odrv4 I__3796 (
            .O(N__25859),
            .I(\ADC_IAC.n12473 ));
    CascadeMux I__3795 (
            .O(N__25854),
            .I(\ADC_VDC.n11676_cascade_ ));
    IoInMux I__3794 (
            .O(N__25851),
            .I(N__25848));
    LocalMux I__3793 (
            .O(N__25848),
            .I(N__25845));
    IoSpan4Mux I__3792 (
            .O(N__25845),
            .I(N__25842));
    Span4Mux_s3_h I__3791 (
            .O(N__25842),
            .I(N__25839));
    Span4Mux_h I__3790 (
            .O(N__25839),
            .I(N__25836));
    Span4Mux_h I__3789 (
            .O(N__25836),
            .I(N__25832));
    InMux I__3788 (
            .O(N__25835),
            .I(N__25829));
    Odrv4 I__3787 (
            .O(N__25832),
            .I(VDC_SCLK));
    LocalMux I__3786 (
            .O(N__25829),
            .I(VDC_SCLK));
    SRMux I__3785 (
            .O(N__25824),
            .I(N__25821));
    LocalMux I__3784 (
            .O(N__25821),
            .I(N__25818));
    Span4Mux_h I__3783 (
            .O(N__25818),
            .I(N__25815));
    Odrv4 I__3782 (
            .O(N__25815),
            .I(\comm_spi.iclk_N_763 ));
    InMux I__3781 (
            .O(N__25812),
            .I(N__25809));
    LocalMux I__3780 (
            .O(N__25809),
            .I(N__25806));
    Span4Mux_v I__3779 (
            .O(N__25806),
            .I(N__25803));
    Span4Mux_v I__3778 (
            .O(N__25803),
            .I(N__25799));
    InMux I__3777 (
            .O(N__25802),
            .I(N__25796));
    Odrv4 I__3776 (
            .O(N__25799),
            .I(cmd_rdadcbuf_33));
    LocalMux I__3775 (
            .O(N__25796),
            .I(cmd_rdadcbuf_33));
    InMux I__3774 (
            .O(N__25791),
            .I(N__25788));
    LocalMux I__3773 (
            .O(N__25788),
            .I(N__25785));
    Span4Mux_v I__3772 (
            .O(N__25785),
            .I(N__25781));
    InMux I__3771 (
            .O(N__25784),
            .I(N__25778));
    Odrv4 I__3770 (
            .O(N__25781),
            .I(cmd_rdadcbuf_11));
    LocalMux I__3769 (
            .O(N__25778),
            .I(cmd_rdadcbuf_11));
    CascadeMux I__3768 (
            .O(N__25773),
            .I(N__25770));
    InMux I__3767 (
            .O(N__25770),
            .I(N__25767));
    LocalMux I__3766 (
            .O(N__25767),
            .I(N__25764));
    Span4Mux_v I__3765 (
            .O(N__25764),
            .I(N__25760));
    InMux I__3764 (
            .O(N__25763),
            .I(N__25757));
    Odrv4 I__3763 (
            .O(N__25760),
            .I(cmd_rdadcbuf_21));
    LocalMux I__3762 (
            .O(N__25757),
            .I(cmd_rdadcbuf_21));
    CascadeMux I__3761 (
            .O(N__25752),
            .I(N__25737));
    InMux I__3760 (
            .O(N__25751),
            .I(N__25720));
    InMux I__3759 (
            .O(N__25750),
            .I(N__25720));
    InMux I__3758 (
            .O(N__25749),
            .I(N__25720));
    InMux I__3757 (
            .O(N__25748),
            .I(N__25720));
    InMux I__3756 (
            .O(N__25747),
            .I(N__25720));
    InMux I__3755 (
            .O(N__25746),
            .I(N__25720));
    InMux I__3754 (
            .O(N__25745),
            .I(N__25720));
    InMux I__3753 (
            .O(N__25744),
            .I(N__25709));
    InMux I__3752 (
            .O(N__25743),
            .I(N__25709));
    InMux I__3751 (
            .O(N__25742),
            .I(N__25709));
    InMux I__3750 (
            .O(N__25741),
            .I(N__25709));
    InMux I__3749 (
            .O(N__25740),
            .I(N__25709));
    InMux I__3748 (
            .O(N__25737),
            .I(N__25702));
    InMux I__3747 (
            .O(N__25736),
            .I(N__25702));
    InMux I__3746 (
            .O(N__25735),
            .I(N__25702));
    LocalMux I__3745 (
            .O(N__25720),
            .I(N__25698));
    LocalMux I__3744 (
            .O(N__25709),
            .I(N__25695));
    LocalMux I__3743 (
            .O(N__25702),
            .I(N__25692));
    InMux I__3742 (
            .O(N__25701),
            .I(N__25689));
    Span4Mux_v I__3741 (
            .O(N__25698),
            .I(N__25679));
    Span4Mux_h I__3740 (
            .O(N__25695),
            .I(N__25676));
    Span4Mux_h I__3739 (
            .O(N__25692),
            .I(N__25673));
    LocalMux I__3738 (
            .O(N__25689),
            .I(N__25670));
    InMux I__3737 (
            .O(N__25688),
            .I(N__25665));
    InMux I__3736 (
            .O(N__25687),
            .I(N__25665));
    InMux I__3735 (
            .O(N__25686),
            .I(N__25660));
    InMux I__3734 (
            .O(N__25685),
            .I(N__25660));
    InMux I__3733 (
            .O(N__25684),
            .I(N__25653));
    InMux I__3732 (
            .O(N__25683),
            .I(N__25653));
    InMux I__3731 (
            .O(N__25682),
            .I(N__25653));
    Odrv4 I__3730 (
            .O(N__25679),
            .I(n13087));
    Odrv4 I__3729 (
            .O(N__25676),
            .I(n13087));
    Odrv4 I__3728 (
            .O(N__25673),
            .I(n13087));
    Odrv4 I__3727 (
            .O(N__25670),
            .I(n13087));
    LocalMux I__3726 (
            .O(N__25665),
            .I(n13087));
    LocalMux I__3725 (
            .O(N__25660),
            .I(n13087));
    LocalMux I__3724 (
            .O(N__25653),
            .I(n13087));
    CascadeMux I__3723 (
            .O(N__25638),
            .I(\ADC_IAC.n20960_cascade_ ));
    CEMux I__3722 (
            .O(N__25635),
            .I(N__25632));
    LocalMux I__3721 (
            .O(N__25632),
            .I(N__25629));
    Span4Mux_h I__3720 (
            .O(N__25629),
            .I(N__25626));
    Odrv4 I__3719 (
            .O(N__25626),
            .I(\ADC_IAC.n20961 ));
    InMux I__3718 (
            .O(N__25623),
            .I(N__25619));
    InMux I__3717 (
            .O(N__25622),
            .I(N__25616));
    LocalMux I__3716 (
            .O(N__25619),
            .I(\ADC_IAC.bit_cnt_2 ));
    LocalMux I__3715 (
            .O(N__25616),
            .I(\ADC_IAC.bit_cnt_2 ));
    InMux I__3714 (
            .O(N__25611),
            .I(N__25607));
    InMux I__3713 (
            .O(N__25610),
            .I(N__25604));
    LocalMux I__3712 (
            .O(N__25607),
            .I(\ADC_IAC.bit_cnt_5 ));
    LocalMux I__3711 (
            .O(N__25604),
            .I(\ADC_IAC.bit_cnt_5 ));
    CascadeMux I__3710 (
            .O(N__25599),
            .I(N__25595));
    InMux I__3709 (
            .O(N__25598),
            .I(N__25592));
    InMux I__3708 (
            .O(N__25595),
            .I(N__25589));
    LocalMux I__3707 (
            .O(N__25592),
            .I(\ADC_IAC.bit_cnt_3 ));
    LocalMux I__3706 (
            .O(N__25589),
            .I(\ADC_IAC.bit_cnt_3 ));
    InMux I__3705 (
            .O(N__25584),
            .I(N__25580));
    InMux I__3704 (
            .O(N__25583),
            .I(N__25577));
    LocalMux I__3703 (
            .O(N__25580),
            .I(\ADC_IAC.bit_cnt_4 ));
    LocalMux I__3702 (
            .O(N__25577),
            .I(\ADC_IAC.bit_cnt_4 ));
    InMux I__3701 (
            .O(N__25572),
            .I(N__25568));
    InMux I__3700 (
            .O(N__25571),
            .I(N__25565));
    LocalMux I__3699 (
            .O(N__25568),
            .I(\ADC_IAC.bit_cnt_1 ));
    LocalMux I__3698 (
            .O(N__25565),
            .I(\ADC_IAC.bit_cnt_1 ));
    InMux I__3697 (
            .O(N__25560),
            .I(N__25556));
    InMux I__3696 (
            .O(N__25559),
            .I(N__25553));
    LocalMux I__3695 (
            .O(N__25556),
            .I(N__25550));
    LocalMux I__3694 (
            .O(N__25553),
            .I(\ADC_IAC.bit_cnt_7 ));
    Odrv4 I__3693 (
            .O(N__25550),
            .I(\ADC_IAC.bit_cnt_7 ));
    CascadeMux I__3692 (
            .O(N__25545),
            .I(\ADC_IAC.n21295_cascade_ ));
    InMux I__3691 (
            .O(N__25542),
            .I(N__25539));
    LocalMux I__3690 (
            .O(N__25539),
            .I(\ADC_IAC.n21294 ));
    InMux I__3689 (
            .O(N__25536),
            .I(N__25532));
    InMux I__3688 (
            .O(N__25535),
            .I(N__25529));
    LocalMux I__3687 (
            .O(N__25532),
            .I(\ADC_VAC.bit_cnt_4 ));
    LocalMux I__3686 (
            .O(N__25529),
            .I(\ADC_VAC.bit_cnt_4 ));
    InMux I__3685 (
            .O(N__25524),
            .I(N__25520));
    InMux I__3684 (
            .O(N__25523),
            .I(N__25517));
    LocalMux I__3683 (
            .O(N__25520),
            .I(\ADC_VAC.bit_cnt_3 ));
    LocalMux I__3682 (
            .O(N__25517),
            .I(\ADC_VAC.bit_cnt_3 ));
    CascadeMux I__3681 (
            .O(N__25512),
            .I(N__25508));
    InMux I__3680 (
            .O(N__25511),
            .I(N__25505));
    InMux I__3679 (
            .O(N__25508),
            .I(N__25502));
    LocalMux I__3678 (
            .O(N__25505),
            .I(\ADC_VAC.bit_cnt_1 ));
    LocalMux I__3677 (
            .O(N__25502),
            .I(\ADC_VAC.bit_cnt_1 ));
    InMux I__3676 (
            .O(N__25497),
            .I(N__25493));
    InMux I__3675 (
            .O(N__25496),
            .I(N__25490));
    LocalMux I__3674 (
            .O(N__25493),
            .I(\ADC_VAC.bit_cnt_2 ));
    LocalMux I__3673 (
            .O(N__25490),
            .I(\ADC_VAC.bit_cnt_2 ));
    InMux I__3672 (
            .O(N__25485),
            .I(N__25481));
    InMux I__3671 (
            .O(N__25484),
            .I(N__25478));
    LocalMux I__3670 (
            .O(N__25481),
            .I(\ADC_VAC.bit_cnt_0 ));
    LocalMux I__3669 (
            .O(N__25478),
            .I(\ADC_VAC.bit_cnt_0 ));
    InMux I__3668 (
            .O(N__25473),
            .I(N__25469));
    InMux I__3667 (
            .O(N__25472),
            .I(N__25466));
    LocalMux I__3666 (
            .O(N__25469),
            .I(\ADC_VAC.bit_cnt_6 ));
    LocalMux I__3665 (
            .O(N__25466),
            .I(\ADC_VAC.bit_cnt_6 ));
    CascadeMux I__3664 (
            .O(N__25461),
            .I(\ADC_VAC.n21029_cascade_ ));
    InMux I__3663 (
            .O(N__25458),
            .I(N__25454));
    InMux I__3662 (
            .O(N__25457),
            .I(N__25451));
    LocalMux I__3661 (
            .O(N__25454),
            .I(\ADC_VAC.bit_cnt_7 ));
    LocalMux I__3660 (
            .O(N__25451),
            .I(\ADC_VAC.bit_cnt_7 ));
    InMux I__3659 (
            .O(N__25446),
            .I(N__25443));
    LocalMux I__3658 (
            .O(N__25443),
            .I(N__25440));
    Odrv4 I__3657 (
            .O(N__25440),
            .I(\ADC_VAC.n21043 ));
    CascadeMux I__3656 (
            .O(N__25437),
            .I(N__25433));
    InMux I__3655 (
            .O(N__25436),
            .I(N__25430));
    InMux I__3654 (
            .O(N__25433),
            .I(N__25427));
    LocalMux I__3653 (
            .O(N__25430),
            .I(\ADC_IAC.bit_cnt_6 ));
    LocalMux I__3652 (
            .O(N__25427),
            .I(\ADC_IAC.bit_cnt_6 ));
    InMux I__3651 (
            .O(N__25422),
            .I(N__25418));
    InMux I__3650 (
            .O(N__25421),
            .I(N__25415));
    LocalMux I__3649 (
            .O(N__25418),
            .I(\ADC_IAC.bit_cnt_0 ));
    LocalMux I__3648 (
            .O(N__25415),
            .I(\ADC_IAC.bit_cnt_0 ));
    InMux I__3647 (
            .O(N__25410),
            .I(N__25407));
    LocalMux I__3646 (
            .O(N__25407),
            .I(\ADC_IAC.n16 ));
    InMux I__3645 (
            .O(N__25404),
            .I(N__25399));
    InMux I__3644 (
            .O(N__25403),
            .I(N__25396));
    CascadeMux I__3643 (
            .O(N__25402),
            .I(N__25393));
    LocalMux I__3642 (
            .O(N__25399),
            .I(N__25386));
    LocalMux I__3641 (
            .O(N__25396),
            .I(N__25386));
    InMux I__3640 (
            .O(N__25393),
            .I(N__25383));
    InMux I__3639 (
            .O(N__25392),
            .I(N__25380));
    InMux I__3638 (
            .O(N__25391),
            .I(N__25377));
    Span4Mux_h I__3637 (
            .O(N__25386),
            .I(N__25374));
    LocalMux I__3636 (
            .O(N__25383),
            .I(acadc_trig));
    LocalMux I__3635 (
            .O(N__25380),
            .I(acadc_trig));
    LocalMux I__3634 (
            .O(N__25377),
            .I(acadc_trig));
    Odrv4 I__3633 (
            .O(N__25374),
            .I(acadc_trig));
    IoInMux I__3632 (
            .O(N__25365),
            .I(N__25362));
    LocalMux I__3631 (
            .O(N__25362),
            .I(N__25359));
    Span4Mux_s1_h I__3630 (
            .O(N__25359),
            .I(N__25356));
    Sp12to4 I__3629 (
            .O(N__25356),
            .I(N__25353));
    Span12Mux_s11_v I__3628 (
            .O(N__25353),
            .I(N__25348));
    InMux I__3627 (
            .O(N__25352),
            .I(N__25343));
    InMux I__3626 (
            .O(N__25351),
            .I(N__25343));
    Odrv12 I__3625 (
            .O(N__25348),
            .I(VAC_FLT1));
    LocalMux I__3624 (
            .O(N__25343),
            .I(VAC_FLT1));
    InMux I__3623 (
            .O(N__25338),
            .I(bfn_9_16_0_));
    InMux I__3622 (
            .O(N__25335),
            .I(\ADC_VAC.n19656 ));
    InMux I__3621 (
            .O(N__25332),
            .I(\ADC_VAC.n19657 ));
    InMux I__3620 (
            .O(N__25329),
            .I(\ADC_VAC.n19658 ));
    InMux I__3619 (
            .O(N__25326),
            .I(\ADC_VAC.n19659 ));
    CascadeMux I__3618 (
            .O(N__25323),
            .I(N__25320));
    InMux I__3617 (
            .O(N__25320),
            .I(N__25317));
    LocalMux I__3616 (
            .O(N__25317),
            .I(N__25313));
    InMux I__3615 (
            .O(N__25316),
            .I(N__25310));
    Sp12to4 I__3614 (
            .O(N__25313),
            .I(N__25307));
    LocalMux I__3613 (
            .O(N__25310),
            .I(N__25302));
    Span12Mux_s10_v I__3612 (
            .O(N__25307),
            .I(N__25302));
    Odrv12 I__3611 (
            .O(N__25302),
            .I(\ADC_VAC.bit_cnt_5 ));
    InMux I__3610 (
            .O(N__25299),
            .I(\ADC_VAC.n19660 ));
    InMux I__3609 (
            .O(N__25296),
            .I(\ADC_VAC.n19661 ));
    InMux I__3608 (
            .O(N__25293),
            .I(\ADC_VAC.n19662 ));
    InMux I__3607 (
            .O(N__25290),
            .I(N__25287));
    LocalMux I__3606 (
            .O(N__25287),
            .I(N__25283));
    InMux I__3605 (
            .O(N__25286),
            .I(N__25279));
    Span4Mux_v I__3604 (
            .O(N__25283),
            .I(N__25276));
    CascadeMux I__3603 (
            .O(N__25282),
            .I(N__25273));
    LocalMux I__3602 (
            .O(N__25279),
            .I(N__25270));
    Sp12to4 I__3601 (
            .O(N__25276),
            .I(N__25267));
    InMux I__3600 (
            .O(N__25273),
            .I(N__25264));
    Span4Mux_v I__3599 (
            .O(N__25270),
            .I(N__25261));
    Span12Mux_h I__3598 (
            .O(N__25267),
            .I(N__25258));
    LocalMux I__3597 (
            .O(N__25264),
            .I(buf_adcdata_vac_19));
    Odrv4 I__3596 (
            .O(N__25261),
            .I(buf_adcdata_vac_19));
    Odrv12 I__3595 (
            .O(N__25258),
            .I(buf_adcdata_vac_19));
    InMux I__3594 (
            .O(N__25251),
            .I(N__25248));
    LocalMux I__3593 (
            .O(N__25248),
            .I(N__25245));
    Odrv4 I__3592 (
            .O(N__25245),
            .I(n22435));
    CascadeMux I__3591 (
            .O(N__25242),
            .I(N__25239));
    InMux I__3590 (
            .O(N__25239),
            .I(N__25236));
    LocalMux I__3589 (
            .O(N__25236),
            .I(N__25232));
    CascadeMux I__3588 (
            .O(N__25235),
            .I(N__25229));
    Span4Mux_v I__3587 (
            .O(N__25232),
            .I(N__25226));
    InMux I__3586 (
            .O(N__25229),
            .I(N__25223));
    Odrv4 I__3585 (
            .O(N__25226),
            .I(buf_adcdata_vdc_19));
    LocalMux I__3584 (
            .O(N__25223),
            .I(buf_adcdata_vdc_19));
    InMux I__3583 (
            .O(N__25218),
            .I(N__25212));
    InMux I__3582 (
            .O(N__25217),
            .I(N__25212));
    LocalMux I__3581 (
            .O(N__25212),
            .I(N__25209));
    Odrv4 I__3580 (
            .O(N__25209),
            .I(cmd_rdadctmp_31));
    InMux I__3579 (
            .O(N__25206),
            .I(N__25202));
    CascadeMux I__3578 (
            .O(N__25205),
            .I(N__25198));
    LocalMux I__3577 (
            .O(N__25202),
            .I(N__25195));
    InMux I__3576 (
            .O(N__25201),
            .I(N__25190));
    InMux I__3575 (
            .O(N__25198),
            .I(N__25190));
    Odrv4 I__3574 (
            .O(N__25195),
            .I(cmd_rdadctmp_29));
    LocalMux I__3573 (
            .O(N__25190),
            .I(cmd_rdadctmp_29));
    CascadeMux I__3572 (
            .O(N__25185),
            .I(N__25180));
    CascadeMux I__3571 (
            .O(N__25184),
            .I(N__25177));
    InMux I__3570 (
            .O(N__25183),
            .I(N__25172));
    InMux I__3569 (
            .O(N__25180),
            .I(N__25172));
    InMux I__3568 (
            .O(N__25177),
            .I(N__25169));
    LocalMux I__3567 (
            .O(N__25172),
            .I(cmd_rdadctmp_30));
    LocalMux I__3566 (
            .O(N__25169),
            .I(cmd_rdadctmp_30));
    InMux I__3565 (
            .O(N__25164),
            .I(N__25161));
    LocalMux I__3564 (
            .O(N__25161),
            .I(N__25158));
    Span4Mux_h I__3563 (
            .O(N__25158),
            .I(N__25154));
    CascadeMux I__3562 (
            .O(N__25157),
            .I(N__25151));
    Sp12to4 I__3561 (
            .O(N__25154),
            .I(N__25147));
    InMux I__3560 (
            .O(N__25151),
            .I(N__25144));
    InMux I__3559 (
            .O(N__25150),
            .I(N__25141));
    Span12Mux_v I__3558 (
            .O(N__25147),
            .I(N__25138));
    LocalMux I__3557 (
            .O(N__25144),
            .I(buf_adcdata_iac_23));
    LocalMux I__3556 (
            .O(N__25141),
            .I(buf_adcdata_iac_23));
    Odrv12 I__3555 (
            .O(N__25138),
            .I(buf_adcdata_iac_23));
    InMux I__3554 (
            .O(N__25131),
            .I(N__25128));
    LocalMux I__3553 (
            .O(N__25128),
            .I(N__25123));
    CascadeMux I__3552 (
            .O(N__25127),
            .I(N__25120));
    InMux I__3551 (
            .O(N__25126),
            .I(N__25117));
    Span4Mux_v I__3550 (
            .O(N__25123),
            .I(N__25114));
    InMux I__3549 (
            .O(N__25120),
            .I(N__25111));
    LocalMux I__3548 (
            .O(N__25117),
            .I(cmd_rdadctmp_23));
    Odrv4 I__3547 (
            .O(N__25114),
            .I(cmd_rdadctmp_23));
    LocalMux I__3546 (
            .O(N__25111),
            .I(cmd_rdadctmp_23));
    InMux I__3545 (
            .O(N__25104),
            .I(N__25101));
    LocalMux I__3544 (
            .O(N__25101),
            .I(n22417));
    InMux I__3543 (
            .O(N__25098),
            .I(N__25095));
    LocalMux I__3542 (
            .O(N__25095),
            .I(N__25092));
    Span4Mux_v I__3541 (
            .O(N__25092),
            .I(N__25087));
    CascadeMux I__3540 (
            .O(N__25091),
            .I(N__25084));
    InMux I__3539 (
            .O(N__25090),
            .I(N__25081));
    Sp12to4 I__3538 (
            .O(N__25087),
            .I(N__25078));
    InMux I__3537 (
            .O(N__25084),
            .I(N__25075));
    LocalMux I__3536 (
            .O(N__25081),
            .I(N__25072));
    Span12Mux_h I__3535 (
            .O(N__25078),
            .I(N__25069));
    LocalMux I__3534 (
            .O(N__25075),
            .I(buf_adcdata_vac_20));
    Odrv4 I__3533 (
            .O(N__25072),
            .I(buf_adcdata_vac_20));
    Odrv12 I__3532 (
            .O(N__25069),
            .I(buf_adcdata_vac_20));
    CascadeMux I__3531 (
            .O(N__25062),
            .I(N__25059));
    InMux I__3530 (
            .O(N__25059),
            .I(N__25055));
    CascadeMux I__3529 (
            .O(N__25058),
            .I(N__25052));
    LocalMux I__3528 (
            .O(N__25055),
            .I(N__25049));
    InMux I__3527 (
            .O(N__25052),
            .I(N__25046));
    Odrv12 I__3526 (
            .O(N__25049),
            .I(buf_adcdata_vdc_20));
    LocalMux I__3525 (
            .O(N__25046),
            .I(buf_adcdata_vdc_20));
    CascadeMux I__3524 (
            .O(N__25041),
            .I(N__25038));
    InMux I__3523 (
            .O(N__25038),
            .I(N__25031));
    InMux I__3522 (
            .O(N__25037),
            .I(N__25031));
    CascadeMux I__3521 (
            .O(N__25036),
            .I(N__25028));
    LocalMux I__3520 (
            .O(N__25031),
            .I(N__25025));
    InMux I__3519 (
            .O(N__25028),
            .I(N__25022));
    Odrv4 I__3518 (
            .O(N__25025),
            .I(cmd_rdadctmp_20));
    LocalMux I__3517 (
            .O(N__25022),
            .I(cmd_rdadctmp_20));
    InMux I__3516 (
            .O(N__25017),
            .I(N__25014));
    LocalMux I__3515 (
            .O(N__25014),
            .I(n21139));
    InMux I__3514 (
            .O(N__25011),
            .I(N__25008));
    LocalMux I__3513 (
            .O(N__25008),
            .I(n22291));
    CascadeMux I__3512 (
            .O(N__25005),
            .I(n21138_cascade_));
    InMux I__3511 (
            .O(N__25002),
            .I(N__24999));
    LocalMux I__3510 (
            .O(N__24999),
            .I(N__24994));
    CascadeMux I__3509 (
            .O(N__24998),
            .I(N__24991));
    CascadeMux I__3508 (
            .O(N__24997),
            .I(N__24988));
    Span12Mux_s9_v I__3507 (
            .O(N__24994),
            .I(N__24985));
    InMux I__3506 (
            .O(N__24991),
            .I(N__24982));
    InMux I__3505 (
            .O(N__24988),
            .I(N__24979));
    Span12Mux_h I__3504 (
            .O(N__24985),
            .I(N__24976));
    LocalMux I__3503 (
            .O(N__24982),
            .I(buf_adcdata_iac_21));
    LocalMux I__3502 (
            .O(N__24979),
            .I(buf_adcdata_iac_21));
    Odrv12 I__3501 (
            .O(N__24976),
            .I(buf_adcdata_iac_21));
    InMux I__3500 (
            .O(N__24969),
            .I(N__24966));
    LocalMux I__3499 (
            .O(N__24966),
            .I(N__24962));
    CascadeMux I__3498 (
            .O(N__24965),
            .I(N__24959));
    Span4Mux_v I__3497 (
            .O(N__24962),
            .I(N__24956));
    InMux I__3496 (
            .O(N__24959),
            .I(N__24953));
    Odrv4 I__3495 (
            .O(N__24956),
            .I(buf_adcdata_vdc_13));
    LocalMux I__3494 (
            .O(N__24953),
            .I(buf_adcdata_vdc_13));
    CascadeMux I__3493 (
            .O(N__24948),
            .I(N__24943));
    CascadeMux I__3492 (
            .O(N__24947),
            .I(N__24940));
    InMux I__3491 (
            .O(N__24946),
            .I(N__24937));
    InMux I__3490 (
            .O(N__24943),
            .I(N__24932));
    InMux I__3489 (
            .O(N__24940),
            .I(N__24932));
    LocalMux I__3488 (
            .O(N__24937),
            .I(cmd_rdadctmp_21_adj_1429));
    LocalMux I__3487 (
            .O(N__24932),
            .I(cmd_rdadctmp_21_adj_1429));
    InMux I__3486 (
            .O(N__24927),
            .I(N__24924));
    LocalMux I__3485 (
            .O(N__24924),
            .I(N__24921));
    Span12Mux_v I__3484 (
            .O(N__24921),
            .I(N__24918));
    Span12Mux_h I__3483 (
            .O(N__24918),
            .I(N__24913));
    InMux I__3482 (
            .O(N__24917),
            .I(N__24908));
    InMux I__3481 (
            .O(N__24916),
            .I(N__24908));
    Odrv12 I__3480 (
            .O(N__24913),
            .I(buf_adcdata_vac_13));
    LocalMux I__3479 (
            .O(N__24908),
            .I(buf_adcdata_vac_13));
    InMux I__3478 (
            .O(N__24903),
            .I(N__24898));
    CascadeMux I__3477 (
            .O(N__24902),
            .I(N__24895));
    InMux I__3476 (
            .O(N__24901),
            .I(N__24892));
    LocalMux I__3475 (
            .O(N__24898),
            .I(N__24889));
    InMux I__3474 (
            .O(N__24895),
            .I(N__24886));
    LocalMux I__3473 (
            .O(N__24892),
            .I(cmd_rdadctmp_22_adj_1428));
    Odrv4 I__3472 (
            .O(N__24889),
            .I(cmd_rdadctmp_22_adj_1428));
    LocalMux I__3471 (
            .O(N__24886),
            .I(cmd_rdadctmp_22_adj_1428));
    CascadeMux I__3470 (
            .O(N__24879),
            .I(N__24874));
    InMux I__3469 (
            .O(N__24878),
            .I(N__24871));
    InMux I__3468 (
            .O(N__24877),
            .I(N__24866));
    InMux I__3467 (
            .O(N__24874),
            .I(N__24866));
    LocalMux I__3466 (
            .O(N__24871),
            .I(cmd_rdadctmp_20_adj_1430));
    LocalMux I__3465 (
            .O(N__24866),
            .I(cmd_rdadctmp_20_adj_1430));
    InMux I__3464 (
            .O(N__24861),
            .I(N__24858));
    LocalMux I__3463 (
            .O(N__24858),
            .I(N__24855));
    Span12Mux_v I__3462 (
            .O(N__24855),
            .I(N__24851));
    InMux I__3461 (
            .O(N__24854),
            .I(N__24847));
    Span12Mux_h I__3460 (
            .O(N__24851),
            .I(N__24844));
    InMux I__3459 (
            .O(N__24850),
            .I(N__24841));
    LocalMux I__3458 (
            .O(N__24847),
            .I(buf_adcdata_vac_12));
    Odrv12 I__3457 (
            .O(N__24844),
            .I(buf_adcdata_vac_12));
    LocalMux I__3456 (
            .O(N__24841),
            .I(buf_adcdata_vac_12));
    InMux I__3455 (
            .O(N__24834),
            .I(N__24830));
    InMux I__3454 (
            .O(N__24833),
            .I(N__24827));
    LocalMux I__3453 (
            .O(N__24830),
            .I(N__24823));
    LocalMux I__3452 (
            .O(N__24827),
            .I(N__24820));
    InMux I__3451 (
            .O(N__24826),
            .I(N__24817));
    Span12Mux_s11_h I__3450 (
            .O(N__24823),
            .I(N__24814));
    Span4Mux_h I__3449 (
            .O(N__24820),
            .I(N__24811));
    LocalMux I__3448 (
            .O(N__24817),
            .I(buf_adcdata_iac_7));
    Odrv12 I__3447 (
            .O(N__24814),
            .I(buf_adcdata_iac_7));
    Odrv4 I__3446 (
            .O(N__24811),
            .I(buf_adcdata_iac_7));
    InMux I__3445 (
            .O(N__24804),
            .I(N__24801));
    LocalMux I__3444 (
            .O(N__24801),
            .I(N__24798));
    Odrv4 I__3443 (
            .O(N__24798),
            .I(n19_adj_1623));
    InMux I__3442 (
            .O(N__24795),
            .I(N__24792));
    LocalMux I__3441 (
            .O(N__24792),
            .I(N__24789));
    Span4Mux_v I__3440 (
            .O(N__24789),
            .I(N__24786));
    Span4Mux_h I__3439 (
            .O(N__24786),
            .I(N__24783));
    Odrv4 I__3438 (
            .O(N__24783),
            .I(buf_data_iac_7));
    CascadeMux I__3437 (
            .O(N__24780),
            .I(n22_adj_1624_cascade_));
    InMux I__3436 (
            .O(N__24777),
            .I(N__24767));
    InMux I__3435 (
            .O(N__24776),
            .I(N__24767));
    InMux I__3434 (
            .O(N__24775),
            .I(N__24767));
    InMux I__3433 (
            .O(N__24774),
            .I(N__24764));
    LocalMux I__3432 (
            .O(N__24767),
            .I(N__24758));
    LocalMux I__3431 (
            .O(N__24764),
            .I(N__24758));
    InMux I__3430 (
            .O(N__24763),
            .I(N__24755));
    Span4Mux_v I__3429 (
            .O(N__24758),
            .I(N__24752));
    LocalMux I__3428 (
            .O(N__24755),
            .I(bit_cnt_0_adj_1456));
    Odrv4 I__3427 (
            .O(N__24752),
            .I(bit_cnt_0_adj_1456));
    CascadeMux I__3426 (
            .O(N__24747),
            .I(N__24744));
    InMux I__3425 (
            .O(N__24744),
            .I(N__24740));
    CascadeMux I__3424 (
            .O(N__24743),
            .I(N__24737));
    LocalMux I__3423 (
            .O(N__24740),
            .I(N__24734));
    InMux I__3422 (
            .O(N__24737),
            .I(N__24731));
    Odrv12 I__3421 (
            .O(N__24734),
            .I(cmd_rdadctmp_7));
    LocalMux I__3420 (
            .O(N__24731),
            .I(cmd_rdadctmp_7));
    IoInMux I__3419 (
            .O(N__24726),
            .I(N__24723));
    LocalMux I__3418 (
            .O(N__24723),
            .I(N__24720));
    IoSpan4Mux I__3417 (
            .O(N__24720),
            .I(N__24717));
    Span4Mux_s3_v I__3416 (
            .O(N__24717),
            .I(N__24714));
    Span4Mux_v I__3415 (
            .O(N__24714),
            .I(N__24711));
    Span4Mux_v I__3414 (
            .O(N__24711),
            .I(N__24708));
    Span4Mux_v I__3413 (
            .O(N__24708),
            .I(N__24704));
    InMux I__3412 (
            .O(N__24707),
            .I(N__24701));
    Odrv4 I__3411 (
            .O(N__24704),
            .I(DDS_MOSI1));
    LocalMux I__3410 (
            .O(N__24701),
            .I(DDS_MOSI1));
    CascadeMux I__3409 (
            .O(N__24696),
            .I(N__24693));
    InMux I__3408 (
            .O(N__24693),
            .I(N__24688));
    InMux I__3407 (
            .O(N__24692),
            .I(N__24685));
    InMux I__3406 (
            .O(N__24691),
            .I(N__24682));
    LocalMux I__3405 (
            .O(N__24688),
            .I(N__24679));
    LocalMux I__3404 (
            .O(N__24685),
            .I(N__24675));
    LocalMux I__3403 (
            .O(N__24682),
            .I(N__24672));
    Span4Mux_v I__3402 (
            .O(N__24679),
            .I(N__24668));
    InMux I__3401 (
            .O(N__24678),
            .I(N__24665));
    Span4Mux_h I__3400 (
            .O(N__24675),
            .I(N__24662));
    Span4Mux_v I__3399 (
            .O(N__24672),
            .I(N__24659));
    InMux I__3398 (
            .O(N__24671),
            .I(N__24656));
    Span4Mux_h I__3397 (
            .O(N__24668),
            .I(N__24651));
    LocalMux I__3396 (
            .O(N__24665),
            .I(N__24651));
    Span4Mux_v I__3395 (
            .O(N__24662),
            .I(N__24646));
    Span4Mux_h I__3394 (
            .O(N__24659),
            .I(N__24646));
    LocalMux I__3393 (
            .O(N__24656),
            .I(N__24641));
    Span4Mux_v I__3392 (
            .O(N__24651),
            .I(N__24641));
    Odrv4 I__3391 (
            .O(N__24646),
            .I(buf_cfgRTD_3));
    Odrv4 I__3390 (
            .O(N__24641),
            .I(buf_cfgRTD_3));
    CascadeMux I__3389 (
            .O(N__24636),
            .I(N__24633));
    InMux I__3388 (
            .O(N__24633),
            .I(N__24630));
    LocalMux I__3387 (
            .O(N__24630),
            .I(N__24626));
    CascadeMux I__3386 (
            .O(N__24629),
            .I(N__24623));
    Span4Mux_h I__3385 (
            .O(N__24626),
            .I(N__24620));
    InMux I__3384 (
            .O(N__24623),
            .I(N__24617));
    Odrv4 I__3383 (
            .O(N__24620),
            .I(buf_readRTD_11));
    LocalMux I__3382 (
            .O(N__24617),
            .I(buf_readRTD_11));
    InMux I__3381 (
            .O(N__24612),
            .I(N__24609));
    LocalMux I__3380 (
            .O(N__24609),
            .I(N__24605));
    CascadeMux I__3379 (
            .O(N__24608),
            .I(N__24602));
    Span4Mux_v I__3378 (
            .O(N__24605),
            .I(N__24599));
    InMux I__3377 (
            .O(N__24602),
            .I(N__24596));
    Odrv4 I__3376 (
            .O(N__24599),
            .I(buf_adcdata_vdc_12));
    LocalMux I__3375 (
            .O(N__24596),
            .I(buf_adcdata_vdc_12));
    InMux I__3374 (
            .O(N__24591),
            .I(N__24588));
    LocalMux I__3373 (
            .O(N__24588),
            .I(n19_adj_1511));
    InMux I__3372 (
            .O(N__24585),
            .I(N__24581));
    InMux I__3371 (
            .O(N__24584),
            .I(N__24578));
    LocalMux I__3370 (
            .O(N__24581),
            .I(cmd_rdadcbuf_32));
    LocalMux I__3369 (
            .O(N__24578),
            .I(cmd_rdadcbuf_32));
    InMux I__3368 (
            .O(N__24573),
            .I(N__24570));
    LocalMux I__3367 (
            .O(N__24570),
            .I(N__24566));
    CascadeMux I__3366 (
            .O(N__24569),
            .I(N__24563));
    Span4Mux_v I__3365 (
            .O(N__24566),
            .I(N__24560));
    InMux I__3364 (
            .O(N__24563),
            .I(N__24557));
    Odrv4 I__3363 (
            .O(N__24560),
            .I(buf_adcdata_vdc_21));
    LocalMux I__3362 (
            .O(N__24557),
            .I(buf_adcdata_vdc_21));
    InMux I__3361 (
            .O(N__24552),
            .I(N__24548));
    InMux I__3360 (
            .O(N__24551),
            .I(N__24545));
    LocalMux I__3359 (
            .O(N__24548),
            .I(cmd_rdadcbuf_31));
    LocalMux I__3358 (
            .O(N__24545),
            .I(cmd_rdadcbuf_31));
    InMux I__3357 (
            .O(N__24540),
            .I(N__24536));
    InMux I__3356 (
            .O(N__24539),
            .I(N__24533));
    LocalMux I__3355 (
            .O(N__24536),
            .I(cmd_rdadcbuf_30));
    LocalMux I__3354 (
            .O(N__24533),
            .I(cmd_rdadcbuf_30));
    InMux I__3353 (
            .O(N__24528),
            .I(N__24524));
    InMux I__3352 (
            .O(N__24527),
            .I(N__24521));
    LocalMux I__3351 (
            .O(N__24524),
            .I(cmd_rdadcbuf_29));
    LocalMux I__3350 (
            .O(N__24521),
            .I(cmd_rdadcbuf_29));
    CascadeMux I__3349 (
            .O(N__24516),
            .I(N__24513));
    InMux I__3348 (
            .O(N__24513),
            .I(N__24510));
    LocalMux I__3347 (
            .O(N__24510),
            .I(N__24506));
    CascadeMux I__3346 (
            .O(N__24509),
            .I(N__24502));
    Span4Mux_v I__3345 (
            .O(N__24506),
            .I(N__24499));
    InMux I__3344 (
            .O(N__24505),
            .I(N__24494));
    InMux I__3343 (
            .O(N__24502),
            .I(N__24494));
    Odrv4 I__3342 (
            .O(N__24499),
            .I(cmd_rdadctmp_23_adj_1427));
    LocalMux I__3341 (
            .O(N__24494),
            .I(cmd_rdadctmp_23_adj_1427));
    CascadeMux I__3340 (
            .O(N__24489),
            .I(N__24486));
    InMux I__3339 (
            .O(N__24486),
            .I(N__24481));
    InMux I__3338 (
            .O(N__24485),
            .I(N__24478));
    CascadeMux I__3337 (
            .O(N__24484),
            .I(N__24475));
    LocalMux I__3336 (
            .O(N__24481),
            .I(N__24472));
    LocalMux I__3335 (
            .O(N__24478),
            .I(N__24469));
    InMux I__3334 (
            .O(N__24475),
            .I(N__24466));
    Span4Mux_v I__3333 (
            .O(N__24472),
            .I(N__24463));
    Span4Mux_h I__3332 (
            .O(N__24469),
            .I(N__24460));
    LocalMux I__3331 (
            .O(N__24466),
            .I(cmd_rdadctmp_26_adj_1424));
    Odrv4 I__3330 (
            .O(N__24463),
            .I(cmd_rdadctmp_26_adj_1424));
    Odrv4 I__3329 (
            .O(N__24460),
            .I(cmd_rdadctmp_26_adj_1424));
    CascadeMux I__3328 (
            .O(N__24453),
            .I(N__24449));
    InMux I__3327 (
            .O(N__24452),
            .I(N__24446));
    InMux I__3326 (
            .O(N__24449),
            .I(N__24443));
    LocalMux I__3325 (
            .O(N__24446),
            .I(buf_adcdata_vdc_17));
    LocalMux I__3324 (
            .O(N__24443),
            .I(buf_adcdata_vdc_17));
    CascadeMux I__3323 (
            .O(N__24438),
            .I(N__24435));
    InMux I__3322 (
            .O(N__24435),
            .I(N__24432));
    LocalMux I__3321 (
            .O(N__24432),
            .I(N__24429));
    Span4Mux_h I__3320 (
            .O(N__24429),
            .I(N__24426));
    Odrv4 I__3319 (
            .O(N__24426),
            .I(n22441));
    CascadeMux I__3318 (
            .O(N__24423),
            .I(N__24420));
    InMux I__3317 (
            .O(N__24420),
            .I(N__24417));
    LocalMux I__3316 (
            .O(N__24417),
            .I(N__24413));
    CascadeMux I__3315 (
            .O(N__24416),
            .I(N__24409));
    Span4Mux_h I__3314 (
            .O(N__24413),
            .I(N__24406));
    InMux I__3313 (
            .O(N__24412),
            .I(N__24403));
    InMux I__3312 (
            .O(N__24409),
            .I(N__24400));
    Odrv4 I__3311 (
            .O(N__24406),
            .I(cmd_rdadctmp_25_adj_1425));
    LocalMux I__3310 (
            .O(N__24403),
            .I(cmd_rdadctmp_25_adj_1425));
    LocalMux I__3309 (
            .O(N__24400),
            .I(cmd_rdadctmp_25_adj_1425));
    InMux I__3308 (
            .O(N__24393),
            .I(N__24390));
    LocalMux I__3307 (
            .O(N__24390),
            .I(N__24387));
    Span4Mux_v I__3306 (
            .O(N__24387),
            .I(N__24384));
    Span4Mux_h I__3305 (
            .O(N__24384),
            .I(N__24381));
    Span4Mux_h I__3304 (
            .O(N__24381),
            .I(N__24376));
    InMux I__3303 (
            .O(N__24380),
            .I(N__24371));
    InMux I__3302 (
            .O(N__24379),
            .I(N__24371));
    Odrv4 I__3301 (
            .O(N__24376),
            .I(buf_adcdata_vac_17));
    LocalMux I__3300 (
            .O(N__24371),
            .I(buf_adcdata_vac_17));
    InMux I__3299 (
            .O(N__24366),
            .I(N__24362));
    InMux I__3298 (
            .O(N__24365),
            .I(N__24359));
    LocalMux I__3297 (
            .O(N__24362),
            .I(cmd_rdadcbuf_24));
    LocalMux I__3296 (
            .O(N__24359),
            .I(cmd_rdadcbuf_24));
    InMux I__3295 (
            .O(N__24354),
            .I(N__24351));
    LocalMux I__3294 (
            .O(N__24351),
            .I(N__24347));
    InMux I__3293 (
            .O(N__24350),
            .I(N__24344));
    Odrv4 I__3292 (
            .O(N__24347),
            .I(cmd_rdadcbuf_17));
    LocalMux I__3291 (
            .O(N__24344),
            .I(cmd_rdadcbuf_17));
    InMux I__3290 (
            .O(N__24339),
            .I(N__24336));
    LocalMux I__3289 (
            .O(N__24336),
            .I(N__24333));
    Span4Mux_h I__3288 (
            .O(N__24333),
            .I(N__24329));
    InMux I__3287 (
            .O(N__24332),
            .I(N__24326));
    Odrv4 I__3286 (
            .O(N__24329),
            .I(buf_adcdata_vdc_6));
    LocalMux I__3285 (
            .O(N__24326),
            .I(buf_adcdata_vdc_6));
    InMux I__3284 (
            .O(N__24321),
            .I(N__24317));
    InMux I__3283 (
            .O(N__24320),
            .I(N__24314));
    LocalMux I__3282 (
            .O(N__24317),
            .I(cmd_rdadcbuf_23));
    LocalMux I__3281 (
            .O(N__24314),
            .I(cmd_rdadcbuf_23));
    InMux I__3280 (
            .O(N__24309),
            .I(N__24305));
    InMux I__3279 (
            .O(N__24308),
            .I(N__24302));
    LocalMux I__3278 (
            .O(N__24305),
            .I(buf_adcdata_vdc_7));
    LocalMux I__3277 (
            .O(N__24302),
            .I(buf_adcdata_vdc_7));
    InMux I__3276 (
            .O(N__24297),
            .I(N__24294));
    LocalMux I__3275 (
            .O(N__24294),
            .I(N__24289));
    InMux I__3274 (
            .O(N__24293),
            .I(N__24286));
    InMux I__3273 (
            .O(N__24292),
            .I(N__24283));
    Span4Mux_h I__3272 (
            .O(N__24289),
            .I(N__24280));
    LocalMux I__3271 (
            .O(N__24286),
            .I(N__24277));
    LocalMux I__3270 (
            .O(N__24283),
            .I(buf_adcdata_vac_7));
    Odrv4 I__3269 (
            .O(N__24280),
            .I(buf_adcdata_vac_7));
    Odrv4 I__3268 (
            .O(N__24277),
            .I(buf_adcdata_vac_7));
    InMux I__3267 (
            .O(N__24270),
            .I(N__24266));
    InMux I__3266 (
            .O(N__24269),
            .I(N__24263));
    LocalMux I__3265 (
            .O(N__24266),
            .I(cmd_rdadcbuf_20));
    LocalMux I__3264 (
            .O(N__24263),
            .I(cmd_rdadcbuf_20));
    InMux I__3263 (
            .O(N__24258),
            .I(N__24254));
    InMux I__3262 (
            .O(N__24257),
            .I(N__24251));
    LocalMux I__3261 (
            .O(N__24254),
            .I(cmd_rdadcbuf_22));
    LocalMux I__3260 (
            .O(N__24251),
            .I(cmd_rdadcbuf_22));
    InMux I__3259 (
            .O(N__24246),
            .I(N__24242));
    InMux I__3258 (
            .O(N__24245),
            .I(N__24239));
    LocalMux I__3257 (
            .O(N__24242),
            .I(cmd_rdadcbuf_28));
    LocalMux I__3256 (
            .O(N__24239),
            .I(cmd_rdadcbuf_28));
    InMux I__3255 (
            .O(N__24234),
            .I(N__24230));
    InMux I__3254 (
            .O(N__24233),
            .I(N__24227));
    LocalMux I__3253 (
            .O(N__24230),
            .I(N__24223));
    LocalMux I__3252 (
            .O(N__24227),
            .I(N__24220));
    InMux I__3251 (
            .O(N__24226),
            .I(N__24217));
    Span12Mux_h I__3250 (
            .O(N__24223),
            .I(N__24212));
    Sp12to4 I__3249 (
            .O(N__24220),
            .I(N__24212));
    LocalMux I__3248 (
            .O(N__24217),
            .I(cmd_rdadcbuf_34));
    Odrv12 I__3247 (
            .O(N__24212),
            .I(cmd_rdadcbuf_34));
    CascadeMux I__3246 (
            .O(N__24207),
            .I(N__24203));
    InMux I__3245 (
            .O(N__24206),
            .I(N__24200));
    InMux I__3244 (
            .O(N__24203),
            .I(N__24197));
    LocalMux I__3243 (
            .O(N__24200),
            .I(buf_adcdata_vdc_23));
    LocalMux I__3242 (
            .O(N__24197),
            .I(buf_adcdata_vdc_23));
    InMux I__3241 (
            .O(N__24192),
            .I(N__24189));
    LocalMux I__3240 (
            .O(N__24189),
            .I(N__24186));
    Span12Mux_s8_h I__3239 (
            .O(N__24186),
            .I(N__24181));
    InMux I__3238 (
            .O(N__24185),
            .I(N__24178));
    InMux I__3237 (
            .O(N__24184),
            .I(N__24175));
    Span12Mux_h I__3236 (
            .O(N__24181),
            .I(N__24172));
    LocalMux I__3235 (
            .O(N__24178),
            .I(N__24169));
    LocalMux I__3234 (
            .O(N__24175),
            .I(buf_adcdata_vac_23));
    Odrv12 I__3233 (
            .O(N__24172),
            .I(buf_adcdata_vac_23));
    Odrv4 I__3232 (
            .O(N__24169),
            .I(buf_adcdata_vac_23));
    InMux I__3231 (
            .O(N__24162),
            .I(N__24157));
    CascadeMux I__3230 (
            .O(N__24161),
            .I(N__24154));
    CascadeMux I__3229 (
            .O(N__24160),
            .I(N__24151));
    LocalMux I__3228 (
            .O(N__24157),
            .I(N__24148));
    InMux I__3227 (
            .O(N__24154),
            .I(N__24145));
    InMux I__3226 (
            .O(N__24151),
            .I(N__24142));
    Odrv4 I__3225 (
            .O(N__24148),
            .I(cmd_rdadctmp_5_adj_1474));
    LocalMux I__3224 (
            .O(N__24145),
            .I(cmd_rdadctmp_5_adj_1474));
    LocalMux I__3223 (
            .O(N__24142),
            .I(cmd_rdadctmp_5_adj_1474));
    CascadeMux I__3222 (
            .O(N__24135),
            .I(N__24132));
    InMux I__3221 (
            .O(N__24132),
            .I(N__24128));
    CascadeMux I__3220 (
            .O(N__24131),
            .I(N__24124));
    LocalMux I__3219 (
            .O(N__24128),
            .I(N__24121));
    InMux I__3218 (
            .O(N__24127),
            .I(N__24118));
    InMux I__3217 (
            .O(N__24124),
            .I(N__24115));
    Odrv4 I__3216 (
            .O(N__24121),
            .I(cmd_rdadctmp_6_adj_1473));
    LocalMux I__3215 (
            .O(N__24118),
            .I(cmd_rdadctmp_6_adj_1473));
    LocalMux I__3214 (
            .O(N__24115),
            .I(cmd_rdadctmp_6_adj_1473));
    InMux I__3213 (
            .O(N__24108),
            .I(N__24101));
    InMux I__3212 (
            .O(N__24107),
            .I(N__24101));
    InMux I__3211 (
            .O(N__24106),
            .I(N__24098));
    LocalMux I__3210 (
            .O(N__24101),
            .I(cmd_rdadctmp_7_adj_1472));
    LocalMux I__3209 (
            .O(N__24098),
            .I(cmd_rdadctmp_7_adj_1472));
    InMux I__3208 (
            .O(N__24093),
            .I(N__24089));
    InMux I__3207 (
            .O(N__24092),
            .I(N__24086));
    LocalMux I__3206 (
            .O(N__24089),
            .I(cmd_rdadcbuf_15));
    LocalMux I__3205 (
            .O(N__24086),
            .I(cmd_rdadcbuf_15));
    InMux I__3204 (
            .O(N__24081),
            .I(N__24077));
    CascadeMux I__3203 (
            .O(N__24080),
            .I(N__24074));
    LocalMux I__3202 (
            .O(N__24077),
            .I(N__24071));
    InMux I__3201 (
            .O(N__24074),
            .I(N__24068));
    Odrv4 I__3200 (
            .O(N__24071),
            .I(buf_adcdata_vdc_4));
    LocalMux I__3199 (
            .O(N__24068),
            .I(buf_adcdata_vdc_4));
    InMux I__3198 (
            .O(N__24063),
            .I(N__24058));
    CascadeMux I__3197 (
            .O(N__24062),
            .I(N__24055));
    InMux I__3196 (
            .O(N__24061),
            .I(N__24052));
    LocalMux I__3195 (
            .O(N__24058),
            .I(N__24049));
    InMux I__3194 (
            .O(N__24055),
            .I(N__24046));
    LocalMux I__3193 (
            .O(N__24052),
            .I(cmd_rdadctmp_12_adj_1467));
    Odrv12 I__3192 (
            .O(N__24049),
            .I(cmd_rdadctmp_12_adj_1467));
    LocalMux I__3191 (
            .O(N__24046),
            .I(cmd_rdadctmp_12_adj_1467));
    CascadeMux I__3190 (
            .O(N__24039),
            .I(N__24034));
    InMux I__3189 (
            .O(N__24038),
            .I(N__24031));
    CascadeMux I__3188 (
            .O(N__24037),
            .I(N__24028));
    InMux I__3187 (
            .O(N__24034),
            .I(N__24025));
    LocalMux I__3186 (
            .O(N__24031),
            .I(N__24022));
    InMux I__3185 (
            .O(N__24028),
            .I(N__24019));
    LocalMux I__3184 (
            .O(N__24025),
            .I(cmd_rdadctmp_13_adj_1466));
    Odrv4 I__3183 (
            .O(N__24022),
            .I(cmd_rdadctmp_13_adj_1466));
    LocalMux I__3182 (
            .O(N__24019),
            .I(cmd_rdadctmp_13_adj_1466));
    CascadeMux I__3181 (
            .O(N__24012),
            .I(N__24007));
    CascadeMux I__3180 (
            .O(N__24011),
            .I(N__24004));
    InMux I__3179 (
            .O(N__24010),
            .I(N__24001));
    InMux I__3178 (
            .O(N__24007),
            .I(N__23998));
    InMux I__3177 (
            .O(N__24004),
            .I(N__23995));
    LocalMux I__3176 (
            .O(N__24001),
            .I(cmd_rdadctmp_9_adj_1470));
    LocalMux I__3175 (
            .O(N__23998),
            .I(cmd_rdadctmp_9_adj_1470));
    LocalMux I__3174 (
            .O(N__23995),
            .I(cmd_rdadctmp_9_adj_1470));
    InMux I__3173 (
            .O(N__23988),
            .I(N__23984));
    CascadeMux I__3172 (
            .O(N__23987),
            .I(N__23980));
    LocalMux I__3171 (
            .O(N__23984),
            .I(N__23977));
    InMux I__3170 (
            .O(N__23983),
            .I(N__23974));
    InMux I__3169 (
            .O(N__23980),
            .I(N__23971));
    Odrv4 I__3168 (
            .O(N__23977),
            .I(cmd_rdadctmp_10_adj_1469));
    LocalMux I__3167 (
            .O(N__23974),
            .I(cmd_rdadctmp_10_adj_1469));
    LocalMux I__3166 (
            .O(N__23971),
            .I(cmd_rdadctmp_10_adj_1469));
    InMux I__3165 (
            .O(N__23964),
            .I(N__23961));
    LocalMux I__3164 (
            .O(N__23961),
            .I(N__23957));
    InMux I__3163 (
            .O(N__23960),
            .I(N__23954));
    Odrv4 I__3162 (
            .O(N__23957),
            .I(cmd_rdadcbuf_14));
    LocalMux I__3161 (
            .O(N__23954),
            .I(cmd_rdadcbuf_14));
    InMux I__3160 (
            .O(N__23949),
            .I(N__23945));
    CascadeMux I__3159 (
            .O(N__23948),
            .I(N__23941));
    LocalMux I__3158 (
            .O(N__23945),
            .I(N__23938));
    InMux I__3157 (
            .O(N__23944),
            .I(N__23935));
    InMux I__3156 (
            .O(N__23941),
            .I(N__23932));
    Odrv4 I__3155 (
            .O(N__23938),
            .I(cmd_rdadctmp_15_adj_1464));
    LocalMux I__3154 (
            .O(N__23935),
            .I(cmd_rdadctmp_15_adj_1464));
    LocalMux I__3153 (
            .O(N__23932),
            .I(cmd_rdadctmp_15_adj_1464));
    CascadeMux I__3152 (
            .O(N__23925),
            .I(N__23922));
    InMux I__3151 (
            .O(N__23922),
            .I(N__23918));
    InMux I__3150 (
            .O(N__23921),
            .I(N__23914));
    LocalMux I__3149 (
            .O(N__23918),
            .I(N__23911));
    CascadeMux I__3148 (
            .O(N__23917),
            .I(N__23908));
    LocalMux I__3147 (
            .O(N__23914),
            .I(N__23903));
    Span4Mux_v I__3146 (
            .O(N__23911),
            .I(N__23903));
    InMux I__3145 (
            .O(N__23908),
            .I(N__23900));
    Odrv4 I__3144 (
            .O(N__23903),
            .I(cmd_rdadctmp_16_adj_1463));
    LocalMux I__3143 (
            .O(N__23900),
            .I(cmd_rdadctmp_16_adj_1463));
    CascadeMux I__3142 (
            .O(N__23895),
            .I(N__23884));
    CascadeMux I__3141 (
            .O(N__23894),
            .I(N__23881));
    CascadeMux I__3140 (
            .O(N__23893),
            .I(N__23877));
    CascadeMux I__3139 (
            .O(N__23892),
            .I(N__23873));
    CascadeMux I__3138 (
            .O(N__23891),
            .I(N__23870));
    CascadeMux I__3137 (
            .O(N__23890),
            .I(N__23866));
    CascadeMux I__3136 (
            .O(N__23889),
            .I(N__23863));
    CascadeMux I__3135 (
            .O(N__23888),
            .I(N__23857));
    InMux I__3134 (
            .O(N__23887),
            .I(N__23852));
    InMux I__3133 (
            .O(N__23884),
            .I(N__23852));
    InMux I__3132 (
            .O(N__23881),
            .I(N__23841));
    InMux I__3131 (
            .O(N__23880),
            .I(N__23841));
    InMux I__3130 (
            .O(N__23877),
            .I(N__23841));
    InMux I__3129 (
            .O(N__23876),
            .I(N__23841));
    InMux I__3128 (
            .O(N__23873),
            .I(N__23841));
    InMux I__3127 (
            .O(N__23870),
            .I(N__23820));
    InMux I__3126 (
            .O(N__23869),
            .I(N__23820));
    InMux I__3125 (
            .O(N__23866),
            .I(N__23820));
    InMux I__3124 (
            .O(N__23863),
            .I(N__23820));
    InMux I__3123 (
            .O(N__23862),
            .I(N__23820));
    InMux I__3122 (
            .O(N__23861),
            .I(N__23820));
    InMux I__3121 (
            .O(N__23860),
            .I(N__23820));
    InMux I__3120 (
            .O(N__23857),
            .I(N__23820));
    LocalMux I__3119 (
            .O(N__23852),
            .I(N__23815));
    LocalMux I__3118 (
            .O(N__23841),
            .I(N__23815));
    CascadeMux I__3117 (
            .O(N__23840),
            .I(N__23811));
    CascadeMux I__3116 (
            .O(N__23839),
            .I(N__23808));
    CascadeMux I__3115 (
            .O(N__23838),
            .I(N__23804));
    CascadeMux I__3114 (
            .O(N__23837),
            .I(N__23801));
    LocalMux I__3113 (
            .O(N__23820),
            .I(N__23797));
    Span4Mux_v I__3112 (
            .O(N__23815),
            .I(N__23794));
    InMux I__3111 (
            .O(N__23814),
            .I(N__23787));
    InMux I__3110 (
            .O(N__23811),
            .I(N__23787));
    InMux I__3109 (
            .O(N__23808),
            .I(N__23787));
    InMux I__3108 (
            .O(N__23807),
            .I(N__23784));
    InMux I__3107 (
            .O(N__23804),
            .I(N__23777));
    InMux I__3106 (
            .O(N__23801),
            .I(N__23777));
    InMux I__3105 (
            .O(N__23800),
            .I(N__23777));
    Odrv4 I__3104 (
            .O(N__23797),
            .I(n12871));
    Odrv4 I__3103 (
            .O(N__23794),
            .I(n12871));
    LocalMux I__3102 (
            .O(N__23787),
            .I(n12871));
    LocalMux I__3101 (
            .O(N__23784),
            .I(n12871));
    LocalMux I__3100 (
            .O(N__23777),
            .I(n12871));
    InMux I__3099 (
            .O(N__23766),
            .I(N__23763));
    LocalMux I__3098 (
            .O(N__23763),
            .I(N__23758));
    CascadeMux I__3097 (
            .O(N__23762),
            .I(N__23755));
    InMux I__3096 (
            .O(N__23761),
            .I(N__23752));
    Span4Mux_v I__3095 (
            .O(N__23758),
            .I(N__23749));
    InMux I__3094 (
            .O(N__23755),
            .I(N__23746));
    LocalMux I__3093 (
            .O(N__23752),
            .I(cmd_rdadctmp_18_adj_1461));
    Odrv4 I__3092 (
            .O(N__23749),
            .I(cmd_rdadctmp_18_adj_1461));
    LocalMux I__3091 (
            .O(N__23746),
            .I(cmd_rdadctmp_18_adj_1461));
    InMux I__3090 (
            .O(N__23739),
            .I(N__23736));
    LocalMux I__3089 (
            .O(N__23736),
            .I(N__23731));
    CascadeMux I__3088 (
            .O(N__23735),
            .I(N__23728));
    CascadeMux I__3087 (
            .O(N__23734),
            .I(N__23725));
    Span4Mux_v I__3086 (
            .O(N__23731),
            .I(N__23722));
    InMux I__3085 (
            .O(N__23728),
            .I(N__23719));
    InMux I__3084 (
            .O(N__23725),
            .I(N__23716));
    Odrv4 I__3083 (
            .O(N__23722),
            .I(cmd_rdadctmp_19_adj_1460));
    LocalMux I__3082 (
            .O(N__23719),
            .I(cmd_rdadctmp_19_adj_1460));
    LocalMux I__3081 (
            .O(N__23716),
            .I(cmd_rdadctmp_19_adj_1460));
    InMux I__3080 (
            .O(N__23709),
            .I(N__23706));
    LocalMux I__3079 (
            .O(N__23706),
            .I(N__23702));
    InMux I__3078 (
            .O(N__23705),
            .I(N__23699));
    Odrv4 I__3077 (
            .O(N__23702),
            .I(cmd_rdadcbuf_25));
    LocalMux I__3076 (
            .O(N__23699),
            .I(cmd_rdadcbuf_25));
    InMux I__3075 (
            .O(N__23694),
            .I(N__23691));
    LocalMux I__3074 (
            .O(N__23691),
            .I(N__23687));
    InMux I__3073 (
            .O(N__23690),
            .I(N__23684));
    Odrv4 I__3072 (
            .O(N__23687),
            .I(cmd_rdadcbuf_19));
    LocalMux I__3071 (
            .O(N__23684),
            .I(cmd_rdadcbuf_19));
    InMux I__3070 (
            .O(N__23679),
            .I(N__23676));
    LocalMux I__3069 (
            .O(N__23676),
            .I(N__23673));
    Span4Mux_v I__3068 (
            .O(N__23673),
            .I(N__23669));
    CascadeMux I__3067 (
            .O(N__23672),
            .I(N__23666));
    Span4Mux_v I__3066 (
            .O(N__23669),
            .I(N__23663));
    InMux I__3065 (
            .O(N__23666),
            .I(N__23660));
    Odrv4 I__3064 (
            .O(N__23663),
            .I(buf_adcdata_vdc_8));
    LocalMux I__3063 (
            .O(N__23660),
            .I(buf_adcdata_vdc_8));
    InMux I__3062 (
            .O(N__23655),
            .I(N__23651));
    InMux I__3061 (
            .O(N__23654),
            .I(N__23648));
    LocalMux I__3060 (
            .O(N__23651),
            .I(cmd_rdadcbuf_12));
    LocalMux I__3059 (
            .O(N__23648),
            .I(cmd_rdadcbuf_12));
    InMux I__3058 (
            .O(N__23643),
            .I(N__23639));
    InMux I__3057 (
            .O(N__23642),
            .I(N__23636));
    LocalMux I__3056 (
            .O(N__23639),
            .I(cmd_rdadcbuf_13));
    LocalMux I__3055 (
            .O(N__23636),
            .I(cmd_rdadcbuf_13));
    InMux I__3054 (
            .O(N__23631),
            .I(N__23627));
    CascadeMux I__3053 (
            .O(N__23630),
            .I(N__23623));
    LocalMux I__3052 (
            .O(N__23627),
            .I(N__23620));
    CascadeMux I__3051 (
            .O(N__23626),
            .I(N__23617));
    InMux I__3050 (
            .O(N__23623),
            .I(N__23614));
    Span4Mux_v I__3049 (
            .O(N__23620),
            .I(N__23611));
    InMux I__3048 (
            .O(N__23617),
            .I(N__23608));
    LocalMux I__3047 (
            .O(N__23614),
            .I(cmd_rdadctmp_14_adj_1465));
    Odrv4 I__3046 (
            .O(N__23611),
            .I(cmd_rdadctmp_14_adj_1465));
    LocalMux I__3045 (
            .O(N__23608),
            .I(cmd_rdadctmp_14_adj_1465));
    CascadeMux I__3044 (
            .O(N__23601),
            .I(N__23596));
    InMux I__3043 (
            .O(N__23600),
            .I(N__23593));
    InMux I__3042 (
            .O(N__23599),
            .I(N__23590));
    InMux I__3041 (
            .O(N__23596),
            .I(N__23587));
    LocalMux I__3040 (
            .O(N__23593),
            .I(cmd_rdadctmp_3_adj_1476));
    LocalMux I__3039 (
            .O(N__23590),
            .I(cmd_rdadctmp_3_adj_1476));
    LocalMux I__3038 (
            .O(N__23587),
            .I(cmd_rdadctmp_3_adj_1476));
    CascadeMux I__3037 (
            .O(N__23580),
            .I(N__23575));
    InMux I__3036 (
            .O(N__23579),
            .I(N__23572));
    InMux I__3035 (
            .O(N__23578),
            .I(N__23569));
    InMux I__3034 (
            .O(N__23575),
            .I(N__23566));
    LocalMux I__3033 (
            .O(N__23572),
            .I(cmd_rdadctmp_4_adj_1475));
    LocalMux I__3032 (
            .O(N__23569),
            .I(cmd_rdadctmp_4_adj_1475));
    LocalMux I__3031 (
            .O(N__23566),
            .I(cmd_rdadctmp_4_adj_1475));
    CascadeMux I__3030 (
            .O(N__23559),
            .I(N__23554));
    InMux I__3029 (
            .O(N__23558),
            .I(N__23551));
    InMux I__3028 (
            .O(N__23557),
            .I(N__23548));
    InMux I__3027 (
            .O(N__23554),
            .I(N__23545));
    LocalMux I__3026 (
            .O(N__23551),
            .I(cmd_rdadctmp_8_adj_1471));
    LocalMux I__3025 (
            .O(N__23548),
            .I(cmd_rdadctmp_8_adj_1471));
    LocalMux I__3024 (
            .O(N__23545),
            .I(cmd_rdadctmp_8_adj_1471));
    InMux I__3023 (
            .O(N__23538),
            .I(N__23534));
    InMux I__3022 (
            .O(N__23537),
            .I(N__23531));
    LocalMux I__3021 (
            .O(N__23534),
            .I(cmd_rdadcbuf_18));
    LocalMux I__3020 (
            .O(N__23531),
            .I(cmd_rdadcbuf_18));
    InMux I__3019 (
            .O(N__23526),
            .I(\ADC_IAC.n19654 ));
    InMux I__3018 (
            .O(N__23523),
            .I(\ADC_IAC.n19655 ));
    SRMux I__3017 (
            .O(N__23520),
            .I(N__23517));
    LocalMux I__3016 (
            .O(N__23517),
            .I(N__23514));
    Sp12to4 I__3015 (
            .O(N__23514),
            .I(N__23511));
    Odrv12 I__3014 (
            .O(N__23511),
            .I(\ADC_IAC.n14806 ));
    CascadeMux I__3013 (
            .O(N__23508),
            .I(\ADC_IAC.n17_cascade_ ));
    CEMux I__3012 (
            .O(N__23505),
            .I(N__23502));
    LocalMux I__3011 (
            .O(N__23502),
            .I(\ADC_IAC.n12 ));
    InMux I__3010 (
            .O(N__23499),
            .I(N__23495));
    InMux I__3009 (
            .O(N__23498),
            .I(N__23492));
    LocalMux I__3008 (
            .O(N__23495),
            .I(\ADC_VDC.avg_cnt_4 ));
    LocalMux I__3007 (
            .O(N__23492),
            .I(\ADC_VDC.avg_cnt_4 ));
    InMux I__3006 (
            .O(N__23487),
            .I(N__23483));
    InMux I__3005 (
            .O(N__23486),
            .I(N__23480));
    LocalMux I__3004 (
            .O(N__23483),
            .I(\ADC_VDC.avg_cnt_7 ));
    LocalMux I__3003 (
            .O(N__23480),
            .I(\ADC_VDC.avg_cnt_7 ));
    CascadeMux I__3002 (
            .O(N__23475),
            .I(N__23471));
    InMux I__3001 (
            .O(N__23474),
            .I(N__23468));
    InMux I__3000 (
            .O(N__23471),
            .I(N__23465));
    LocalMux I__2999 (
            .O(N__23468),
            .I(\ADC_VDC.avg_cnt_3 ));
    LocalMux I__2998 (
            .O(N__23465),
            .I(\ADC_VDC.avg_cnt_3 ));
    InMux I__2997 (
            .O(N__23460),
            .I(N__23456));
    InMux I__2996 (
            .O(N__23459),
            .I(N__23453));
    LocalMux I__2995 (
            .O(N__23456),
            .I(\ADC_VDC.avg_cnt_5 ));
    LocalMux I__2994 (
            .O(N__23453),
            .I(\ADC_VDC.avg_cnt_5 ));
    InMux I__2993 (
            .O(N__23448),
            .I(N__23445));
    LocalMux I__2992 (
            .O(N__23445),
            .I(\ADC_VDC.n20 ));
    InMux I__2991 (
            .O(N__23442),
            .I(N__23438));
    InMux I__2990 (
            .O(N__23441),
            .I(N__23435));
    LocalMux I__2989 (
            .O(N__23438),
            .I(\ADC_VDC.avg_cnt_11 ));
    LocalMux I__2988 (
            .O(N__23435),
            .I(\ADC_VDC.avg_cnt_11 ));
    InMux I__2987 (
            .O(N__23430),
            .I(N__23426));
    InMux I__2986 (
            .O(N__23429),
            .I(N__23423));
    LocalMux I__2985 (
            .O(N__23426),
            .I(\ADC_VDC.avg_cnt_2 ));
    LocalMux I__2984 (
            .O(N__23423),
            .I(\ADC_VDC.avg_cnt_2 ));
    CascadeMux I__2983 (
            .O(N__23418),
            .I(N__23414));
    InMux I__2982 (
            .O(N__23417),
            .I(N__23411));
    InMux I__2981 (
            .O(N__23414),
            .I(N__23408));
    LocalMux I__2980 (
            .O(N__23411),
            .I(\ADC_VDC.avg_cnt_1 ));
    LocalMux I__2979 (
            .O(N__23408),
            .I(\ADC_VDC.avg_cnt_1 ));
    InMux I__2978 (
            .O(N__23403),
            .I(N__23399));
    InMux I__2977 (
            .O(N__23402),
            .I(N__23396));
    LocalMux I__2976 (
            .O(N__23399),
            .I(\ADC_VDC.avg_cnt_6 ));
    LocalMux I__2975 (
            .O(N__23396),
            .I(\ADC_VDC.avg_cnt_6 ));
    InMux I__2974 (
            .O(N__23391),
            .I(N__23388));
    LocalMux I__2973 (
            .O(N__23388),
            .I(\ADC_VDC.n21 ));
    InMux I__2972 (
            .O(N__23385),
            .I(N__23382));
    LocalMux I__2971 (
            .O(N__23382),
            .I(N__23379));
    Span4Mux_h I__2970 (
            .O(N__23379),
            .I(N__23375));
    InMux I__2969 (
            .O(N__23378),
            .I(N__23372));
    Odrv4 I__2968 (
            .O(N__23375),
            .I(cmd_rdadcbuf_27));
    LocalMux I__2967 (
            .O(N__23372),
            .I(cmd_rdadcbuf_27));
    InMux I__2966 (
            .O(N__23367),
            .I(N__23364));
    LocalMux I__2965 (
            .O(N__23364),
            .I(N__23360));
    CascadeMux I__2964 (
            .O(N__23363),
            .I(N__23357));
    Sp12to4 I__2963 (
            .O(N__23360),
            .I(N__23354));
    InMux I__2962 (
            .O(N__23357),
            .I(N__23351));
    Odrv12 I__2961 (
            .O(N__23354),
            .I(buf_adcdata_vdc_16));
    LocalMux I__2960 (
            .O(N__23351),
            .I(buf_adcdata_vdc_16));
    CascadeMux I__2959 (
            .O(N__23346),
            .I(N__23343));
    InMux I__2958 (
            .O(N__23343),
            .I(N__23340));
    LocalMux I__2957 (
            .O(N__23340),
            .I(N__23335));
    InMux I__2956 (
            .O(N__23339),
            .I(N__23330));
    InMux I__2955 (
            .O(N__23338),
            .I(N__23330));
    Span4Mux_v I__2954 (
            .O(N__23335),
            .I(N__23327));
    LocalMux I__2953 (
            .O(N__23330),
            .I(cmd_rdadctmp_18));
    Odrv4 I__2952 (
            .O(N__23327),
            .I(cmd_rdadctmp_18));
    IoInMux I__2951 (
            .O(N__23322),
            .I(N__23319));
    LocalMux I__2950 (
            .O(N__23319),
            .I(N__23316));
    IoSpan4Mux I__2949 (
            .O(N__23316),
            .I(N__23313));
    Span4Mux_s3_v I__2948 (
            .O(N__23313),
            .I(N__23310));
    Sp12to4 I__2947 (
            .O(N__23310),
            .I(N__23307));
    Span12Mux_s10_v I__2946 (
            .O(N__23307),
            .I(N__23303));
    InMux I__2945 (
            .O(N__23306),
            .I(N__23300));
    Odrv12 I__2944 (
            .O(N__23303),
            .I(IAC_SCLK));
    LocalMux I__2943 (
            .O(N__23300),
            .I(IAC_SCLK));
    InMux I__2942 (
            .O(N__23295),
            .I(bfn_8_17_0_));
    InMux I__2941 (
            .O(N__23292),
            .I(\ADC_IAC.n19649 ));
    InMux I__2940 (
            .O(N__23289),
            .I(\ADC_IAC.n19650 ));
    InMux I__2939 (
            .O(N__23286),
            .I(\ADC_IAC.n19651 ));
    InMux I__2938 (
            .O(N__23283),
            .I(\ADC_IAC.n19652 ));
    InMux I__2937 (
            .O(N__23280),
            .I(\ADC_IAC.n19653 ));
    CascadeMux I__2936 (
            .O(N__23277),
            .I(N__23273));
    InMux I__2935 (
            .O(N__23276),
            .I(N__23270));
    InMux I__2934 (
            .O(N__23273),
            .I(N__23267));
    LocalMux I__2933 (
            .O(N__23270),
            .I(buf_readRTD_8));
    LocalMux I__2932 (
            .O(N__23267),
            .I(buf_readRTD_8));
    CascadeMux I__2931 (
            .O(N__23262),
            .I(N__23258));
    InMux I__2930 (
            .O(N__23261),
            .I(N__23254));
    InMux I__2929 (
            .O(N__23258),
            .I(N__23251));
    CascadeMux I__2928 (
            .O(N__23257),
            .I(N__23248));
    LocalMux I__2927 (
            .O(N__23254),
            .I(N__23245));
    LocalMux I__2926 (
            .O(N__23251),
            .I(N__23242));
    InMux I__2925 (
            .O(N__23248),
            .I(N__23239));
    Span4Mux_h I__2924 (
            .O(N__23245),
            .I(N__23236));
    Span4Mux_v I__2923 (
            .O(N__23242),
            .I(N__23233));
    LocalMux I__2922 (
            .O(N__23239),
            .I(N__23230));
    Span4Mux_v I__2921 (
            .O(N__23236),
            .I(N__23227));
    Span4Mux_v I__2920 (
            .O(N__23233),
            .I(N__23224));
    Span4Mux_h I__2919 (
            .O(N__23230),
            .I(N__23221));
    Span4Mux_v I__2918 (
            .O(N__23227),
            .I(N__23216));
    Span4Mux_h I__2917 (
            .O(N__23224),
            .I(N__23213));
    Span4Mux_v I__2916 (
            .O(N__23221),
            .I(N__23210));
    InMux I__2915 (
            .O(N__23220),
            .I(N__23205));
    InMux I__2914 (
            .O(N__23219),
            .I(N__23205));
    Odrv4 I__2913 (
            .O(N__23216),
            .I(buf_cfgRTD_0));
    Odrv4 I__2912 (
            .O(N__23213),
            .I(buf_cfgRTD_0));
    Odrv4 I__2911 (
            .O(N__23210),
            .I(buf_cfgRTD_0));
    LocalMux I__2910 (
            .O(N__23205),
            .I(buf_cfgRTD_0));
    CascadeMux I__2909 (
            .O(N__23196),
            .I(N__23193));
    InMux I__2908 (
            .O(N__23193),
            .I(N__23190));
    LocalMux I__2907 (
            .O(N__23190),
            .I(n21202));
    IoInMux I__2906 (
            .O(N__23187),
            .I(N__23184));
    LocalMux I__2905 (
            .O(N__23184),
            .I(N__23181));
    Span4Mux_s0_h I__2904 (
            .O(N__23181),
            .I(N__23178));
    Sp12to4 I__2903 (
            .O(N__23178),
            .I(N__23175));
    Span12Mux_s11_v I__2902 (
            .O(N__23175),
            .I(N__23170));
    InMux I__2901 (
            .O(N__23174),
            .I(N__23167));
    InMux I__2900 (
            .O(N__23173),
            .I(N__23164));
    Odrv12 I__2899 (
            .O(N__23170),
            .I(VAC_OSR1));
    LocalMux I__2898 (
            .O(N__23167),
            .I(VAC_OSR1));
    LocalMux I__2897 (
            .O(N__23164),
            .I(VAC_OSR1));
    InMux I__2896 (
            .O(N__23157),
            .I(N__23153));
    InMux I__2895 (
            .O(N__23156),
            .I(N__23150));
    LocalMux I__2894 (
            .O(N__23153),
            .I(N__23147));
    LocalMux I__2893 (
            .O(N__23150),
            .I(N__23144));
    Span4Mux_h I__2892 (
            .O(N__23147),
            .I(N__23140));
    Span4Mux_v I__2891 (
            .O(N__23144),
            .I(N__23137));
    InMux I__2890 (
            .O(N__23143),
            .I(N__23134));
    Odrv4 I__2889 (
            .O(N__23140),
            .I(cmd_rdadctmp_16));
    Odrv4 I__2888 (
            .O(N__23137),
            .I(cmd_rdadctmp_16));
    LocalMux I__2887 (
            .O(N__23134),
            .I(cmd_rdadctmp_16));
    CascadeMux I__2886 (
            .O(N__23127),
            .I(N__23124));
    InMux I__2885 (
            .O(N__23124),
            .I(N__23117));
    InMux I__2884 (
            .O(N__23123),
            .I(N__23117));
    CascadeMux I__2883 (
            .O(N__23122),
            .I(N__23114));
    LocalMux I__2882 (
            .O(N__23117),
            .I(N__23111));
    InMux I__2881 (
            .O(N__23114),
            .I(N__23108));
    Odrv4 I__2880 (
            .O(N__23111),
            .I(cmd_rdadctmp_17));
    LocalMux I__2879 (
            .O(N__23108),
            .I(cmd_rdadctmp_17));
    CascadeMux I__2878 (
            .O(N__23103),
            .I(N__23096));
    InMux I__2877 (
            .O(N__23102),
            .I(N__23093));
    InMux I__2876 (
            .O(N__23101),
            .I(N__23090));
    InMux I__2875 (
            .O(N__23100),
            .I(N__23087));
    InMux I__2874 (
            .O(N__23099),
            .I(N__23084));
    InMux I__2873 (
            .O(N__23096),
            .I(N__23081));
    LocalMux I__2872 (
            .O(N__23093),
            .I(N__23072));
    LocalMux I__2871 (
            .O(N__23090),
            .I(N__23072));
    LocalMux I__2870 (
            .O(N__23087),
            .I(N__23072));
    LocalMux I__2869 (
            .O(N__23084),
            .I(N__23072));
    LocalMux I__2868 (
            .O(N__23081),
            .I(N__23069));
    Span4Mux_v I__2867 (
            .O(N__23072),
            .I(N__23066));
    Span12Mux_v I__2866 (
            .O(N__23069),
            .I(N__23061));
    Sp12to4 I__2865 (
            .O(N__23066),
            .I(N__23061));
    Odrv12 I__2864 (
            .O(N__23061),
            .I(VAC_DRDY));
    IoInMux I__2863 (
            .O(N__23058),
            .I(N__23055));
    LocalMux I__2862 (
            .O(N__23055),
            .I(N__23052));
    Span12Mux_s8_h I__2861 (
            .O(N__23052),
            .I(N__23048));
    InMux I__2860 (
            .O(N__23051),
            .I(N__23044));
    Span12Mux_v I__2859 (
            .O(N__23048),
            .I(N__23041));
    InMux I__2858 (
            .O(N__23047),
            .I(N__23038));
    LocalMux I__2857 (
            .O(N__23044),
            .I(N__23035));
    Odrv12 I__2856 (
            .O(N__23041),
            .I(AMPV_POW));
    LocalMux I__2855 (
            .O(N__23038),
            .I(AMPV_POW));
    Odrv4 I__2854 (
            .O(N__23035),
            .I(AMPV_POW));
    CascadeMux I__2853 (
            .O(N__23028),
            .I(n23_adj_1540_cascade_));
    InMux I__2852 (
            .O(N__23025),
            .I(N__23022));
    LocalMux I__2851 (
            .O(N__23022),
            .I(n21123));
    InMux I__2850 (
            .O(N__23019),
            .I(N__23016));
    LocalMux I__2849 (
            .O(N__23016),
            .I(N__23013));
    Span4Mux_v I__2848 (
            .O(N__23013),
            .I(N__23010));
    Sp12to4 I__2847 (
            .O(N__23010),
            .I(N__23007));
    Span12Mux_h I__2846 (
            .O(N__23007),
            .I(N__23004));
    Span12Mux_v I__2845 (
            .O(N__23004),
            .I(N__23001));
    Odrv12 I__2844 (
            .O(N__23001),
            .I(EIS_SYNCCLK));
    IoInMux I__2843 (
            .O(N__22998),
            .I(N__22995));
    LocalMux I__2842 (
            .O(N__22995),
            .I(N__22991));
    IoInMux I__2841 (
            .O(N__22994),
            .I(N__22988));
    IoSpan4Mux I__2840 (
            .O(N__22991),
            .I(N__22985));
    LocalMux I__2839 (
            .O(N__22988),
            .I(N__22982));
    Span4Mux_s2_h I__2838 (
            .O(N__22985),
            .I(N__22979));
    IoSpan4Mux I__2837 (
            .O(N__22982),
            .I(N__22976));
    Span4Mux_h I__2836 (
            .O(N__22979),
            .I(N__22973));
    Span4Mux_s2_v I__2835 (
            .O(N__22976),
            .I(N__22970));
    Span4Mux_h I__2834 (
            .O(N__22973),
            .I(N__22967));
    Sp12to4 I__2833 (
            .O(N__22970),
            .I(N__22964));
    Span4Mux_v I__2832 (
            .O(N__22967),
            .I(N__22961));
    Odrv12 I__2831 (
            .O(N__22964),
            .I(IAC_CLK));
    Odrv4 I__2830 (
            .O(N__22961),
            .I(IAC_CLK));
    CascadeMux I__2829 (
            .O(N__22956),
            .I(N__22953));
    InMux I__2828 (
            .O(N__22953),
            .I(N__22950));
    LocalMux I__2827 (
            .O(N__22950),
            .I(N__22947));
    Span4Mux_h I__2826 (
            .O(N__22947),
            .I(N__22942));
    InMux I__2825 (
            .O(N__22946),
            .I(N__22937));
    InMux I__2824 (
            .O(N__22945),
            .I(N__22937));
    Odrv4 I__2823 (
            .O(N__22942),
            .I(cmd_rdadctmp_15));
    LocalMux I__2822 (
            .O(N__22937),
            .I(cmd_rdadctmp_15));
    InMux I__2821 (
            .O(N__22932),
            .I(N__22929));
    LocalMux I__2820 (
            .O(N__22929),
            .I(N__22926));
    Span4Mux_h I__2819 (
            .O(N__22926),
            .I(N__22923));
    Odrv4 I__2818 (
            .O(N__22923),
            .I(n21082));
    InMux I__2817 (
            .O(N__22920),
            .I(N__22917));
    LocalMux I__2816 (
            .O(N__22917),
            .I(N__22914));
    Odrv12 I__2815 (
            .O(N__22914),
            .I(n21201));
    CascadeMux I__2814 (
            .O(N__22911),
            .I(n22315_cascade_));
    InMux I__2813 (
            .O(N__22908),
            .I(N__22905));
    LocalMux I__2812 (
            .O(N__22905),
            .I(n22318));
    CascadeMux I__2811 (
            .O(N__22902),
            .I(N__22899));
    InMux I__2810 (
            .O(N__22899),
            .I(N__22896));
    LocalMux I__2809 (
            .O(N__22896),
            .I(N__22892));
    CascadeMux I__2808 (
            .O(N__22895),
            .I(N__22888));
    Span4Mux_h I__2807 (
            .O(N__22892),
            .I(N__22885));
    InMux I__2806 (
            .O(N__22891),
            .I(N__22880));
    InMux I__2805 (
            .O(N__22888),
            .I(N__22880));
    Odrv4 I__2804 (
            .O(N__22885),
            .I(cmd_rdadctmp_22));
    LocalMux I__2803 (
            .O(N__22880),
            .I(cmd_rdadctmp_22));
    CascadeMux I__2802 (
            .O(N__22875),
            .I(N__22871));
    CascadeMux I__2801 (
            .O(N__22874),
            .I(N__22868));
    InMux I__2800 (
            .O(N__22871),
            .I(N__22865));
    InMux I__2799 (
            .O(N__22868),
            .I(N__22862));
    LocalMux I__2798 (
            .O(N__22865),
            .I(cmd_rdadctmp_31_adj_1419));
    LocalMux I__2797 (
            .O(N__22862),
            .I(cmd_rdadctmp_31_adj_1419));
    CascadeMux I__2796 (
            .O(N__22857),
            .I(N__22852));
    InMux I__2795 (
            .O(N__22856),
            .I(N__22847));
    InMux I__2794 (
            .O(N__22855),
            .I(N__22847));
    InMux I__2793 (
            .O(N__22852),
            .I(N__22844));
    LocalMux I__2792 (
            .O(N__22847),
            .I(cmd_rdadctmp_30_adj_1420));
    LocalMux I__2791 (
            .O(N__22844),
            .I(cmd_rdadctmp_30_adj_1420));
    InMux I__2790 (
            .O(N__22839),
            .I(N__22836));
    LocalMux I__2789 (
            .O(N__22836),
            .I(N__22833));
    Odrv4 I__2788 (
            .O(N__22833),
            .I(n22405));
    InMux I__2787 (
            .O(N__22830),
            .I(N__22827));
    LocalMux I__2786 (
            .O(N__22827),
            .I(N__22824));
    Span4Mux_v I__2785 (
            .O(N__22824),
            .I(N__22821));
    Span4Mux_v I__2784 (
            .O(N__22821),
            .I(N__22817));
    CascadeMux I__2783 (
            .O(N__22820),
            .I(N__22814));
    Span4Mux_h I__2782 (
            .O(N__22817),
            .I(N__22811));
    InMux I__2781 (
            .O(N__22814),
            .I(N__22807));
    Span4Mux_h I__2780 (
            .O(N__22811),
            .I(N__22804));
    InMux I__2779 (
            .O(N__22810),
            .I(N__22801));
    LocalMux I__2778 (
            .O(N__22807),
            .I(N__22798));
    Span4Mux_h I__2777 (
            .O(N__22804),
            .I(N__22795));
    LocalMux I__2776 (
            .O(N__22801),
            .I(buf_adcdata_vac_21));
    Odrv4 I__2775 (
            .O(N__22798),
            .I(buf_adcdata_vac_21));
    Odrv4 I__2774 (
            .O(N__22795),
            .I(buf_adcdata_vac_21));
    InMux I__2773 (
            .O(N__22788),
            .I(N__22785));
    LocalMux I__2772 (
            .O(N__22785),
            .I(n21097));
    InMux I__2771 (
            .O(N__22782),
            .I(N__22778));
    CascadeMux I__2770 (
            .O(N__22781),
            .I(N__22774));
    LocalMux I__2769 (
            .O(N__22778),
            .I(N__22771));
    InMux I__2768 (
            .O(N__22777),
            .I(N__22768));
    InMux I__2767 (
            .O(N__22774),
            .I(N__22765));
    Sp12to4 I__2766 (
            .O(N__22771),
            .I(N__22760));
    LocalMux I__2765 (
            .O(N__22768),
            .I(N__22760));
    LocalMux I__2764 (
            .O(N__22765),
            .I(N__22757));
    Span12Mux_v I__2763 (
            .O(N__22760),
            .I(N__22752));
    Span4Mux_h I__2762 (
            .O(N__22757),
            .I(N__22749));
    InMux I__2761 (
            .O(N__22756),
            .I(N__22744));
    InMux I__2760 (
            .O(N__22755),
            .I(N__22744));
    Odrv12 I__2759 (
            .O(N__22752),
            .I(buf_cfgRTD_4));
    Odrv4 I__2758 (
            .O(N__22749),
            .I(buf_cfgRTD_4));
    LocalMux I__2757 (
            .O(N__22744),
            .I(buf_cfgRTD_4));
    CascadeMux I__2756 (
            .O(N__22737),
            .I(N__22734));
    InMux I__2755 (
            .O(N__22734),
            .I(N__22731));
    LocalMux I__2754 (
            .O(N__22731),
            .I(N__22728));
    Span4Mux_h I__2753 (
            .O(N__22728),
            .I(N__22724));
    CascadeMux I__2752 (
            .O(N__22727),
            .I(N__22721));
    Span4Mux_v I__2751 (
            .O(N__22724),
            .I(N__22718));
    InMux I__2750 (
            .O(N__22721),
            .I(N__22715));
    Odrv4 I__2749 (
            .O(N__22718),
            .I(buf_readRTD_12));
    LocalMux I__2748 (
            .O(N__22715),
            .I(buf_readRTD_12));
    CascadeMux I__2747 (
            .O(N__22710),
            .I(N__22707));
    InMux I__2746 (
            .O(N__22707),
            .I(N__22704));
    LocalMux I__2745 (
            .O(N__22704),
            .I(N__22701));
    Span4Mux_v I__2744 (
            .O(N__22701),
            .I(N__22697));
    CascadeMux I__2743 (
            .O(N__22700),
            .I(N__22694));
    Span4Mux_v I__2742 (
            .O(N__22697),
            .I(N__22691));
    InMux I__2741 (
            .O(N__22694),
            .I(N__22688));
    Odrv4 I__2740 (
            .O(N__22691),
            .I(buf_readRTD_4));
    LocalMux I__2739 (
            .O(N__22688),
            .I(buf_readRTD_4));
    InMux I__2738 (
            .O(N__22683),
            .I(N__22680));
    LocalMux I__2737 (
            .O(N__22680),
            .I(N__22676));
    InMux I__2736 (
            .O(N__22679),
            .I(N__22672));
    Span12Mux_h I__2735 (
            .O(N__22676),
            .I(N__22669));
    InMux I__2734 (
            .O(N__22675),
            .I(N__22666));
    LocalMux I__2733 (
            .O(N__22672),
            .I(buf_adcdata_vac_16));
    Odrv12 I__2732 (
            .O(N__22669),
            .I(buf_adcdata_vac_16));
    LocalMux I__2731 (
            .O(N__22666),
            .I(buf_adcdata_vac_16));
    InMux I__2730 (
            .O(N__22659),
            .I(N__22656));
    LocalMux I__2729 (
            .O(N__22656),
            .I(N__22652));
    CascadeMux I__2728 (
            .O(N__22655),
            .I(N__22649));
    Span4Mux_v I__2727 (
            .O(N__22652),
            .I(N__22646));
    InMux I__2726 (
            .O(N__22649),
            .I(N__22643));
    Odrv4 I__2725 (
            .O(N__22646),
            .I(cmd_rdadctmp_3));
    LocalMux I__2724 (
            .O(N__22643),
            .I(cmd_rdadctmp_3));
    InMux I__2723 (
            .O(N__22638),
            .I(N__22633));
    CascadeMux I__2722 (
            .O(N__22637),
            .I(N__22630));
    InMux I__2721 (
            .O(N__22636),
            .I(N__22627));
    LocalMux I__2720 (
            .O(N__22633),
            .I(N__22624));
    InMux I__2719 (
            .O(N__22630),
            .I(N__22621));
    LocalMux I__2718 (
            .O(N__22627),
            .I(cmd_rdadctmp_27_adj_1423));
    Odrv12 I__2717 (
            .O(N__22624),
            .I(cmd_rdadctmp_27_adj_1423));
    LocalMux I__2716 (
            .O(N__22621),
            .I(cmd_rdadctmp_27_adj_1423));
    CascadeMux I__2715 (
            .O(N__22614),
            .I(N__22609));
    InMux I__2714 (
            .O(N__22613),
            .I(N__22606));
    InMux I__2713 (
            .O(N__22612),
            .I(N__22601));
    InMux I__2712 (
            .O(N__22609),
            .I(N__22601));
    LocalMux I__2711 (
            .O(N__22606),
            .I(cmd_rdadctmp_28_adj_1422));
    LocalMux I__2710 (
            .O(N__22601),
            .I(cmd_rdadctmp_28_adj_1422));
    InMux I__2709 (
            .O(N__22596),
            .I(N__22592));
    CascadeMux I__2708 (
            .O(N__22595),
            .I(N__22589));
    LocalMux I__2707 (
            .O(N__22592),
            .I(N__22586));
    InMux I__2706 (
            .O(N__22589),
            .I(N__22582));
    Span4Mux_v I__2705 (
            .O(N__22586),
            .I(N__22579));
    InMux I__2704 (
            .O(N__22585),
            .I(N__22576));
    LocalMux I__2703 (
            .O(N__22582),
            .I(cmd_rdadctmp_29_adj_1421));
    Odrv4 I__2702 (
            .O(N__22579),
            .I(cmd_rdadctmp_29_adj_1421));
    LocalMux I__2701 (
            .O(N__22576),
            .I(cmd_rdadctmp_29_adj_1421));
    CascadeMux I__2700 (
            .O(N__22569),
            .I(N__22566));
    InMux I__2699 (
            .O(N__22566),
            .I(N__22563));
    LocalMux I__2698 (
            .O(N__22563),
            .I(N__22559));
    CascadeMux I__2697 (
            .O(N__22562),
            .I(N__22556));
    Span4Mux_h I__2696 (
            .O(N__22559),
            .I(N__22553));
    InMux I__2695 (
            .O(N__22556),
            .I(N__22550));
    Odrv4 I__2694 (
            .O(N__22553),
            .I(cmd_rdadctmp_7_adj_1443));
    LocalMux I__2693 (
            .O(N__22550),
            .I(cmd_rdadctmp_7_adj_1443));
    InMux I__2692 (
            .O(N__22545),
            .I(\ADC_VDC.n19688 ));
    InMux I__2691 (
            .O(N__22542),
            .I(\ADC_VDC.n19689 ));
    InMux I__2690 (
            .O(N__22539),
            .I(\ADC_VDC.n19690 ));
    InMux I__2689 (
            .O(N__22536),
            .I(\ADC_VDC.n19691 ));
    InMux I__2688 (
            .O(N__22533),
            .I(\ADC_VDC.n19692 ));
    InMux I__2687 (
            .O(N__22530),
            .I(\ADC_VDC.n19693 ));
    InMux I__2686 (
            .O(N__22527),
            .I(bfn_8_10_0_));
    InMux I__2685 (
            .O(N__22524),
            .I(\ADC_VDC.n19695 ));
    CEMux I__2684 (
            .O(N__22521),
            .I(N__22516));
    CEMux I__2683 (
            .O(N__22520),
            .I(N__22510));
    CEMux I__2682 (
            .O(N__22519),
            .I(N__22507));
    LocalMux I__2681 (
            .O(N__22516),
            .I(N__22503));
    CEMux I__2680 (
            .O(N__22515),
            .I(N__22500));
    CEMux I__2679 (
            .O(N__22514),
            .I(N__22497));
    CEMux I__2678 (
            .O(N__22513),
            .I(N__22494));
    LocalMux I__2677 (
            .O(N__22510),
            .I(N__22489));
    LocalMux I__2676 (
            .O(N__22507),
            .I(N__22489));
    CEMux I__2675 (
            .O(N__22506),
            .I(N__22486));
    Span4Mux_h I__2674 (
            .O(N__22503),
            .I(N__22483));
    LocalMux I__2673 (
            .O(N__22500),
            .I(N__22480));
    LocalMux I__2672 (
            .O(N__22497),
            .I(N__22477));
    LocalMux I__2671 (
            .O(N__22494),
            .I(N__22474));
    Span4Mux_v I__2670 (
            .O(N__22489),
            .I(N__22467));
    LocalMux I__2669 (
            .O(N__22486),
            .I(N__22467));
    Span4Mux_h I__2668 (
            .O(N__22483),
            .I(N__22467));
    Span4Mux_v I__2667 (
            .O(N__22480),
            .I(N__22462));
    Span4Mux_v I__2666 (
            .O(N__22477),
            .I(N__22462));
    Odrv4 I__2665 (
            .O(N__22474),
            .I(\ADC_VDC.n13010 ));
    Odrv4 I__2664 (
            .O(N__22467),
            .I(\ADC_VDC.n13010 ));
    Odrv4 I__2663 (
            .O(N__22462),
            .I(\ADC_VDC.n13010 ));
    SRMux I__2662 (
            .O(N__22455),
            .I(N__22448));
    SRMux I__2661 (
            .O(N__22454),
            .I(N__22444));
    SRMux I__2660 (
            .O(N__22453),
            .I(N__22440));
    SRMux I__2659 (
            .O(N__22452),
            .I(N__22437));
    SRMux I__2658 (
            .O(N__22451),
            .I(N__22434));
    LocalMux I__2657 (
            .O(N__22448),
            .I(N__22431));
    SRMux I__2656 (
            .O(N__22447),
            .I(N__22428));
    LocalMux I__2655 (
            .O(N__22444),
            .I(N__22425));
    SRMux I__2654 (
            .O(N__22443),
            .I(N__22422));
    LocalMux I__2653 (
            .O(N__22440),
            .I(N__22419));
    LocalMux I__2652 (
            .O(N__22437),
            .I(N__22416));
    LocalMux I__2651 (
            .O(N__22434),
            .I(N__22413));
    Span4Mux_v I__2650 (
            .O(N__22431),
            .I(N__22408));
    LocalMux I__2649 (
            .O(N__22428),
            .I(N__22408));
    Span4Mux_v I__2648 (
            .O(N__22425),
            .I(N__22401));
    LocalMux I__2647 (
            .O(N__22422),
            .I(N__22401));
    Span4Mux_h I__2646 (
            .O(N__22419),
            .I(N__22401));
    Span4Mux_h I__2645 (
            .O(N__22416),
            .I(N__22398));
    Odrv12 I__2644 (
            .O(N__22413),
            .I(\ADC_VDC.n14915 ));
    Odrv4 I__2643 (
            .O(N__22408),
            .I(\ADC_VDC.n14915 ));
    Odrv4 I__2642 (
            .O(N__22401),
            .I(\ADC_VDC.n14915 ));
    Odrv4 I__2641 (
            .O(N__22398),
            .I(\ADC_VDC.n14915 ));
    InMux I__2640 (
            .O(N__22389),
            .I(\ADC_VDC.n19696 ));
    InMux I__2639 (
            .O(N__22386),
            .I(N__22383));
    LocalMux I__2638 (
            .O(N__22383),
            .I(N__22380));
    Odrv12 I__2637 (
            .O(N__22380),
            .I(\ADC_VDC.cmd_rdadcbuf_35_N_1138_34 ));
    CascadeMux I__2636 (
            .O(N__22377),
            .I(N__22372));
    InMux I__2635 (
            .O(N__22376),
            .I(N__22367));
    InMux I__2634 (
            .O(N__22375),
            .I(N__22367));
    InMux I__2633 (
            .O(N__22372),
            .I(N__22364));
    LocalMux I__2632 (
            .O(N__22367),
            .I(cmd_rdadctmp_17_adj_1462));
    LocalMux I__2631 (
            .O(N__22364),
            .I(cmd_rdadctmp_17_adj_1462));
    InMux I__2630 (
            .O(N__22359),
            .I(\ADC_VDC.n19679 ));
    InMux I__2629 (
            .O(N__22356),
            .I(\ADC_VDC.n19680 ));
    InMux I__2628 (
            .O(N__22353),
            .I(\ADC_VDC.n19681 ));
    CascadeMux I__2627 (
            .O(N__22350),
            .I(N__22346));
    CascadeMux I__2626 (
            .O(N__22349),
            .I(N__22342));
    InMux I__2625 (
            .O(N__22346),
            .I(N__22339));
    InMux I__2624 (
            .O(N__22345),
            .I(N__22336));
    InMux I__2623 (
            .O(N__22342),
            .I(N__22333));
    LocalMux I__2622 (
            .O(N__22339),
            .I(cmd_rdadctmp_20_adj_1459));
    LocalMux I__2621 (
            .O(N__22336),
            .I(cmd_rdadctmp_20_adj_1459));
    LocalMux I__2620 (
            .O(N__22333),
            .I(cmd_rdadctmp_20_adj_1459));
    InMux I__2619 (
            .O(N__22326),
            .I(\ADC_VDC.n19682 ));
    CascadeMux I__2618 (
            .O(N__22323),
            .I(N__22318));
    InMux I__2617 (
            .O(N__22322),
            .I(N__22313));
    InMux I__2616 (
            .O(N__22321),
            .I(N__22313));
    InMux I__2615 (
            .O(N__22318),
            .I(N__22310));
    LocalMux I__2614 (
            .O(N__22313),
            .I(cmd_rdadctmp_21_adj_1458));
    LocalMux I__2613 (
            .O(N__22310),
            .I(cmd_rdadctmp_21_adj_1458));
    InMux I__2612 (
            .O(N__22305),
            .I(\ADC_VDC.n19683 ));
    InMux I__2611 (
            .O(N__22302),
            .I(\ADC_VDC.n19684 ));
    InMux I__2610 (
            .O(N__22299),
            .I(\ADC_VDC.n19685 ));
    InMux I__2609 (
            .O(N__22296),
            .I(bfn_8_9_0_));
    InMux I__2608 (
            .O(N__22293),
            .I(\ADC_VDC.n19687 ));
    InMux I__2607 (
            .O(N__22290),
            .I(N__22287));
    LocalMux I__2606 (
            .O(N__22287),
            .I(\ADC_VDC.cmd_rdadcbuf_9 ));
    InMux I__2605 (
            .O(N__22284),
            .I(\ADC_VDC.n19671 ));
    InMux I__2604 (
            .O(N__22281),
            .I(N__22278));
    LocalMux I__2603 (
            .O(N__22278),
            .I(\ADC_VDC.cmd_rdadcbuf_10 ));
    InMux I__2602 (
            .O(N__22275),
            .I(\ADC_VDC.n19672 ));
    CascadeMux I__2601 (
            .O(N__22272),
            .I(N__22268));
    CascadeMux I__2600 (
            .O(N__22271),
            .I(N__22264));
    InMux I__2599 (
            .O(N__22268),
            .I(N__22259));
    InMux I__2598 (
            .O(N__22267),
            .I(N__22259));
    InMux I__2597 (
            .O(N__22264),
            .I(N__22256));
    LocalMux I__2596 (
            .O(N__22259),
            .I(cmd_rdadctmp_11_adj_1468));
    LocalMux I__2595 (
            .O(N__22256),
            .I(cmd_rdadctmp_11_adj_1468));
    InMux I__2594 (
            .O(N__22251),
            .I(\ADC_VDC.n19673 ));
    InMux I__2593 (
            .O(N__22248),
            .I(\ADC_VDC.n19674 ));
    InMux I__2592 (
            .O(N__22245),
            .I(\ADC_VDC.n19675 ));
    InMux I__2591 (
            .O(N__22242),
            .I(\ADC_VDC.n19676 ));
    InMux I__2590 (
            .O(N__22239),
            .I(\ADC_VDC.n19677 ));
    InMux I__2589 (
            .O(N__22236),
            .I(N__22233));
    LocalMux I__2588 (
            .O(N__22233),
            .I(N__22229));
    InMux I__2587 (
            .O(N__22232),
            .I(N__22226));
    Odrv4 I__2586 (
            .O(N__22229),
            .I(cmd_rdadcbuf_16));
    LocalMux I__2585 (
            .O(N__22226),
            .I(cmd_rdadcbuf_16));
    InMux I__2584 (
            .O(N__22221),
            .I(bfn_8_8_0_));
    InMux I__2583 (
            .O(N__22218),
            .I(N__22215));
    LocalMux I__2582 (
            .O(N__22215),
            .I(\ADC_VDC.cmd_rdadcbuf_0 ));
    CascadeMux I__2581 (
            .O(N__22212),
            .I(N__22207));
    InMux I__2580 (
            .O(N__22211),
            .I(N__22202));
    InMux I__2579 (
            .O(N__22210),
            .I(N__22202));
    InMux I__2578 (
            .O(N__22207),
            .I(N__22199));
    LocalMux I__2577 (
            .O(N__22202),
            .I(cmd_rdadctmp_1_adj_1478));
    LocalMux I__2576 (
            .O(N__22199),
            .I(cmd_rdadctmp_1_adj_1478));
    InMux I__2575 (
            .O(N__22194),
            .I(N__22191));
    LocalMux I__2574 (
            .O(N__22191),
            .I(\ADC_VDC.cmd_rdadcbuf_1 ));
    InMux I__2573 (
            .O(N__22188),
            .I(\ADC_VDC.n19663 ));
    CascadeMux I__2572 (
            .O(N__22185),
            .I(N__22180));
    InMux I__2571 (
            .O(N__22184),
            .I(N__22175));
    InMux I__2570 (
            .O(N__22183),
            .I(N__22175));
    InMux I__2569 (
            .O(N__22180),
            .I(N__22172));
    LocalMux I__2568 (
            .O(N__22175),
            .I(cmd_rdadctmp_2_adj_1477));
    LocalMux I__2567 (
            .O(N__22172),
            .I(cmd_rdadctmp_2_adj_1477));
    InMux I__2566 (
            .O(N__22167),
            .I(N__22164));
    LocalMux I__2565 (
            .O(N__22164),
            .I(\ADC_VDC.cmd_rdadcbuf_2 ));
    InMux I__2564 (
            .O(N__22161),
            .I(\ADC_VDC.n19664 ));
    InMux I__2563 (
            .O(N__22158),
            .I(N__22155));
    LocalMux I__2562 (
            .O(N__22155),
            .I(\ADC_VDC.cmd_rdadcbuf_3 ));
    InMux I__2561 (
            .O(N__22152),
            .I(\ADC_VDC.n19665 ));
    InMux I__2560 (
            .O(N__22149),
            .I(N__22146));
    LocalMux I__2559 (
            .O(N__22146),
            .I(\ADC_VDC.cmd_rdadcbuf_4 ));
    InMux I__2558 (
            .O(N__22143),
            .I(\ADC_VDC.n19666 ));
    InMux I__2557 (
            .O(N__22140),
            .I(N__22137));
    LocalMux I__2556 (
            .O(N__22137),
            .I(\ADC_VDC.cmd_rdadcbuf_5 ));
    InMux I__2555 (
            .O(N__22134),
            .I(\ADC_VDC.n19667 ));
    InMux I__2554 (
            .O(N__22131),
            .I(N__22128));
    LocalMux I__2553 (
            .O(N__22128),
            .I(\ADC_VDC.cmd_rdadcbuf_6 ));
    InMux I__2552 (
            .O(N__22125),
            .I(\ADC_VDC.n19668 ));
    CascadeMux I__2551 (
            .O(N__22122),
            .I(N__22119));
    InMux I__2550 (
            .O(N__22119),
            .I(N__22116));
    LocalMux I__2549 (
            .O(N__22116),
            .I(\ADC_VDC.cmd_rdadcbuf_7 ));
    InMux I__2548 (
            .O(N__22113),
            .I(\ADC_VDC.n19669 ));
    InMux I__2547 (
            .O(N__22110),
            .I(N__22107));
    LocalMux I__2546 (
            .O(N__22107),
            .I(\ADC_VDC.cmd_rdadcbuf_8 ));
    InMux I__2545 (
            .O(N__22104),
            .I(bfn_8_7_0_));
    InMux I__2544 (
            .O(N__22101),
            .I(N__22097));
    InMux I__2543 (
            .O(N__22100),
            .I(N__22094));
    LocalMux I__2542 (
            .O(N__22097),
            .I(N__22091));
    LocalMux I__2541 (
            .O(N__22094),
            .I(\ADC_VDC.avg_cnt_10 ));
    Odrv4 I__2540 (
            .O(N__22091),
            .I(\ADC_VDC.avg_cnt_10 ));
    InMux I__2539 (
            .O(N__22086),
            .I(\ADC_VDC.n19707 ));
    InMux I__2538 (
            .O(N__22083),
            .I(\ADC_VDC.n19708 ));
    CascadeMux I__2537 (
            .O(N__22080),
            .I(\ADC_VDC.n13010_cascade_ ));
    CascadeMux I__2536 (
            .O(N__22077),
            .I(n12871_cascade_));
    CascadeMux I__2535 (
            .O(N__22074),
            .I(N__22069));
    InMux I__2534 (
            .O(N__22073),
            .I(N__22064));
    InMux I__2533 (
            .O(N__22072),
            .I(N__22064));
    InMux I__2532 (
            .O(N__22069),
            .I(N__22061));
    LocalMux I__2531 (
            .O(N__22064),
            .I(cmd_rdadctmp_0_adj_1479));
    LocalMux I__2530 (
            .O(N__22061),
            .I(cmd_rdadctmp_0_adj_1479));
    InMux I__2529 (
            .O(N__22056),
            .I(\ADC_VDC.n19698 ));
    InMux I__2528 (
            .O(N__22053),
            .I(\ADC_VDC.n19699 ));
    InMux I__2527 (
            .O(N__22050),
            .I(\ADC_VDC.n19700 ));
    InMux I__2526 (
            .O(N__22047),
            .I(\ADC_VDC.n19701 ));
    InMux I__2525 (
            .O(N__22044),
            .I(\ADC_VDC.n19702 ));
    InMux I__2524 (
            .O(N__22041),
            .I(\ADC_VDC.n19703 ));
    InMux I__2523 (
            .O(N__22038),
            .I(\ADC_VDC.n19704 ));
    CascadeMux I__2522 (
            .O(N__22035),
            .I(N__22032));
    InMux I__2521 (
            .O(N__22032),
            .I(N__22028));
    InMux I__2520 (
            .O(N__22031),
            .I(N__22025));
    LocalMux I__2519 (
            .O(N__22028),
            .I(N__22022));
    LocalMux I__2518 (
            .O(N__22025),
            .I(\ADC_VDC.avg_cnt_8 ));
    Odrv4 I__2517 (
            .O(N__22022),
            .I(\ADC_VDC.avg_cnt_8 ));
    InMux I__2516 (
            .O(N__22017),
            .I(bfn_8_4_0_));
    InMux I__2515 (
            .O(N__22014),
            .I(N__22010));
    InMux I__2514 (
            .O(N__22013),
            .I(N__22007));
    LocalMux I__2513 (
            .O(N__22010),
            .I(N__22004));
    LocalMux I__2512 (
            .O(N__22007),
            .I(\ADC_VDC.avg_cnt_9 ));
    Odrv4 I__2511 (
            .O(N__22004),
            .I(\ADC_VDC.avg_cnt_9 ));
    InMux I__2510 (
            .O(N__21999),
            .I(\ADC_VDC.n19706 ));
    CascadeMux I__2509 (
            .O(N__21996),
            .I(\ADC_VDC.n19_cascade_ ));
    CascadeMux I__2508 (
            .O(N__21993),
            .I(\ADC_VDC.n18563_cascade_ ));
    InMux I__2507 (
            .O(N__21990),
            .I(N__21987));
    LocalMux I__2506 (
            .O(N__21987),
            .I(\ADC_VDC.n18563 ));
    CascadeMux I__2505 (
            .O(N__21984),
            .I(\ADC_VDC.n21384_cascade_ ));
    CEMux I__2504 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__2503 (
            .O(N__21978),
            .I(N__21975));
    Odrv4 I__2502 (
            .O(N__21975),
            .I(\ADC_VDC.n13034 ));
    InMux I__2501 (
            .O(N__21972),
            .I(N__21968));
    InMux I__2500 (
            .O(N__21971),
            .I(N__21965));
    LocalMux I__2499 (
            .O(N__21968),
            .I(\ADC_VDC.avg_cnt_0 ));
    LocalMux I__2498 (
            .O(N__21965),
            .I(\ADC_VDC.avg_cnt_0 ));
    InMux I__2497 (
            .O(N__21960),
            .I(bfn_8_3_0_));
    IoInMux I__2496 (
            .O(N__21957),
            .I(N__21954));
    LocalMux I__2495 (
            .O(N__21954),
            .I(N__21951));
    IoSpan4Mux I__2494 (
            .O(N__21951),
            .I(N__21948));
    Span4Mux_s3_h I__2493 (
            .O(N__21948),
            .I(N__21944));
    CascadeMux I__2492 (
            .O(N__21947),
            .I(N__21941));
    Span4Mux_h I__2491 (
            .O(N__21944),
            .I(N__21938));
    InMux I__2490 (
            .O(N__21941),
            .I(N__21935));
    Odrv4 I__2489 (
            .O(N__21938),
            .I(VAC_SCLK));
    LocalMux I__2488 (
            .O(N__21935),
            .I(VAC_SCLK));
    InMux I__2487 (
            .O(N__21930),
            .I(N__21927));
    LocalMux I__2486 (
            .O(N__21927),
            .I(N__21923));
    InMux I__2485 (
            .O(N__21926),
            .I(N__21920));
    Odrv4 I__2484 (
            .O(N__21923),
            .I(cmd_rdadctmp_5_adj_1445));
    LocalMux I__2483 (
            .O(N__21920),
            .I(cmd_rdadctmp_5_adj_1445));
    CascadeMux I__2482 (
            .O(N__21915),
            .I(N__21911));
    InMux I__2481 (
            .O(N__21914),
            .I(N__21906));
    InMux I__2480 (
            .O(N__21911),
            .I(N__21906));
    LocalMux I__2479 (
            .O(N__21906),
            .I(cmd_rdadctmp_6_adj_1444));
    InMux I__2478 (
            .O(N__21903),
            .I(N__21900));
    LocalMux I__2477 (
            .O(N__21900),
            .I(\ADC_VAC.n21312 ));
    CascadeMux I__2476 (
            .O(N__21897),
            .I(\ADC_VAC.n20958_cascade_ ));
    CEMux I__2475 (
            .O(N__21894),
            .I(N__21891));
    LocalMux I__2474 (
            .O(N__21891),
            .I(N__21888));
    Span4Mux_h I__2473 (
            .O(N__21888),
            .I(N__21885));
    Odrv4 I__2472 (
            .O(N__21885),
            .I(\ADC_VAC.n20959 ));
    InMux I__2471 (
            .O(N__21882),
            .I(N__21878));
    CascadeMux I__2470 (
            .O(N__21881),
            .I(N__21874));
    LocalMux I__2469 (
            .O(N__21878),
            .I(N__21871));
    CascadeMux I__2468 (
            .O(N__21877),
            .I(N__21868));
    InMux I__2467 (
            .O(N__21874),
            .I(N__21865));
    Span4Mux_v I__2466 (
            .O(N__21871),
            .I(N__21862));
    InMux I__2465 (
            .O(N__21868),
            .I(N__21859));
    LocalMux I__2464 (
            .O(N__21865),
            .I(N__21856));
    Span4Mux_h I__2463 (
            .O(N__21862),
            .I(N__21851));
    LocalMux I__2462 (
            .O(N__21859),
            .I(N__21851));
    Span4Mux_v I__2461 (
            .O(N__21856),
            .I(N__21848));
    Span4Mux_v I__2460 (
            .O(N__21851),
            .I(N__21845));
    Span4Mux_h I__2459 (
            .O(N__21848),
            .I(N__21840));
    Sp12to4 I__2458 (
            .O(N__21845),
            .I(N__21837));
    InMux I__2457 (
            .O(N__21844),
            .I(N__21834));
    InMux I__2456 (
            .O(N__21843),
            .I(N__21831));
    Odrv4 I__2455 (
            .O(N__21840),
            .I(buf_cfgRTD_2));
    Odrv12 I__2454 (
            .O(N__21837),
            .I(buf_cfgRTD_2));
    LocalMux I__2453 (
            .O(N__21834),
            .I(buf_cfgRTD_2));
    LocalMux I__2452 (
            .O(N__21831),
            .I(buf_cfgRTD_2));
    CascadeMux I__2451 (
            .O(N__21822),
            .I(N__21818));
    InMux I__2450 (
            .O(N__21821),
            .I(N__21815));
    InMux I__2449 (
            .O(N__21818),
            .I(N__21812));
    LocalMux I__2448 (
            .O(N__21815),
            .I(N__21808));
    LocalMux I__2447 (
            .O(N__21812),
            .I(N__21805));
    CascadeMux I__2446 (
            .O(N__21811),
            .I(N__21802));
    Span4Mux_v I__2445 (
            .O(N__21808),
            .I(N__21797));
    Span4Mux_v I__2444 (
            .O(N__21805),
            .I(N__21797));
    InMux I__2443 (
            .O(N__21802),
            .I(N__21794));
    Span4Mux_v I__2442 (
            .O(N__21797),
            .I(N__21790));
    LocalMux I__2441 (
            .O(N__21794),
            .I(N__21786));
    InMux I__2440 (
            .O(N__21793),
            .I(N__21783));
    Span4Mux_h I__2439 (
            .O(N__21790),
            .I(N__21780));
    InMux I__2438 (
            .O(N__21789),
            .I(N__21777));
    Span4Mux_v I__2437 (
            .O(N__21786),
            .I(N__21772));
    LocalMux I__2436 (
            .O(N__21783),
            .I(N__21772));
    Odrv4 I__2435 (
            .O(N__21780),
            .I(buf_cfgRTD_5));
    LocalMux I__2434 (
            .O(N__21777),
            .I(buf_cfgRTD_5));
    Odrv4 I__2433 (
            .O(N__21772),
            .I(buf_cfgRTD_5));
    InMux I__2432 (
            .O(N__21765),
            .I(N__21760));
    CascadeMux I__2431 (
            .O(N__21764),
            .I(N__21757));
    CascadeMux I__2430 (
            .O(N__21763),
            .I(N__21754));
    LocalMux I__2429 (
            .O(N__21760),
            .I(N__21751));
    InMux I__2428 (
            .O(N__21757),
            .I(N__21746));
    InMux I__2427 (
            .O(N__21754),
            .I(N__21746));
    Odrv4 I__2426 (
            .O(N__21751),
            .I(cmd_rdadctmp_24_adj_1426));
    LocalMux I__2425 (
            .O(N__21746),
            .I(cmd_rdadctmp_24_adj_1426));
    CascadeMux I__2424 (
            .O(N__21741),
            .I(n22321_cascade_));
    InMux I__2423 (
            .O(N__21738),
            .I(N__21735));
    LocalMux I__2422 (
            .O(N__21735),
            .I(N__21730));
    InMux I__2421 (
            .O(N__21734),
            .I(N__21725));
    InMux I__2420 (
            .O(N__21733),
            .I(N__21725));
    Odrv4 I__2419 (
            .O(N__21730),
            .I(read_buf_8));
    LocalMux I__2418 (
            .O(N__21725),
            .I(read_buf_8));
    InMux I__2417 (
            .O(N__21720),
            .I(N__21713));
    InMux I__2416 (
            .O(N__21719),
            .I(N__21713));
    InMux I__2415 (
            .O(N__21718),
            .I(N__21705));
    LocalMux I__2414 (
            .O(N__21713),
            .I(N__21698));
    InMux I__2413 (
            .O(N__21712),
            .I(N__21693));
    InMux I__2412 (
            .O(N__21711),
            .I(N__21693));
    InMux I__2411 (
            .O(N__21710),
            .I(N__21688));
    InMux I__2410 (
            .O(N__21709),
            .I(N__21688));
    InMux I__2409 (
            .O(N__21708),
            .I(N__21685));
    LocalMux I__2408 (
            .O(N__21705),
            .I(N__21680));
    InMux I__2407 (
            .O(N__21704),
            .I(N__21671));
    InMux I__2406 (
            .O(N__21703),
            .I(N__21671));
    InMux I__2405 (
            .O(N__21702),
            .I(N__21671));
    InMux I__2404 (
            .O(N__21701),
            .I(N__21671));
    Span4Mux_v I__2403 (
            .O(N__21698),
            .I(N__21663));
    LocalMux I__2402 (
            .O(N__21693),
            .I(N__21663));
    LocalMux I__2401 (
            .O(N__21688),
            .I(N__21663));
    LocalMux I__2400 (
            .O(N__21685),
            .I(N__21660));
    InMux I__2399 (
            .O(N__21684),
            .I(N__21655));
    InMux I__2398 (
            .O(N__21683),
            .I(N__21655));
    Span4Mux_v I__2397 (
            .O(N__21680),
            .I(N__21650));
    LocalMux I__2396 (
            .O(N__21671),
            .I(N__21650));
    InMux I__2395 (
            .O(N__21670),
            .I(N__21647));
    Span4Mux_v I__2394 (
            .O(N__21663),
            .I(N__21640));
    Span4Mux_h I__2393 (
            .O(N__21660),
            .I(N__21640));
    LocalMux I__2392 (
            .O(N__21655),
            .I(N__21640));
    Span4Mux_h I__2391 (
            .O(N__21650),
            .I(N__21634));
    LocalMux I__2390 (
            .O(N__21647),
            .I(N__21634));
    Span4Mux_h I__2389 (
            .O(N__21640),
            .I(N__21631));
    InMux I__2388 (
            .O(N__21639),
            .I(N__21628));
    Span4Mux_v I__2387 (
            .O(N__21634),
            .I(N__21625));
    Span4Mux_h I__2386 (
            .O(N__21631),
            .I(N__21622));
    LocalMux I__2385 (
            .O(N__21628),
            .I(N__21619));
    Odrv4 I__2384 (
            .O(N__21625),
            .I(n11714));
    Odrv4 I__2383 (
            .O(N__21622),
            .I(n11714));
    Odrv12 I__2382 (
            .O(N__21619),
            .I(n11714));
    CascadeMux I__2381 (
            .O(N__21612),
            .I(N__21608));
    CascadeMux I__2380 (
            .O(N__21611),
            .I(N__21605));
    InMux I__2379 (
            .O(N__21608),
            .I(N__21602));
    InMux I__2378 (
            .O(N__21605),
            .I(N__21599));
    LocalMux I__2377 (
            .O(N__21602),
            .I(N__21596));
    LocalMux I__2376 (
            .O(N__21599),
            .I(N__21593));
    Span4Mux_v I__2375 (
            .O(N__21596),
            .I(N__21589));
    Span4Mux_h I__2374 (
            .O(N__21593),
            .I(N__21586));
    InMux I__2373 (
            .O(N__21592),
            .I(N__21583));
    Odrv4 I__2372 (
            .O(N__21589),
            .I(cmd_rdadctmp_13_adj_1437));
    Odrv4 I__2371 (
            .O(N__21586),
            .I(cmd_rdadctmp_13_adj_1437));
    LocalMux I__2370 (
            .O(N__21583),
            .I(cmd_rdadctmp_13_adj_1437));
    InMux I__2369 (
            .O(N__21576),
            .I(N__21573));
    LocalMux I__2368 (
            .O(N__21573),
            .I(N__21570));
    Span12Mux_s11_h I__2367 (
            .O(N__21570),
            .I(N__21565));
    InMux I__2366 (
            .O(N__21569),
            .I(N__21562));
    InMux I__2365 (
            .O(N__21568),
            .I(N__21559));
    Span12Mux_v I__2364 (
            .O(N__21565),
            .I(N__21556));
    LocalMux I__2363 (
            .O(N__21562),
            .I(N__21553));
    LocalMux I__2362 (
            .O(N__21559),
            .I(buf_adcdata_vac_8));
    Odrv12 I__2361 (
            .O(N__21556),
            .I(buf_adcdata_vac_8));
    Odrv4 I__2360 (
            .O(N__21553),
            .I(buf_adcdata_vac_8));
    InMux I__2359 (
            .O(N__21546),
            .I(N__21543));
    LocalMux I__2358 (
            .O(N__21543),
            .I(N__21539));
    CascadeMux I__2357 (
            .O(N__21542),
            .I(N__21535));
    Span4Mux_h I__2356 (
            .O(N__21539),
            .I(N__21532));
    InMux I__2355 (
            .O(N__21538),
            .I(N__21529));
    InMux I__2354 (
            .O(N__21535),
            .I(N__21526));
    Span4Mux_v I__2353 (
            .O(N__21532),
            .I(N__21523));
    LocalMux I__2352 (
            .O(N__21529),
            .I(N__21520));
    LocalMux I__2351 (
            .O(N__21526),
            .I(buf_adcdata_vac_6));
    Odrv4 I__2350 (
            .O(N__21523),
            .I(buf_adcdata_vac_6));
    Odrv12 I__2349 (
            .O(N__21520),
            .I(buf_adcdata_vac_6));
    CascadeMux I__2348 (
            .O(N__21513),
            .I(N__21509));
    InMux I__2347 (
            .O(N__21512),
            .I(N__21501));
    InMux I__2346 (
            .O(N__21509),
            .I(N__21501));
    InMux I__2345 (
            .O(N__21508),
            .I(N__21501));
    LocalMux I__2344 (
            .O(N__21501),
            .I(cmd_rdadctmp_14_adj_1436));
    CascadeMux I__2343 (
            .O(N__21498),
            .I(N__21495));
    InMux I__2342 (
            .O(N__21495),
            .I(N__21489));
    InMux I__2341 (
            .O(N__21494),
            .I(N__21489));
    LocalMux I__2340 (
            .O(N__21489),
            .I(N__21486));
    Span4Mux_h I__2339 (
            .O(N__21486),
            .I(N__21482));
    InMux I__2338 (
            .O(N__21485),
            .I(N__21479));
    Odrv4 I__2337 (
            .O(N__21482),
            .I(cmd_rdadctmp_15_adj_1435));
    LocalMux I__2336 (
            .O(N__21479),
            .I(cmd_rdadctmp_15_adj_1435));
    CascadeMux I__2335 (
            .O(N__21474),
            .I(N__21470));
    CascadeMux I__2334 (
            .O(N__21473),
            .I(N__21466));
    InMux I__2333 (
            .O(N__21470),
            .I(N__21459));
    InMux I__2332 (
            .O(N__21469),
            .I(N__21459));
    InMux I__2331 (
            .O(N__21466),
            .I(N__21459));
    LocalMux I__2330 (
            .O(N__21459),
            .I(cmd_rdadctmp_16_adj_1434));
    InMux I__2329 (
            .O(N__21456),
            .I(N__21453));
    LocalMux I__2328 (
            .O(N__21453),
            .I(N__21450));
    Odrv4 I__2327 (
            .O(N__21450),
            .I(buf_data_iac_4));
    InMux I__2326 (
            .O(N__21447),
            .I(N__21444));
    LocalMux I__2325 (
            .O(N__21444),
            .I(n22_adj_1633));
    InMux I__2324 (
            .O(N__21441),
            .I(N__21437));
    InMux I__2323 (
            .O(N__21440),
            .I(N__21434));
    LocalMux I__2322 (
            .O(N__21437),
            .I(bit_cnt_3));
    LocalMux I__2321 (
            .O(N__21434),
            .I(bit_cnt_3));
    InMux I__2320 (
            .O(N__21429),
            .I(N__21426));
    LocalMux I__2319 (
            .O(N__21426),
            .I(n21456));
    CascadeMux I__2318 (
            .O(N__21423),
            .I(N__21417));
    InMux I__2317 (
            .O(N__21422),
            .I(N__21410));
    InMux I__2316 (
            .O(N__21421),
            .I(N__21410));
    InMux I__2315 (
            .O(N__21420),
            .I(N__21410));
    InMux I__2314 (
            .O(N__21417),
            .I(N__21407));
    LocalMux I__2313 (
            .O(N__21410),
            .I(bit_cnt_1));
    LocalMux I__2312 (
            .O(N__21407),
            .I(bit_cnt_1));
    CascadeMux I__2311 (
            .O(N__21402),
            .I(N__21399));
    InMux I__2310 (
            .O(N__21399),
            .I(N__21392));
    InMux I__2309 (
            .O(N__21398),
            .I(N__21392));
    InMux I__2308 (
            .O(N__21397),
            .I(N__21389));
    LocalMux I__2307 (
            .O(N__21392),
            .I(bit_cnt_2));
    LocalMux I__2306 (
            .O(N__21389),
            .I(bit_cnt_2));
    InMux I__2305 (
            .O(N__21384),
            .I(N__21381));
    LocalMux I__2304 (
            .O(N__21381),
            .I(n8_adj_1602));
    CEMux I__2303 (
            .O(N__21378),
            .I(N__21374));
    CEMux I__2302 (
            .O(N__21377),
            .I(N__21371));
    LocalMux I__2301 (
            .O(N__21374),
            .I(N__21368));
    LocalMux I__2300 (
            .O(N__21371),
            .I(N__21365));
    Span4Mux_v I__2299 (
            .O(N__21368),
            .I(N__21362));
    Odrv12 I__2298 (
            .O(N__21365),
            .I(\CLK_DDS.n9 ));
    Odrv4 I__2297 (
            .O(N__21362),
            .I(\CLK_DDS.n9 ));
    InMux I__2296 (
            .O(N__21357),
            .I(N__21354));
    LocalMux I__2295 (
            .O(N__21354),
            .I(n19_adj_1626));
    InMux I__2294 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__2293 (
            .O(N__21348),
            .I(n20867));
    CascadeMux I__2292 (
            .O(N__21345),
            .I(n20867_cascade_));
    InMux I__2291 (
            .O(N__21342),
            .I(N__21339));
    LocalMux I__2290 (
            .O(N__21339),
            .I(N__21336));
    Span4Mux_v I__2289 (
            .O(N__21336),
            .I(N__21333));
    Span4Mux_v I__2288 (
            .O(N__21333),
            .I(N__21330));
    IoSpan4Mux I__2287 (
            .O(N__21330),
            .I(N__21327));
    Odrv4 I__2286 (
            .O(N__21327),
            .I(IAC_MISO));
    CascadeMux I__2285 (
            .O(N__21324),
            .I(n12498_cascade_));
    InMux I__2284 (
            .O(N__21321),
            .I(N__21315));
    InMux I__2283 (
            .O(N__21320),
            .I(N__21315));
    LocalMux I__2282 (
            .O(N__21315),
            .I(cmd_rdadctmp_0));
    CascadeMux I__2281 (
            .O(N__21312),
            .I(N__21308));
    InMux I__2280 (
            .O(N__21311),
            .I(N__21303));
    InMux I__2279 (
            .O(N__21308),
            .I(N__21303));
    LocalMux I__2278 (
            .O(N__21303),
            .I(cmd_rdadctmp_1));
    CascadeMux I__2277 (
            .O(N__21300),
            .I(N__21296));
    InMux I__2276 (
            .O(N__21299),
            .I(N__21293));
    InMux I__2275 (
            .O(N__21296),
            .I(N__21290));
    LocalMux I__2274 (
            .O(N__21293),
            .I(N__21287));
    LocalMux I__2273 (
            .O(N__21290),
            .I(cmd_rdadctmp_2));
    Odrv12 I__2272 (
            .O(N__21287),
            .I(cmd_rdadctmp_2));
    IoInMux I__2271 (
            .O(N__21282),
            .I(N__21279));
    LocalMux I__2270 (
            .O(N__21279),
            .I(N__21276));
    Span4Mux_s3_v I__2269 (
            .O(N__21276),
            .I(N__21273));
    Span4Mux_h I__2268 (
            .O(N__21273),
            .I(N__21270));
    Span4Mux_v I__2267 (
            .O(N__21270),
            .I(N__21267));
    Odrv4 I__2266 (
            .O(N__21267),
            .I(AC_ADC_SYNC));
    InMux I__2265 (
            .O(N__21264),
            .I(N__21260));
    CascadeMux I__2264 (
            .O(N__21263),
            .I(N__21257));
    LocalMux I__2263 (
            .O(N__21260),
            .I(N__21254));
    InMux I__2262 (
            .O(N__21257),
            .I(N__21251));
    Odrv4 I__2261 (
            .O(N__21254),
            .I(buf_adcdata_vdc_5));
    LocalMux I__2260 (
            .O(N__21251),
            .I(buf_adcdata_vdc_5));
    CascadeMux I__2259 (
            .O(N__21246),
            .I(N__21242));
    CascadeMux I__2258 (
            .O(N__21245),
            .I(N__21239));
    InMux I__2257 (
            .O(N__21242),
            .I(N__21234));
    InMux I__2256 (
            .O(N__21239),
            .I(N__21234));
    LocalMux I__2255 (
            .O(N__21234),
            .I(cmd_rdadctmp_4_adj_1446));
    InMux I__2254 (
            .O(N__21231),
            .I(N__21228));
    LocalMux I__2253 (
            .O(N__21228),
            .I(n20864));
    CascadeMux I__2252 (
            .O(N__21225),
            .I(n20864_cascade_));
    CascadeMux I__2251 (
            .O(N__21222),
            .I(\ADC_VAC.n17_cascade_ ));
    CEMux I__2250 (
            .O(N__21219),
            .I(N__21216));
    LocalMux I__2249 (
            .O(N__21216),
            .I(\ADC_VAC.n12 ));
    IoInMux I__2248 (
            .O(N__21213),
            .I(N__21210));
    LocalMux I__2247 (
            .O(N__21210),
            .I(N__21207));
    IoSpan4Mux I__2246 (
            .O(N__21207),
            .I(N__21204));
    Span4Mux_s2_v I__2245 (
            .O(N__21204),
            .I(N__21200));
    CascadeMux I__2244 (
            .O(N__21203),
            .I(N__21197));
    Span4Mux_v I__2243 (
            .O(N__21200),
            .I(N__21194));
    InMux I__2242 (
            .O(N__21197),
            .I(N__21191));
    Odrv4 I__2241 (
            .O(N__21194),
            .I(IAC_CS));
    LocalMux I__2240 (
            .O(N__21191),
            .I(IAC_CS));
    InMux I__2239 (
            .O(N__21186),
            .I(N__21183));
    LocalMux I__2238 (
            .O(N__21183),
            .I(n14_adj_1612));
    InMux I__2237 (
            .O(N__21180),
            .I(N__21175));
    InMux I__2236 (
            .O(N__21179),
            .I(N__21172));
    CascadeMux I__2235 (
            .O(N__21178),
            .I(N__21169));
    LocalMux I__2234 (
            .O(N__21175),
            .I(N__21166));
    LocalMux I__2233 (
            .O(N__21172),
            .I(N__21163));
    InMux I__2232 (
            .O(N__21169),
            .I(N__21160));
    Span4Mux_v I__2231 (
            .O(N__21166),
            .I(N__21157));
    Span4Mux_h I__2230 (
            .O(N__21163),
            .I(N__21152));
    LocalMux I__2229 (
            .O(N__21160),
            .I(N__21152));
    Span4Mux_v I__2228 (
            .O(N__21157),
            .I(N__21147));
    Span4Mux_v I__2227 (
            .O(N__21152),
            .I(N__21144));
    InMux I__2226 (
            .O(N__21151),
            .I(N__21141));
    InMux I__2225 (
            .O(N__21150),
            .I(N__21138));
    Odrv4 I__2224 (
            .O(N__21147),
            .I(buf_cfgRTD_1));
    Odrv4 I__2223 (
            .O(N__21144),
            .I(buf_cfgRTD_1));
    LocalMux I__2222 (
            .O(N__21141),
            .I(buf_cfgRTD_1));
    LocalMux I__2221 (
            .O(N__21138),
            .I(buf_cfgRTD_1));
    CascadeMux I__2220 (
            .O(N__21129),
            .I(n14_adj_1610_cascade_));
    IoInMux I__2219 (
            .O(N__21126),
            .I(N__21123));
    LocalMux I__2218 (
            .O(N__21123),
            .I(N__21120));
    Span4Mux_s2_h I__2217 (
            .O(N__21120),
            .I(N__21117));
    Span4Mux_h I__2216 (
            .O(N__21117),
            .I(N__21113));
    CascadeMux I__2215 (
            .O(N__21116),
            .I(N__21110));
    Span4Mux_v I__2214 (
            .O(N__21113),
            .I(N__21107));
    InMux I__2213 (
            .O(N__21110),
            .I(N__21104));
    Odrv4 I__2212 (
            .O(N__21107),
            .I(VAC_CS));
    LocalMux I__2211 (
            .O(N__21104),
            .I(VAC_CS));
    CascadeMux I__2210 (
            .O(N__21099),
            .I(N__21096));
    InMux I__2209 (
            .O(N__21096),
            .I(N__21092));
    CascadeMux I__2208 (
            .O(N__21095),
            .I(N__21089));
    LocalMux I__2207 (
            .O(N__21092),
            .I(N__21086));
    InMux I__2206 (
            .O(N__21089),
            .I(N__21082));
    Sp12to4 I__2205 (
            .O(N__21086),
            .I(N__21079));
    InMux I__2204 (
            .O(N__21085),
            .I(N__21076));
    LocalMux I__2203 (
            .O(N__21082),
            .I(cmd_rdadctmp_14));
    Odrv12 I__2202 (
            .O(N__21079),
            .I(cmd_rdadctmp_14));
    LocalMux I__2201 (
            .O(N__21076),
            .I(cmd_rdadctmp_14));
    InMux I__2200 (
            .O(N__21069),
            .I(N__21065));
    CascadeMux I__2199 (
            .O(N__21068),
            .I(N__21062));
    LocalMux I__2198 (
            .O(N__21065),
            .I(N__21059));
    InMux I__2197 (
            .O(N__21062),
            .I(N__21056));
    Odrv4 I__2196 (
            .O(N__21059),
            .I(cmd_rdadctmp_2_adj_1448));
    LocalMux I__2195 (
            .O(N__21056),
            .I(cmd_rdadctmp_2_adj_1448));
    CascadeMux I__2194 (
            .O(N__21051),
            .I(N__21047));
    InMux I__2193 (
            .O(N__21050),
            .I(N__21042));
    InMux I__2192 (
            .O(N__21047),
            .I(N__21042));
    LocalMux I__2191 (
            .O(N__21042),
            .I(cmd_rdadctmp_3_adj_1447));
    InMux I__2190 (
            .O(N__21039),
            .I(N__21036));
    LocalMux I__2189 (
            .O(N__21036),
            .I(N__21033));
    Span4Mux_v I__2188 (
            .O(N__21033),
            .I(N__21028));
    InMux I__2187 (
            .O(N__21032),
            .I(N__21025));
    InMux I__2186 (
            .O(N__21031),
            .I(N__21022));
    Odrv4 I__2185 (
            .O(N__21028),
            .I(read_buf_7));
    LocalMux I__2184 (
            .O(N__21025),
            .I(read_buf_7));
    LocalMux I__2183 (
            .O(N__21022),
            .I(read_buf_7));
    InMux I__2182 (
            .O(N__21015),
            .I(N__21012));
    LocalMux I__2181 (
            .O(N__21012),
            .I(N__21008));
    CascadeMux I__2180 (
            .O(N__21011),
            .I(N__21005));
    Span4Mux_v I__2179 (
            .O(N__21008),
            .I(N__21002));
    InMux I__2178 (
            .O(N__21005),
            .I(N__20999));
    Odrv4 I__2177 (
            .O(N__21002),
            .I(buf_readRTD_10));
    LocalMux I__2176 (
            .O(N__20999),
            .I(buf_readRTD_10));
    InMux I__2175 (
            .O(N__20994),
            .I(N__20980));
    InMux I__2174 (
            .O(N__20993),
            .I(N__20975));
    InMux I__2173 (
            .O(N__20992),
            .I(N__20975));
    InMux I__2172 (
            .O(N__20991),
            .I(N__20968));
    InMux I__2171 (
            .O(N__20990),
            .I(N__20968));
    InMux I__2170 (
            .O(N__20989),
            .I(N__20968));
    InMux I__2169 (
            .O(N__20988),
            .I(N__20961));
    InMux I__2168 (
            .O(N__20987),
            .I(N__20961));
    InMux I__2167 (
            .O(N__20986),
            .I(N__20961));
    InMux I__2166 (
            .O(N__20985),
            .I(N__20958));
    InMux I__2165 (
            .O(N__20984),
            .I(N__20953));
    InMux I__2164 (
            .O(N__20983),
            .I(N__20953));
    LocalMux I__2163 (
            .O(N__20980),
            .I(N__20941));
    LocalMux I__2162 (
            .O(N__20975),
            .I(N__20941));
    LocalMux I__2161 (
            .O(N__20968),
            .I(N__20941));
    LocalMux I__2160 (
            .O(N__20961),
            .I(N__20941));
    LocalMux I__2159 (
            .O(N__20958),
            .I(N__20936));
    LocalMux I__2158 (
            .O(N__20953),
            .I(N__20936));
    InMux I__2157 (
            .O(N__20952),
            .I(N__20931));
    InMux I__2156 (
            .O(N__20951),
            .I(N__20931));
    InMux I__2155 (
            .O(N__20950),
            .I(N__20928));
    Span4Mux_v I__2154 (
            .O(N__20941),
            .I(N__20925));
    Span4Mux_h I__2153 (
            .O(N__20936),
            .I(N__20922));
    LocalMux I__2152 (
            .O(N__20931),
            .I(n1_adj_1606));
    LocalMux I__2151 (
            .O(N__20928),
            .I(n1_adj_1606));
    Odrv4 I__2150 (
            .O(N__20925),
            .I(n1_adj_1606));
    Odrv4 I__2149 (
            .O(N__20922),
            .I(n1_adj_1606));
    CascadeMux I__2148 (
            .O(N__20913),
            .I(N__20908));
    CascadeMux I__2147 (
            .O(N__20912),
            .I(N__20905));
    CascadeMux I__2146 (
            .O(N__20911),
            .I(N__20900));
    InMux I__2145 (
            .O(N__20908),
            .I(N__20888));
    InMux I__2144 (
            .O(N__20905),
            .I(N__20888));
    InMux I__2143 (
            .O(N__20904),
            .I(N__20883));
    InMux I__2142 (
            .O(N__20903),
            .I(N__20883));
    InMux I__2141 (
            .O(N__20900),
            .I(N__20880));
    InMux I__2140 (
            .O(N__20899),
            .I(N__20871));
    InMux I__2139 (
            .O(N__20898),
            .I(N__20871));
    InMux I__2138 (
            .O(N__20897),
            .I(N__20871));
    InMux I__2137 (
            .O(N__20896),
            .I(N__20871));
    InMux I__2136 (
            .O(N__20895),
            .I(N__20864));
    InMux I__2135 (
            .O(N__20894),
            .I(N__20864));
    InMux I__2134 (
            .O(N__20893),
            .I(N__20864));
    LocalMux I__2133 (
            .O(N__20888),
            .I(N__20855));
    LocalMux I__2132 (
            .O(N__20883),
            .I(N__20855));
    LocalMux I__2131 (
            .O(N__20880),
            .I(N__20852));
    LocalMux I__2130 (
            .O(N__20871),
            .I(N__20847));
    LocalMux I__2129 (
            .O(N__20864),
            .I(N__20847));
    InMux I__2128 (
            .O(N__20863),
            .I(N__20842));
    InMux I__2127 (
            .O(N__20862),
            .I(N__20842));
    InMux I__2126 (
            .O(N__20861),
            .I(N__20837));
    InMux I__2125 (
            .O(N__20860),
            .I(N__20837));
    Span4Mux_h I__2124 (
            .O(N__20855),
            .I(N__20834));
    Span4Mux_v I__2123 (
            .O(N__20852),
            .I(N__20829));
    Span4Mux_v I__2122 (
            .O(N__20847),
            .I(N__20829));
    LocalMux I__2121 (
            .O(N__20842),
            .I(n13293));
    LocalMux I__2120 (
            .O(N__20837),
            .I(n13293));
    Odrv4 I__2119 (
            .O(N__20834),
            .I(n13293));
    Odrv4 I__2118 (
            .O(N__20829),
            .I(n13293));
    InMux I__2117 (
            .O(N__20820),
            .I(N__20817));
    LocalMux I__2116 (
            .O(N__20817),
            .I(N__20812));
    InMux I__2115 (
            .O(N__20816),
            .I(N__20807));
    InMux I__2114 (
            .O(N__20815),
            .I(N__20807));
    Odrv12 I__2113 (
            .O(N__20812),
            .I(read_buf_10));
    LocalMux I__2112 (
            .O(N__20807),
            .I(read_buf_10));
    CascadeMux I__2111 (
            .O(N__20802),
            .I(N__20797));
    InMux I__2110 (
            .O(N__20801),
            .I(N__20794));
    InMux I__2109 (
            .O(N__20800),
            .I(N__20791));
    InMux I__2108 (
            .O(N__20797),
            .I(N__20788));
    LocalMux I__2107 (
            .O(N__20794),
            .I(read_buf_11));
    LocalMux I__2106 (
            .O(N__20791),
            .I(read_buf_11));
    LocalMux I__2105 (
            .O(N__20788),
            .I(read_buf_11));
    CascadeMux I__2104 (
            .O(N__20781),
            .I(N__20776));
    InMux I__2103 (
            .O(N__20780),
            .I(N__20773));
    InMux I__2102 (
            .O(N__20779),
            .I(N__20768));
    InMux I__2101 (
            .O(N__20776),
            .I(N__20768));
    LocalMux I__2100 (
            .O(N__20773),
            .I(read_buf_13));
    LocalMux I__2099 (
            .O(N__20768),
            .I(read_buf_13));
    CascadeMux I__2098 (
            .O(N__20763),
            .I(N__20759));
    CascadeMux I__2097 (
            .O(N__20762),
            .I(N__20756));
    InMux I__2096 (
            .O(N__20759),
            .I(N__20753));
    InMux I__2095 (
            .O(N__20756),
            .I(N__20750));
    LocalMux I__2094 (
            .O(N__20753),
            .I(buf_readRTD_13));
    LocalMux I__2093 (
            .O(N__20750),
            .I(buf_readRTD_13));
    CascadeMux I__2092 (
            .O(N__20745),
            .I(N__20741));
    CascadeMux I__2091 (
            .O(N__20744),
            .I(N__20737));
    InMux I__2090 (
            .O(N__20741),
            .I(N__20734));
    InMux I__2089 (
            .O(N__20740),
            .I(N__20729));
    InMux I__2088 (
            .O(N__20737),
            .I(N__20729));
    LocalMux I__2087 (
            .O(N__20734),
            .I(read_buf_9));
    LocalMux I__2086 (
            .O(N__20729),
            .I(read_buf_9));
    CascadeMux I__2085 (
            .O(N__20724),
            .I(N__20721));
    InMux I__2084 (
            .O(N__20721),
            .I(N__20717));
    InMux I__2083 (
            .O(N__20720),
            .I(N__20714));
    LocalMux I__2082 (
            .O(N__20717),
            .I(buf_readRTD_9));
    LocalMux I__2081 (
            .O(N__20714),
            .I(buf_readRTD_9));
    CascadeMux I__2080 (
            .O(N__20709),
            .I(N__20705));
    CascadeMux I__2079 (
            .O(N__20708),
            .I(N__20702));
    InMux I__2078 (
            .O(N__20705),
            .I(N__20690));
    InMux I__2077 (
            .O(N__20702),
            .I(N__20690));
    InMux I__2076 (
            .O(N__20701),
            .I(N__20690));
    InMux I__2075 (
            .O(N__20700),
            .I(N__20690));
    InMux I__2074 (
            .O(N__20699),
            .I(N__20687));
    LocalMux I__2073 (
            .O(N__20690),
            .I(\RTD.bit_cnt_0 ));
    LocalMux I__2072 (
            .O(N__20687),
            .I(\RTD.bit_cnt_0 ));
    CEMux I__2071 (
            .O(N__20682),
            .I(N__20679));
    LocalMux I__2070 (
            .O(N__20679),
            .I(N__20676));
    Span4Mux_v I__2069 (
            .O(N__20676),
            .I(N__20673));
    Odrv4 I__2068 (
            .O(N__20673),
            .I(\RTD.n11740 ));
    SRMux I__2067 (
            .O(N__20670),
            .I(N__20667));
    LocalMux I__2066 (
            .O(N__20667),
            .I(N__20664));
    Odrv4 I__2065 (
            .O(N__20664),
            .I(\CLK_DDS.n16894 ));
    InMux I__2064 (
            .O(N__20661),
            .I(N__20657));
    InMux I__2063 (
            .O(N__20660),
            .I(N__20654));
    LocalMux I__2062 (
            .O(N__20657),
            .I(read_buf_15));
    LocalMux I__2061 (
            .O(N__20654),
            .I(read_buf_15));
    InMux I__2060 (
            .O(N__20649),
            .I(N__20645));
    InMux I__2059 (
            .O(N__20648),
            .I(N__20641));
    LocalMux I__2058 (
            .O(N__20645),
            .I(N__20638));
    InMux I__2057 (
            .O(N__20644),
            .I(N__20635));
    LocalMux I__2056 (
            .O(N__20641),
            .I(buf_adcdata_iac_6));
    Odrv4 I__2055 (
            .O(N__20638),
            .I(buf_adcdata_iac_6));
    LocalMux I__2054 (
            .O(N__20635),
            .I(buf_adcdata_iac_6));
    InMux I__2053 (
            .O(N__20628),
            .I(N__20625));
    LocalMux I__2052 (
            .O(N__20625),
            .I(n22_adj_1627));
    CascadeMux I__2051 (
            .O(N__20622),
            .I(N__20619));
    InMux I__2050 (
            .O(N__20619),
            .I(N__20610));
    InMux I__2049 (
            .O(N__20618),
            .I(N__20610));
    InMux I__2048 (
            .O(N__20617),
            .I(N__20610));
    LocalMux I__2047 (
            .O(N__20610),
            .I(cmd_rdadctmp_12));
    CascadeMux I__2046 (
            .O(N__20607),
            .I(N__20603));
    CascadeMux I__2045 (
            .O(N__20606),
            .I(N__20600));
    InMux I__2044 (
            .O(N__20603),
            .I(N__20596));
    InMux I__2043 (
            .O(N__20600),
            .I(N__20591));
    InMux I__2042 (
            .O(N__20599),
            .I(N__20591));
    LocalMux I__2041 (
            .O(N__20596),
            .I(cmd_rdadctmp_13));
    LocalMux I__2040 (
            .O(N__20591),
            .I(cmd_rdadctmp_13));
    InMux I__2039 (
            .O(N__20586),
            .I(N__20582));
    InMux I__2038 (
            .O(N__20585),
            .I(N__20579));
    LocalMux I__2037 (
            .O(N__20582),
            .I(N__20575));
    LocalMux I__2036 (
            .O(N__20579),
            .I(N__20571));
    InMux I__2035 (
            .O(N__20578),
            .I(N__20568));
    Span4Mux_h I__2034 (
            .O(N__20575),
            .I(N__20565));
    InMux I__2033 (
            .O(N__20574),
            .I(N__20562));
    Odrv4 I__2032 (
            .O(N__20571),
            .I(\RTD.n17799 ));
    LocalMux I__2031 (
            .O(N__20568),
            .I(\RTD.n17799 ));
    Odrv4 I__2030 (
            .O(N__20565),
            .I(\RTD.n17799 ));
    LocalMux I__2029 (
            .O(N__20562),
            .I(\RTD.n17799 ));
    InMux I__2028 (
            .O(N__20553),
            .I(N__20546));
    InMux I__2027 (
            .O(N__20552),
            .I(N__20546));
    InMux I__2026 (
            .O(N__20551),
            .I(N__20541));
    LocalMux I__2025 (
            .O(N__20546),
            .I(N__20538));
    InMux I__2024 (
            .O(N__20545),
            .I(N__20535));
    InMux I__2023 (
            .O(N__20544),
            .I(N__20532));
    LocalMux I__2022 (
            .O(N__20541),
            .I(N__20529));
    Span4Mux_h I__2021 (
            .O(N__20538),
            .I(N__20524));
    LocalMux I__2020 (
            .O(N__20535),
            .I(N__20524));
    LocalMux I__2019 (
            .O(N__20532),
            .I(\RTD.bit_cnt_3 ));
    Odrv4 I__2018 (
            .O(N__20529),
            .I(\RTD.bit_cnt_3 ));
    Odrv4 I__2017 (
            .O(N__20524),
            .I(\RTD.bit_cnt_3 ));
    InMux I__2016 (
            .O(N__20517),
            .I(N__20507));
    InMux I__2015 (
            .O(N__20516),
            .I(N__20507));
    InMux I__2014 (
            .O(N__20515),
            .I(N__20507));
    InMux I__2013 (
            .O(N__20514),
            .I(N__20504));
    LocalMux I__2012 (
            .O(N__20507),
            .I(\RTD.bit_cnt_1 ));
    LocalMux I__2011 (
            .O(N__20504),
            .I(\RTD.bit_cnt_1 ));
    InMux I__2010 (
            .O(N__20499),
            .I(N__20492));
    InMux I__2009 (
            .O(N__20498),
            .I(N__20492));
    InMux I__2008 (
            .O(N__20497),
            .I(N__20489));
    LocalMux I__2007 (
            .O(N__20492),
            .I(\RTD.bit_cnt_2 ));
    LocalMux I__2006 (
            .O(N__20489),
            .I(\RTD.bit_cnt_2 ));
    InMux I__2005 (
            .O(N__20484),
            .I(N__20481));
    LocalMux I__2004 (
            .O(N__20481),
            .I(N__20478));
    Span4Mux_h I__2003 (
            .O(N__20478),
            .I(N__20473));
    InMux I__2002 (
            .O(N__20477),
            .I(N__20468));
    InMux I__2001 (
            .O(N__20476),
            .I(N__20468));
    Odrv4 I__2000 (
            .O(N__20473),
            .I(buf_adcdata_vac_5));
    LocalMux I__1999 (
            .O(N__20468),
            .I(buf_adcdata_vac_5));
    InMux I__1998 (
            .O(N__20463),
            .I(N__20460));
    LocalMux I__1997 (
            .O(N__20460),
            .I(N__20457));
    Span4Mux_h I__1996 (
            .O(N__20457),
            .I(N__20452));
    InMux I__1995 (
            .O(N__20456),
            .I(N__20447));
    InMux I__1994 (
            .O(N__20455),
            .I(N__20447));
    Odrv4 I__1993 (
            .O(N__20452),
            .I(buf_adcdata_iac_5));
    LocalMux I__1992 (
            .O(N__20447),
            .I(buf_adcdata_iac_5));
    CascadeMux I__1991 (
            .O(N__20442),
            .I(n19_adj_1629_cascade_));
    InMux I__1990 (
            .O(N__20439),
            .I(N__20436));
    LocalMux I__1989 (
            .O(N__20436),
            .I(N__20433));
    Odrv4 I__1988 (
            .O(N__20433),
            .I(buf_data_iac_6));
    InMux I__1987 (
            .O(N__20430),
            .I(N__20426));
    InMux I__1986 (
            .O(N__20429),
            .I(N__20422));
    LocalMux I__1985 (
            .O(N__20426),
            .I(N__20419));
    InMux I__1984 (
            .O(N__20425),
            .I(N__20416));
    LocalMux I__1983 (
            .O(N__20422),
            .I(buf_adcdata_vac_4));
    Odrv4 I__1982 (
            .O(N__20419),
            .I(buf_adcdata_vac_4));
    LocalMux I__1981 (
            .O(N__20416),
            .I(buf_adcdata_vac_4));
    CascadeMux I__1980 (
            .O(N__20409),
            .I(n19_adj_1632_cascade_));
    InMux I__1979 (
            .O(N__20406),
            .I(N__20403));
    LocalMux I__1978 (
            .O(N__20403),
            .I(N__20400));
    Span4Mux_h I__1977 (
            .O(N__20400),
            .I(N__20395));
    InMux I__1976 (
            .O(N__20399),
            .I(N__20390));
    InMux I__1975 (
            .O(N__20398),
            .I(N__20390));
    Odrv4 I__1974 (
            .O(N__20395),
            .I(buf_adcdata_iac_4));
    LocalMux I__1973 (
            .O(N__20390),
            .I(buf_adcdata_iac_4));
    CascadeMux I__1972 (
            .O(N__20385),
            .I(N__20380));
    InMux I__1971 (
            .O(N__20384),
            .I(N__20377));
    InMux I__1970 (
            .O(N__20383),
            .I(N__20372));
    InMux I__1969 (
            .O(N__20380),
            .I(N__20372));
    LocalMux I__1968 (
            .O(N__20377),
            .I(read_buf_12));
    LocalMux I__1967 (
            .O(N__20372),
            .I(read_buf_12));
    CascadeMux I__1966 (
            .O(N__20367),
            .I(N__20363));
    CascadeMux I__1965 (
            .O(N__20366),
            .I(N__20359));
    InMux I__1964 (
            .O(N__20363),
            .I(N__20352));
    InMux I__1963 (
            .O(N__20362),
            .I(N__20352));
    InMux I__1962 (
            .O(N__20359),
            .I(N__20352));
    LocalMux I__1961 (
            .O(N__20352),
            .I(read_buf_14));
    CascadeMux I__1960 (
            .O(N__20349),
            .I(N__20346));
    InMux I__1959 (
            .O(N__20346),
            .I(N__20343));
    LocalMux I__1958 (
            .O(N__20343),
            .I(N__20340));
    Span4Mux_v I__1957 (
            .O(N__20340),
            .I(N__20337));
    Sp12to4 I__1956 (
            .O(N__20337),
            .I(N__20334));
    Odrv12 I__1955 (
            .O(N__20334),
            .I(VAC_MISO));
    InMux I__1954 (
            .O(N__20331),
            .I(N__20328));
    LocalMux I__1953 (
            .O(N__20328),
            .I(N__20324));
    InMux I__1952 (
            .O(N__20327),
            .I(N__20321));
    Odrv4 I__1951 (
            .O(N__20324),
            .I(cmd_rdadctmp_0_adj_1450));
    LocalMux I__1950 (
            .O(N__20321),
            .I(cmd_rdadctmp_0_adj_1450));
    CascadeMux I__1949 (
            .O(N__20316),
            .I(N__20312));
    InMux I__1948 (
            .O(N__20315),
            .I(N__20307));
    InMux I__1947 (
            .O(N__20312),
            .I(N__20307));
    LocalMux I__1946 (
            .O(N__20307),
            .I(cmd_rdadctmp_1_adj_1449));
    IoInMux I__1945 (
            .O(N__20304),
            .I(N__20301));
    LocalMux I__1944 (
            .O(N__20301),
            .I(N__20298));
    IoSpan4Mux I__1943 (
            .O(N__20298),
            .I(N__20295));
    Span4Mux_s3_v I__1942 (
            .O(N__20295),
            .I(N__20292));
    Span4Mux_v I__1941 (
            .O(N__20292),
            .I(N__20289));
    Odrv4 I__1940 (
            .O(N__20289),
            .I(DDS_CS1));
    CEMux I__1939 (
            .O(N__20286),
            .I(N__20283));
    LocalMux I__1938 (
            .O(N__20283),
            .I(N__20280));
    Span4Mux_v I__1937 (
            .O(N__20280),
            .I(N__20277));
    Odrv4 I__1936 (
            .O(N__20277),
            .I(\CLK_DDS.n9_adj_1394 ));
    InMux I__1935 (
            .O(N__20274),
            .I(N__20270));
    InMux I__1934 (
            .O(N__20273),
            .I(N__20267));
    LocalMux I__1933 (
            .O(N__20270),
            .I(N__20262));
    LocalMux I__1932 (
            .O(N__20267),
            .I(N__20262));
    Span4Mux_h I__1931 (
            .O(N__20262),
            .I(N__20258));
    InMux I__1930 (
            .O(N__20261),
            .I(N__20255));
    Odrv4 I__1929 (
            .O(N__20258),
            .I(read_buf_0));
    LocalMux I__1928 (
            .O(N__20255),
            .I(read_buf_0));
    InMux I__1927 (
            .O(N__20250),
            .I(N__20246));
    CascadeMux I__1926 (
            .O(N__20249),
            .I(N__20242));
    LocalMux I__1925 (
            .O(N__20246),
            .I(N__20239));
    InMux I__1924 (
            .O(N__20245),
            .I(N__20234));
    InMux I__1923 (
            .O(N__20242),
            .I(N__20234));
    Odrv4 I__1922 (
            .O(N__20239),
            .I(read_buf_1));
    LocalMux I__1921 (
            .O(N__20234),
            .I(read_buf_1));
    CascadeMux I__1920 (
            .O(N__20229),
            .I(N__20224));
    InMux I__1919 (
            .O(N__20228),
            .I(N__20221));
    InMux I__1918 (
            .O(N__20227),
            .I(N__20218));
    InMux I__1917 (
            .O(N__20224),
            .I(N__20215));
    LocalMux I__1916 (
            .O(N__20221),
            .I(read_buf_5));
    LocalMux I__1915 (
            .O(N__20218),
            .I(read_buf_5));
    LocalMux I__1914 (
            .O(N__20215),
            .I(read_buf_5));
    CascadeMux I__1913 (
            .O(N__20208),
            .I(N__20203));
    InMux I__1912 (
            .O(N__20207),
            .I(N__20200));
    InMux I__1911 (
            .O(N__20206),
            .I(N__20195));
    InMux I__1910 (
            .O(N__20203),
            .I(N__20195));
    LocalMux I__1909 (
            .O(N__20200),
            .I(read_buf_6));
    LocalMux I__1908 (
            .O(N__20195),
            .I(read_buf_6));
    InMux I__1907 (
            .O(N__20190),
            .I(N__20187));
    LocalMux I__1906 (
            .O(N__20187),
            .I(\RTD.cfg_tmp_1 ));
    InMux I__1905 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__1904 (
            .O(N__20181),
            .I(\RTD.cfg_tmp_2 ));
    InMux I__1903 (
            .O(N__20178),
            .I(N__20175));
    LocalMux I__1902 (
            .O(N__20175),
            .I(\RTD.cfg_tmp_3 ));
    InMux I__1901 (
            .O(N__20172),
            .I(N__20169));
    LocalMux I__1900 (
            .O(N__20169),
            .I(\RTD.cfg_tmp_4 ));
    InMux I__1899 (
            .O(N__20166),
            .I(N__20163));
    LocalMux I__1898 (
            .O(N__20163),
            .I(\RTD.cfg_tmp_5 ));
    InMux I__1897 (
            .O(N__20160),
            .I(N__20157));
    LocalMux I__1896 (
            .O(N__20157),
            .I(\RTD.cfg_tmp_6 ));
    CascadeMux I__1895 (
            .O(N__20154),
            .I(N__20151));
    InMux I__1894 (
            .O(N__20151),
            .I(N__20148));
    LocalMux I__1893 (
            .O(N__20148),
            .I(N__20145));
    Span4Mux_v I__1892 (
            .O(N__20145),
            .I(N__20141));
    InMux I__1891 (
            .O(N__20144),
            .I(N__20138));
    Odrv4 I__1890 (
            .O(N__20141),
            .I(\RTD.cfg_tmp_7 ));
    LocalMux I__1889 (
            .O(N__20138),
            .I(\RTD.cfg_tmp_7 ));
    InMux I__1888 (
            .O(N__20133),
            .I(N__20130));
    LocalMux I__1887 (
            .O(N__20130),
            .I(\RTD.cfg_tmp_0 ));
    CEMux I__1886 (
            .O(N__20127),
            .I(N__20124));
    LocalMux I__1885 (
            .O(N__20124),
            .I(N__20121));
    Odrv12 I__1884 (
            .O(N__20121),
            .I(\RTD.n11704 ));
    SRMux I__1883 (
            .O(N__20118),
            .I(N__20115));
    LocalMux I__1882 (
            .O(N__20115),
            .I(N__20112));
    Odrv12 I__1881 (
            .O(N__20112),
            .I(\RTD.n14999 ));
    InMux I__1880 (
            .O(N__20109),
            .I(N__20106));
    LocalMux I__1879 (
            .O(N__20106),
            .I(N__20102));
    InMux I__1878 (
            .O(N__20105),
            .I(N__20099));
    Span4Mux_v I__1877 (
            .O(N__20102),
            .I(N__20096));
    LocalMux I__1876 (
            .O(N__20099),
            .I(N__20093));
    Span4Mux_h I__1875 (
            .O(N__20096),
            .I(N__20089));
    Span4Mux_h I__1874 (
            .O(N__20093),
            .I(N__20086));
    InMux I__1873 (
            .O(N__20092),
            .I(N__20083));
    Odrv4 I__1872 (
            .O(N__20089),
            .I(read_buf_4));
    Odrv4 I__1871 (
            .O(N__20086),
            .I(read_buf_4));
    LocalMux I__1870 (
            .O(N__20083),
            .I(read_buf_4));
    CascadeMux I__1869 (
            .O(N__20076),
            .I(N__20073));
    InMux I__1868 (
            .O(N__20073),
            .I(N__20069));
    CascadeMux I__1867 (
            .O(N__20072),
            .I(N__20065));
    LocalMux I__1866 (
            .O(N__20069),
            .I(N__20062));
    InMux I__1865 (
            .O(N__20068),
            .I(N__20057));
    InMux I__1864 (
            .O(N__20065),
            .I(N__20057));
    Span4Mux_h I__1863 (
            .O(N__20062),
            .I(N__20051));
    LocalMux I__1862 (
            .O(N__20057),
            .I(N__20051));
    InMux I__1861 (
            .O(N__20056),
            .I(N__20048));
    Odrv4 I__1860 (
            .O(N__20051),
            .I(\RTD.mode ));
    LocalMux I__1859 (
            .O(N__20048),
            .I(\RTD.mode ));
    InMux I__1858 (
            .O(N__20043),
            .I(N__20038));
    CascadeMux I__1857 (
            .O(N__20042),
            .I(N__20035));
    CascadeMux I__1856 (
            .O(N__20041),
            .I(N__20032));
    LocalMux I__1855 (
            .O(N__20038),
            .I(N__20029));
    InMux I__1854 (
            .O(N__20035),
            .I(N__20026));
    InMux I__1853 (
            .O(N__20032),
            .I(N__20023));
    Span4Mux_v I__1852 (
            .O(N__20029),
            .I(N__20018));
    LocalMux I__1851 (
            .O(N__20026),
            .I(N__20018));
    LocalMux I__1850 (
            .O(N__20023),
            .I(N__20015));
    Span4Mux_v I__1849 (
            .O(N__20018),
            .I(N__20012));
    Span4Mux_v I__1848 (
            .O(N__20015),
            .I(N__20009));
    Span4Mux_v I__1847 (
            .O(N__20012),
            .I(N__20006));
    Span4Mux_v I__1846 (
            .O(N__20009),
            .I(N__20003));
    Sp12to4 I__1845 (
            .O(N__20006),
            .I(N__19998));
    Sp12to4 I__1844 (
            .O(N__20003),
            .I(N__19998));
    Odrv12 I__1843 (
            .O(N__19998),
            .I(RTD_DRDY));
    InMux I__1842 (
            .O(N__19995),
            .I(N__19992));
    LocalMux I__1841 (
            .O(N__19992),
            .I(N__19986));
    InMux I__1840 (
            .O(N__19991),
            .I(N__19983));
    InMux I__1839 (
            .O(N__19990),
            .I(N__19976));
    InMux I__1838 (
            .O(N__19989),
            .I(N__19976));
    Span4Mux_v I__1837 (
            .O(N__19986),
            .I(N__19971));
    LocalMux I__1836 (
            .O(N__19983),
            .I(N__19971));
    InMux I__1835 (
            .O(N__19982),
            .I(N__19966));
    InMux I__1834 (
            .O(N__19981),
            .I(N__19966));
    LocalMux I__1833 (
            .O(N__19976),
            .I(\RTD.adress_7_N_1339_7 ));
    Odrv4 I__1832 (
            .O(N__19971),
            .I(\RTD.adress_7_N_1339_7 ));
    LocalMux I__1831 (
            .O(N__19966),
            .I(\RTD.adress_7_N_1339_7 ));
    InMux I__1830 (
            .O(N__19959),
            .I(N__19956));
    LocalMux I__1829 (
            .O(N__19956),
            .I(N__19953));
    Odrv12 I__1828 (
            .O(N__19953),
            .I(\RTD.n16638 ));
    CascadeMux I__1827 (
            .O(N__19950),
            .I(\RTD.n16638_cascade_ ));
    CascadeMux I__1826 (
            .O(N__19947),
            .I(N__19944));
    InMux I__1825 (
            .O(N__19944),
            .I(N__19941));
    LocalMux I__1824 (
            .O(N__19941),
            .I(N__19938));
    Span4Mux_h I__1823 (
            .O(N__19938),
            .I(N__19934));
    InMux I__1822 (
            .O(N__19937),
            .I(N__19931));
    Odrv4 I__1821 (
            .O(N__19934),
            .I(\RTD.n20787 ));
    LocalMux I__1820 (
            .O(N__19931),
            .I(\RTD.n20787 ));
    InMux I__1819 (
            .O(N__19926),
            .I(N__19923));
    LocalMux I__1818 (
            .O(N__19923),
            .I(\RTD.n17835 ));
    InMux I__1817 (
            .O(N__19920),
            .I(N__19917));
    LocalMux I__1816 (
            .O(N__19917),
            .I(\RTD.n7 ));
    CEMux I__1815 (
            .O(N__19914),
            .I(N__19911));
    LocalMux I__1814 (
            .O(N__19911),
            .I(N__19908));
    Span4Mux_h I__1813 (
            .O(N__19908),
            .I(N__19904));
    CEMux I__1812 (
            .O(N__19907),
            .I(N__19901));
    Odrv4 I__1811 (
            .O(N__19904),
            .I(\RTD.n11726 ));
    LocalMux I__1810 (
            .O(N__19901),
            .I(\RTD.n11726 ));
    InMux I__1809 (
            .O(N__19896),
            .I(N__19893));
    LocalMux I__1808 (
            .O(N__19893),
            .I(\RTD.n19787 ));
    CascadeMux I__1807 (
            .O(N__19890),
            .I(\RTD.n14_cascade_ ));
    InMux I__1806 (
            .O(N__19887),
            .I(N__19884));
    LocalMux I__1805 (
            .O(N__19884),
            .I(N__19881));
    Span4Mux_v I__1804 (
            .O(N__19881),
            .I(N__19877));
    InMux I__1803 (
            .O(N__19880),
            .I(N__19874));
    Odrv4 I__1802 (
            .O(N__19877),
            .I(\RTD.n20832 ));
    LocalMux I__1801 (
            .O(N__19874),
            .I(\RTD.n20832 ));
    CascadeMux I__1800 (
            .O(N__19869),
            .I(\RTD.n11704_cascade_ ));
    CascadeMux I__1799 (
            .O(N__19866),
            .I(N__19863));
    InMux I__1798 (
            .O(N__19863),
            .I(N__19857));
    InMux I__1797 (
            .O(N__19862),
            .I(N__19857));
    LocalMux I__1796 (
            .O(N__19857),
            .I(adress_4));
    CascadeMux I__1795 (
            .O(N__19854),
            .I(\RTD.n21362_cascade_ ));
    InMux I__1794 (
            .O(N__19851),
            .I(N__19847));
    InMux I__1793 (
            .O(N__19850),
            .I(N__19844));
    LocalMux I__1792 (
            .O(N__19847),
            .I(N__19839));
    LocalMux I__1791 (
            .O(N__19844),
            .I(N__19836));
    InMux I__1790 (
            .O(N__19843),
            .I(N__19833));
    InMux I__1789 (
            .O(N__19842),
            .I(N__19830));
    Span4Mux_h I__1788 (
            .O(N__19839),
            .I(N__19827));
    Odrv4 I__1787 (
            .O(N__19836),
            .I(\RTD.n1 ));
    LocalMux I__1786 (
            .O(N__19833),
            .I(\RTD.n1 ));
    LocalMux I__1785 (
            .O(N__19830),
            .I(\RTD.n1 ));
    Odrv4 I__1784 (
            .O(N__19827),
            .I(\RTD.n1 ));
    CascadeMux I__1783 (
            .O(N__19818),
            .I(N__19813));
    CascadeMux I__1782 (
            .O(N__19817),
            .I(N__19809));
    InMux I__1781 (
            .O(N__19816),
            .I(N__19805));
    InMux I__1780 (
            .O(N__19813),
            .I(N__19796));
    InMux I__1779 (
            .O(N__19812),
            .I(N__19796));
    InMux I__1778 (
            .O(N__19809),
            .I(N__19796));
    InMux I__1777 (
            .O(N__19808),
            .I(N__19796));
    LocalMux I__1776 (
            .O(N__19805),
            .I(n14479));
    LocalMux I__1775 (
            .O(N__19796),
            .I(n14479));
    CascadeMux I__1774 (
            .O(N__19791),
            .I(N__19788));
    InMux I__1773 (
            .O(N__19788),
            .I(N__19784));
    InMux I__1772 (
            .O(N__19787),
            .I(N__19781));
    LocalMux I__1771 (
            .O(N__19784),
            .I(adress_2));
    LocalMux I__1770 (
            .O(N__19781),
            .I(adress_2));
    CEMux I__1769 (
            .O(N__19776),
            .I(N__19773));
    LocalMux I__1768 (
            .O(N__19773),
            .I(N__19770));
    Span4Mux_h I__1767 (
            .O(N__19770),
            .I(N__19762));
    InMux I__1766 (
            .O(N__19769),
            .I(N__19759));
    InMux I__1765 (
            .O(N__19768),
            .I(N__19750));
    InMux I__1764 (
            .O(N__19767),
            .I(N__19750));
    InMux I__1763 (
            .O(N__19766),
            .I(N__19750));
    InMux I__1762 (
            .O(N__19765),
            .I(N__19750));
    Odrv4 I__1761 (
            .O(N__19762),
            .I(n13165));
    LocalMux I__1760 (
            .O(N__19759),
            .I(n13165));
    LocalMux I__1759 (
            .O(N__19750),
            .I(n13165));
    InMux I__1758 (
            .O(N__19743),
            .I(N__19740));
    LocalMux I__1757 (
            .O(N__19740),
            .I(N__19736));
    InMux I__1756 (
            .O(N__19739),
            .I(N__19733));
    Odrv4 I__1755 (
            .O(N__19736),
            .I(adress_3));
    LocalMux I__1754 (
            .O(N__19733),
            .I(adress_3));
    CEMux I__1753 (
            .O(N__19728),
            .I(N__19725));
    LocalMux I__1752 (
            .O(N__19725),
            .I(N__19722));
    Odrv12 I__1751 (
            .O(N__19722),
            .I(\RTD.n11687 ));
    InMux I__1750 (
            .O(N__19719),
            .I(N__19713));
    InMux I__1749 (
            .O(N__19718),
            .I(N__19713));
    LocalMux I__1748 (
            .O(N__19713),
            .I(adress_5));
    InMux I__1747 (
            .O(N__19710),
            .I(N__19706));
    InMux I__1746 (
            .O(N__19709),
            .I(N__19703));
    LocalMux I__1745 (
            .O(N__19706),
            .I(N__19698));
    LocalMux I__1744 (
            .O(N__19703),
            .I(N__19698));
    Odrv4 I__1743 (
            .O(N__19698),
            .I(adress_6));
    CascadeMux I__1742 (
            .O(N__19695),
            .I(\RTD.n19_cascade_ ));
    InMux I__1741 (
            .O(N__19692),
            .I(N__19689));
    LocalMux I__1740 (
            .O(N__19689),
            .I(N__19686));
    Span4Mux_v I__1739 (
            .O(N__19686),
            .I(N__19683));
    Odrv4 I__1738 (
            .O(N__19683),
            .I(adress_0));
    CascadeMux I__1737 (
            .O(N__19680),
            .I(n13165_cascade_));
    InMux I__1736 (
            .O(N__19677),
            .I(N__19673));
    InMux I__1735 (
            .O(N__19676),
            .I(N__19670));
    LocalMux I__1734 (
            .O(N__19673),
            .I(adress_1));
    LocalMux I__1733 (
            .O(N__19670),
            .I(adress_1));
    CascadeMux I__1732 (
            .O(N__19665),
            .I(n14479_cascade_));
    CascadeMux I__1731 (
            .O(N__19662),
            .I(n1_adj_1606_cascade_));
    SRMux I__1730 (
            .O(N__19659),
            .I(N__19655));
    SRMux I__1729 (
            .O(N__19658),
            .I(N__19652));
    LocalMux I__1728 (
            .O(N__19655),
            .I(N__19649));
    LocalMux I__1727 (
            .O(N__19652),
            .I(N__19646));
    Span4Mux_h I__1726 (
            .O(N__19649),
            .I(N__19643));
    Span4Mux_v I__1725 (
            .O(N__19646),
            .I(N__19640));
    Odrv4 I__1724 (
            .O(N__19643),
            .I(\RTD.n20160 ));
    Odrv4 I__1723 (
            .O(N__19640),
            .I(\RTD.n20160 ));
    InMux I__1722 (
            .O(N__19635),
            .I(N__19631));
    CascadeMux I__1721 (
            .O(N__19634),
            .I(N__19627));
    LocalMux I__1720 (
            .O(N__19631),
            .I(N__19624));
    InMux I__1719 (
            .O(N__19630),
            .I(N__19619));
    InMux I__1718 (
            .O(N__19627),
            .I(N__19619));
    Odrv4 I__1717 (
            .O(N__19624),
            .I(read_buf_3));
    LocalMux I__1716 (
            .O(N__19619),
            .I(read_buf_3));
    CascadeMux I__1715 (
            .O(N__19614),
            .I(N__19609));
    InMux I__1714 (
            .O(N__19613),
            .I(N__19606));
    InMux I__1713 (
            .O(N__19612),
            .I(N__19601));
    InMux I__1712 (
            .O(N__19609),
            .I(N__19601));
    LocalMux I__1711 (
            .O(N__19606),
            .I(read_buf_2));
    LocalMux I__1710 (
            .O(N__19601),
            .I(read_buf_2));
    IoInMux I__1709 (
            .O(N__19596),
            .I(N__19593));
    LocalMux I__1708 (
            .O(N__19593),
            .I(N__19590));
    Span4Mux_s2_v I__1707 (
            .O(N__19590),
            .I(N__19587));
    Span4Mux_v I__1706 (
            .O(N__19587),
            .I(N__19584));
    Odrv4 I__1705 (
            .O(N__19584),
            .I(DDS_MCLK1));
    IoInMux I__1704 (
            .O(N__19581),
            .I(N__19578));
    LocalMux I__1703 (
            .O(N__19578),
            .I(N__19575));
    Span4Mux_s3_h I__1702 (
            .O(N__19575),
            .I(N__19572));
    Sp12to4 I__1701 (
            .O(N__19572),
            .I(N__19569));
    Span12Mux_s10_v I__1700 (
            .O(N__19569),
            .I(N__19566));
    Odrv12 I__1699 (
            .O(N__19566),
            .I(RTD_CS));
    CascadeMux I__1698 (
            .O(N__19563),
            .I(\RTD.n4_cascade_ ));
    InMux I__1697 (
            .O(N__19560),
            .I(N__19556));
    InMux I__1696 (
            .O(N__19559),
            .I(N__19553));
    LocalMux I__1695 (
            .O(N__19556),
            .I(\RTD.cfg_buf_7 ));
    LocalMux I__1694 (
            .O(N__19553),
            .I(\RTD.cfg_buf_7 ));
    InMux I__1693 (
            .O(N__19548),
            .I(N__19544));
    InMux I__1692 (
            .O(N__19547),
            .I(N__19541));
    LocalMux I__1691 (
            .O(N__19544),
            .I(cfg_buf_1));
    LocalMux I__1690 (
            .O(N__19541),
            .I(cfg_buf_1));
    InMux I__1689 (
            .O(N__19536),
            .I(N__19533));
    LocalMux I__1688 (
            .O(N__19533),
            .I(N__19530));
    Odrv4 I__1687 (
            .O(N__19530),
            .I(\RTD.n12 ));
    InMux I__1686 (
            .O(N__19527),
            .I(N__19524));
    LocalMux I__1685 (
            .O(N__19524),
            .I(\RTD.n11 ));
    InMux I__1684 (
            .O(N__19521),
            .I(N__19518));
    LocalMux I__1683 (
            .O(N__19518),
            .I(\RTD.n11_adj_1403 ));
    CascadeMux I__1682 (
            .O(N__19515),
            .I(N__19512));
    InMux I__1681 (
            .O(N__19512),
            .I(N__19509));
    LocalMux I__1680 (
            .O(N__19509),
            .I(\RTD.n32 ));
    CascadeMux I__1679 (
            .O(N__19506),
            .I(\RTD.n32_cascade_ ));
    InMux I__1678 (
            .O(N__19503),
            .I(N__19500));
    LocalMux I__1677 (
            .O(N__19500),
            .I(\RTD.n21555 ));
    InMux I__1676 (
            .O(N__19497),
            .I(N__19494));
    LocalMux I__1675 (
            .O(N__19494),
            .I(\RTD.n6 ));
    CascadeMux I__1674 (
            .O(N__19491),
            .I(N__19488));
    InMux I__1673 (
            .O(N__19488),
            .I(N__19485));
    LocalMux I__1672 (
            .O(N__19485),
            .I(N__19482));
    Span12Mux_s7_h I__1671 (
            .O(N__19482),
            .I(N__19479));
    Span12Mux_v I__1670 (
            .O(N__19479),
            .I(N__19476));
    Odrv12 I__1669 (
            .O(N__19476),
            .I(RTD_SDO));
    CascadeMux I__1668 (
            .O(N__19473),
            .I(N__19470));
    InMux I__1667 (
            .O(N__19470),
            .I(N__19467));
    LocalMux I__1666 (
            .O(N__19467),
            .I(N__19463));
    InMux I__1665 (
            .O(N__19466),
            .I(N__19460));
    Odrv4 I__1664 (
            .O(N__19463),
            .I(\RTD.cfg_buf_6 ));
    LocalMux I__1663 (
            .O(N__19460),
            .I(\RTD.cfg_buf_6 ));
    CascadeMux I__1662 (
            .O(N__19455),
            .I(N__19452));
    InMux I__1661 (
            .O(N__19452),
            .I(N__19448));
    InMux I__1660 (
            .O(N__19451),
            .I(N__19445));
    LocalMux I__1659 (
            .O(N__19448),
            .I(cfg_buf_0));
    LocalMux I__1658 (
            .O(N__19445),
            .I(cfg_buf_0));
    CascadeMux I__1657 (
            .O(N__19440),
            .I(\RTD.n9_cascade_ ));
    CascadeMux I__1656 (
            .O(N__19437),
            .I(\RTD.adress_7_N_1339_7_cascade_ ));
    InMux I__1655 (
            .O(N__19434),
            .I(N__19430));
    InMux I__1654 (
            .O(N__19433),
            .I(N__19427));
    LocalMux I__1653 (
            .O(N__19430),
            .I(\RTD.cfg_buf_5 ));
    LocalMux I__1652 (
            .O(N__19427),
            .I(\RTD.cfg_buf_5 ));
    InMux I__1651 (
            .O(N__19422),
            .I(N__19418));
    InMux I__1650 (
            .O(N__19421),
            .I(N__19415));
    LocalMux I__1649 (
            .O(N__19418),
            .I(\RTD.cfg_buf_3 ));
    LocalMux I__1648 (
            .O(N__19415),
            .I(\RTD.cfg_buf_3 ));
    InMux I__1647 (
            .O(N__19410),
            .I(N__19407));
    LocalMux I__1646 (
            .O(N__19407),
            .I(\RTD.n11_adj_1405 ));
    CascadeMux I__1645 (
            .O(N__19404),
            .I(N__19401));
    InMux I__1644 (
            .O(N__19401),
            .I(N__19397));
    InMux I__1643 (
            .O(N__19400),
            .I(N__19394));
    LocalMux I__1642 (
            .O(N__19397),
            .I(\RTD.cfg_buf_4 ));
    LocalMux I__1641 (
            .O(N__19394),
            .I(\RTD.cfg_buf_4 ));
    CascadeMux I__1640 (
            .O(N__19389),
            .I(N__19386));
    InMux I__1639 (
            .O(N__19386),
            .I(N__19382));
    InMux I__1638 (
            .O(N__19385),
            .I(N__19379));
    LocalMux I__1637 (
            .O(N__19382),
            .I(\RTD.cfg_buf_2 ));
    LocalMux I__1636 (
            .O(N__19379),
            .I(\RTD.cfg_buf_2 ));
    InMux I__1635 (
            .O(N__19374),
            .I(N__19371));
    LocalMux I__1634 (
            .O(N__19371),
            .I(\RTD.n10 ));
    InMux I__1633 (
            .O(N__19368),
            .I(N__19364));
    InMux I__1632 (
            .O(N__19367),
            .I(N__19361));
    LocalMux I__1631 (
            .O(N__19364),
            .I(\RTD.adress_7 ));
    LocalMux I__1630 (
            .O(N__19361),
            .I(\RTD.adress_7 ));
    InMux I__1629 (
            .O(N__19356),
            .I(N__19353));
    LocalMux I__1628 (
            .O(N__19353),
            .I(N__19350));
    Odrv4 I__1627 (
            .O(N__19350),
            .I(\RTD.n7318 ));
    CascadeMux I__1626 (
            .O(N__19347),
            .I(\RTD.n7318_cascade_ ));
    CascadeMux I__1625 (
            .O(N__19344),
            .I(\RTD.n21_cascade_ ));
    CascadeMux I__1624 (
            .O(N__19341),
            .I(n13176_cascade_));
    InMux I__1623 (
            .O(N__19338),
            .I(N__19319));
    InMux I__1622 (
            .O(N__19337),
            .I(N__19319));
    InMux I__1621 (
            .O(N__19336),
            .I(N__19319));
    InMux I__1620 (
            .O(N__19335),
            .I(N__19319));
    InMux I__1619 (
            .O(N__19334),
            .I(N__19319));
    InMux I__1618 (
            .O(N__19333),
            .I(N__19319));
    InMux I__1617 (
            .O(N__19332),
            .I(N__19316));
    LocalMux I__1616 (
            .O(N__19319),
            .I(n18755));
    LocalMux I__1615 (
            .O(N__19316),
            .I(n18755));
    CascadeMux I__1614 (
            .O(N__19311),
            .I(N__19306));
    CascadeMux I__1613 (
            .O(N__19310),
            .I(N__19303));
    CascadeMux I__1612 (
            .O(N__19309),
            .I(N__19298));
    InMux I__1611 (
            .O(N__19306),
            .I(N__19282));
    InMux I__1610 (
            .O(N__19303),
            .I(N__19282));
    InMux I__1609 (
            .O(N__19302),
            .I(N__19282));
    InMux I__1608 (
            .O(N__19301),
            .I(N__19282));
    InMux I__1607 (
            .O(N__19298),
            .I(N__19282));
    InMux I__1606 (
            .O(N__19297),
            .I(N__19282));
    InMux I__1605 (
            .O(N__19296),
            .I(N__19277));
    InMux I__1604 (
            .O(N__19295),
            .I(N__19277));
    LocalMux I__1603 (
            .O(N__19282),
            .I(n13176));
    LocalMux I__1602 (
            .O(N__19277),
            .I(n13176));
    CascadeMux I__1601 (
            .O(N__19272),
            .I(n18755_cascade_));
    InMux I__1600 (
            .O(N__19269),
            .I(N__19266));
    LocalMux I__1599 (
            .O(N__19266),
            .I(\RTD.n16 ));
    CEMux I__1598 (
            .O(N__19263),
            .I(N__19260));
    LocalMux I__1597 (
            .O(N__19260),
            .I(N__19257));
    Odrv12 I__1596 (
            .O(N__19257),
            .I(\RTD.n8 ));
    IoInMux I__1595 (
            .O(N__19254),
            .I(N__19251));
    LocalMux I__1594 (
            .O(N__19251),
            .I(N__19248));
    Span4Mux_s0_h I__1593 (
            .O(N__19248),
            .I(N__19245));
    Sp12to4 I__1592 (
            .O(N__19245),
            .I(N__19242));
    Span12Mux_v I__1591 (
            .O(N__19242),
            .I(N__19239));
    Odrv12 I__1590 (
            .O(N__19239),
            .I(RTD_SDI));
    CEMux I__1589 (
            .O(N__19236),
            .I(N__19233));
    LocalMux I__1588 (
            .O(N__19233),
            .I(N__19230));
    Span4Mux_h I__1587 (
            .O(N__19230),
            .I(N__19227));
    Odrv4 I__1586 (
            .O(N__19227),
            .I(\RTD.n11718 ));
    IoInMux I__1585 (
            .O(N__19224),
            .I(N__19221));
    LocalMux I__1584 (
            .O(N__19221),
            .I(N__19218));
    IoSpan4Mux I__1583 (
            .O(N__19218),
            .I(N__19215));
    IoSpan4Mux I__1582 (
            .O(N__19215),
            .I(N__19212));
    Span4Mux_s2_h I__1581 (
            .O(N__19212),
            .I(N__19209));
    Odrv4 I__1580 (
            .O(N__19209),
            .I(RTD_SCLK));
    IoInMux I__1579 (
            .O(N__19206),
            .I(N__19203));
    LocalMux I__1578 (
            .O(N__19203),
            .I(N__19200));
    IoSpan4Mux I__1577 (
            .O(N__19200),
            .I(N__19197));
    IoSpan4Mux I__1576 (
            .O(N__19197),
            .I(N__19194));
    Odrv4 I__1575 (
            .O(N__19194),
            .I(ICE_SYSCLK));
    IoInMux I__1574 (
            .O(N__19191),
            .I(N__19188));
    LocalMux I__1573 (
            .O(N__19188),
            .I(N__19185));
    IoSpan4Mux I__1572 (
            .O(N__19185),
            .I(N__19182));
    Span4Mux_s3_v I__1571 (
            .O(N__19182),
            .I(N__19179));
    Sp12to4 I__1570 (
            .O(N__19179),
            .I(N__19176));
    Span12Mux_h I__1569 (
            .O(N__19176),
            .I(N__19173));
    Odrv12 I__1568 (
            .O(N__19173),
            .I(ICE_GPMO_2));
    INV \INVADC_VDC.genclk.t0on_i8C  (
            .O(\INVADC_VDC.genclk.t0on_i8C_net ),
            .I(N__38755));
    INV \INVADC_VDC.genclk.t0on_i0C  (
            .O(\INVADC_VDC.genclk.t0on_i0C_net ),
            .I(N__38754));
    INV \INVADC_VDC.genclk.div_state_i0C  (
            .O(\INVADC_VDC.genclk.div_state_i0C_net ),
            .I(N__38753));
    INV \INVADC_VDC.genclk.div_state_i1C  (
            .O(\INVADC_VDC.genclk.div_state_i1C_net ),
            .I(N__38749));
    INV \INVADC_VDC.genclk.t0off_i8C  (
            .O(\INVADC_VDC.genclk.t0off_i8C_net ),
            .I(N__38752));
    INV \INVADC_VDC.genclk.t0off_i0C  (
            .O(\INVADC_VDC.genclk.t0off_i0C_net ),
            .I(N__38750));
    INV INVdata_cntvec_i0_i8C (
            .O(INVdata_cntvec_i0_i8C_net),
            .I(N__54400));
    INV INVdata_cntvec_i0_i0C (
            .O(INVdata_cntvec_i0_i0C_net),
            .I(N__54388));
    INV \INVcomm_spi.data_valid_85C  (
            .O(\INVcomm_spi.data_valid_85C_net ),
            .I(N__54295));
    INV INVacadc_skipcnt_i0_i9C (
            .O(INVacadc_skipcnt_i0_i9C_net),
            .I(N__54393));
    INV INVacadc_skipcnt_i0_i1C (
            .O(INVacadc_skipcnt_i0_i1C_net),
            .I(N__54381));
    INV INVacadc_skipcnt_i0_i0C (
            .O(INVacadc_skipcnt_i0_i0C_net),
            .I(N__54366));
    INV \INVcomm_spi.imiso_83_12192_12193_setC  (
            .O(\INVcomm_spi.imiso_83_12192_12193_setC_net ),
            .I(N__52601));
    INV INVdds0_mclk_294C (
            .O(INVdds0_mclk_294C_net),
            .I(N__38745));
    INV \INVcomm_spi.MISO_48_12186_12187_setC  (
            .O(\INVcomm_spi.MISO_48_12186_12187_setC_net ),
            .I(N__54271));
    INV \INVcomm_spi.imiso_83_12192_12193_resetC  (
            .O(\INVcomm_spi.imiso_83_12192_12193_resetC_net ),
            .I(N__52502));
    INV INVdds0_mclkcnt_i7_3772__i0C (
            .O(INVdds0_mclkcnt_i7_3772__i0C_net),
            .I(N__38739));
    INV INVeis_state_i2C (
            .O(INVeis_state_i2C_net),
            .I(N__54398));
    INV INVeis_end_299C (
            .O(INVeis_end_299C_net),
            .I(N__54359));
    INV INVdata_count_i0_i8C (
            .O(INVdata_count_i0_i8C_net),
            .I(N__54331));
    INV INVdata_count_i0_i0C (
            .O(INVdata_count_i0_i0C_net),
            .I(N__54318));
    INV \INVcomm_spi.MISO_48_12186_12187_resetC  (
            .O(\INVcomm_spi.MISO_48_12186_12187_resetC_net ),
            .I(N__54269));
    INV INVeis_state_i0C (
            .O(INVeis_state_i0C_net),
            .I(N__54384));
    INV \INVcomm_spi.bit_cnt_3767__i3C  (
            .O(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .I(N__52498));
    INV INVacadc_trig_300C (
            .O(INVacadc_trig_300C_net),
            .I(N__54412));
    INV INViac_raw_buf_vac_raw_buf_merged2WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .I(N__54380));
    INV INViac_raw_buf_vac_raw_buf_merged7WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .I(N__54438));
    INV INViac_raw_buf_vac_raw_buf_merged1WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .I(N__54298));
    INV INViac_raw_buf_vac_raw_buf_merged6WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .I(N__54436));
    INV INViac_raw_buf_vac_raw_buf_merged0WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .I(N__54285));
    INV INViac_raw_buf_vac_raw_buf_merged5WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .I(N__54434));
    INV INViac_raw_buf_vac_raw_buf_merged9WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .I(N__54338));
    INV INViac_raw_buf_vac_raw_buf_merged4WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .I(N__54426));
    INV INViac_raw_buf_vac_raw_buf_merged8WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .I(N__54312));
    INV INViac_raw_buf_vac_raw_buf_merged10WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .I(N__54326));
    INV INViac_raw_buf_vac_raw_buf_merged3WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .I(N__54407));
    INV INViac_raw_buf_vac_raw_buf_merged11WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .I(N__54352));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(n19757),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(n19765),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(n19610_THRU_CRY_6_THRU_CO),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(n19618),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(n19602),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(n19593),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(n19641),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(n19632),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_19_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_8_0_ (
            .carryinitin(\ADC_VDC.genclk.n19716 ),
            .carryinitout(bfn_19_8_0_));
    defparam IN_MUX_bfv_22_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_7_0_));
    defparam IN_MUX_bfv_22_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_8_0_ (
            .carryinitin(\ADC_VDC.genclk.n19731 ),
            .carryinitout(bfn_22_8_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(\ADC_VDC.n19705 ),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\ADC_VDC.n19670 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\ADC_VDC.n19678 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\ADC_VDC.n19686 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\ADC_VDC.n19694 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \RTD.SCLK_51_LC_2_5_3 .C_ON=1'b0;
    defparam \RTD.SCLK_51_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \RTD.SCLK_51_LC_2_5_3 .LUT_INIT=16'b0100010110100110;
    LogicCell40 \RTD.SCLK_51_LC_2_5_3  (
            .in0(N__26783),
            .in1(N__26596),
            .in2(N__26277),
            .in3(N__26415),
            .lcout(RTD_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30472),
            .ce(N__19263),
            .sr(_gnd_net_));
    defparam \RTD.i19375_4_lut_4_lut_LC_2_6_0 .C_ON=1'b0;
    defparam \RTD.i19375_4_lut_4_lut_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i19375_4_lut_4_lut_LC_2_6_0 .LUT_INIT=16'b1011111111011111;
    LogicCell40 \RTD.i19375_4_lut_4_lut_LC_2_6_0  (
            .in0(N__26782),
            .in1(N__26559),
            .in2(N__26441),
            .in3(N__26272),
            .lcout(\RTD.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i7_LC_2_7_0 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i7_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i7_LC_2_7_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \RTD.cfg_buf_i7_LC_2_7_0  (
            .in0(N__19338),
            .in1(N__31301),
            .in2(N__19311),
            .in3(N__19560),
            .lcout(\RTD.cfg_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30518),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_40_LC_2_7_2 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_40_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_40_LC_2_7_2 .LUT_INIT=16'b1110000010000000;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_40_LC_2_7_2  (
            .in0(N__26533),
            .in1(N__26735),
            .in2(N__26391),
            .in3(N__26271),
            .lcout(n11714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i4_LC_2_7_3 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i4_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i4_LC_2_7_3 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \RTD.cfg_buf_i4_LC_2_7_3  (
            .in0(N__22782),
            .in1(N__19302),
            .in2(N__19404),
            .in3(N__19336),
            .lcout(\RTD.cfg_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30518),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i5_LC_2_7_4 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i5_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i5_LC_2_7_4 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \RTD.cfg_buf_i5_LC_2_7_4  (
            .in0(N__19337),
            .in1(N__21821),
            .in2(N__19310),
            .in3(N__19434),
            .lcout(\RTD.cfg_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30518),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i2_LC_2_7_5 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i2_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i2_LC_2_7_5 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \RTD.cfg_buf_i2_LC_2_7_5  (
            .in0(N__21882),
            .in1(N__19301),
            .in2(N__19389),
            .in3(N__19335),
            .lcout(\RTD.cfg_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30518),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i1_LC_2_7_6 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i1_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i1_LC_2_7_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \RTD.cfg_buf_i1_LC_2_7_6  (
            .in0(N__19334),
            .in1(N__21180),
            .in2(N__19309),
            .in3(N__19548),
            .lcout(cfg_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30518),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i0_LC_2_7_7 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i0_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i0_LC_2_7_7 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \RTD.cfg_buf_i0_LC_2_7_7  (
            .in0(N__23261),
            .in1(N__19297),
            .in2(N__19455),
            .in3(N__19333),
            .lcout(cfg_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30518),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.MOSI_59_LC_2_8_1 .C_ON=1'b0;
    defparam \RTD.MOSI_59_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.MOSI_59_LC_2_8_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \RTD.MOSI_59_LC_2_8_1  (
            .in0(N__19367),
            .in1(N__26778),
            .in2(N__20154),
            .in3(N__26273),
            .lcout(RTD_SDI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30508),
            .ce(N__19236),
            .sr(N__19659));
    defparam \RTD.i27_4_lut_4_lut_LC_2_9_6 .C_ON=1'b0;
    defparam \RTD.i27_4_lut_4_lut_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i27_4_lut_4_lut_LC_2_9_6 .LUT_INIT=16'b1010101010000110;
    LogicCell40 \RTD.i27_4_lut_4_lut_LC_2_9_6  (
            .in0(N__26724),
            .in1(N__26541),
            .in2(N__26421),
            .in3(N__26252),
            .lcout(\RTD.n11718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i2_LC_2_11_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i2_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i2_LC_2_11_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i2_LC_2_11_3  (
            .in0(N__19613),
            .in1(N__21639),
            .in2(N__46664),
            .in3(N__26836),
            .lcout(buf_readRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30528),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i6_LC_3_6_0 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i6_LC_3_6_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i6_LC_3_6_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \RTD.cfg_buf_i6_LC_3_6_0  (
            .in0(N__31378),
            .in1(N__19296),
            .in2(N__19473),
            .in3(N__19332),
            .lcout(\RTD.cfg_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30509),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_34_LC_3_6_2 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_34_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_34_LC_3_6_2 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \RTD.i1_4_lut_adj_34_LC_3_6_2  (
            .in0(N__26268),
            .in1(N__19356),
            .in2(N__20041),
            .in3(N__19981),
            .lcout(),
            .ltout(\RTD.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_35_LC_3_6_3 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_35_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_35_LC_3_6_3 .LUT_INIT=16'b0010000010101000;
    LogicCell40 \RTD.i1_4_lut_adj_35_LC_3_6_3  (
            .in0(N__20056),
            .in1(N__26426),
            .in2(N__19344),
            .in3(N__26750),
            .lcout(\RTD.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i22_4_lut_4_lut_LC_3_6_4 .C_ON=1'b0;
    defparam \RTD.i22_4_lut_4_lut_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i22_4_lut_4_lut_LC_3_6_4 .LUT_INIT=16'b1000010110000000;
    LogicCell40 \RTD.i22_4_lut_4_lut_LC_3_6_4  (
            .in0(N__26749),
            .in1(N__19851),
            .in2(N__26443),
            .in3(N__19880),
            .lcout(n13176),
            .ltout(n13176_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_3_lut_LC_3_6_5 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_LC_3_6_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_LC_3_6_5 .LUT_INIT=16'b0011111100001111;
    LogicCell40 \RTD.i1_3_lut_LC_3_6_5  (
            .in0(_gnd_net_),
            .in1(N__26425),
            .in2(N__19341),
            .in3(N__26269),
            .lcout(n18755),
            .ltout(n18755_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i3_LC_3_6_6 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i3_LC_3_6_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i3_LC_3_6_6 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \RTD.cfg_buf_i3_LC_3_6_6  (
            .in0(N__24692),
            .in1(N__19295),
            .in2(N__19272),
            .in3(N__19422),
            .lcout(\RTD.cfg_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30509),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.mode_53_LC_3_6_7 .C_ON=1'b0;
    defparam \RTD.mode_53_LC_3_6_7 .SEQ_MODE=4'b1000;
    defparam \RTD.mode_53_LC_3_6_7 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \RTD.mode_53_LC_3_6_7  (
            .in0(N__19982),
            .in1(N__26270),
            .in2(N__19947),
            .in3(N__19269),
            .lcout(\RTD.mode ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30509),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i7_LC_3_7_0 .C_ON=1'b0;
    defparam \RTD.adress_i7_LC_3_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i7_LC_3_7_0 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \RTD.adress_i7_LC_3_7_0  (
            .in0(N__19990),
            .in1(N__19710),
            .in2(N__26585),
            .in3(N__26260),
            .lcout(\RTD.adress_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30517),
            .ce(N__19776),
            .sr(N__19658));
    defparam \RTD.i1_4_lut_adj_37_LC_3_7_1 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_37_LC_3_7_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_37_LC_3_7_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i1_4_lut_adj_37_LC_3_7_1  (
            .in0(N__31386),
            .in1(N__19466),
            .in2(N__23262),
            .in3(N__19451),
            .lcout(),
            .ltout(\RTD.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i7_4_lut_LC_3_7_2 .C_ON=1'b0;
    defparam \RTD.i7_4_lut_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i7_4_lut_LC_3_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \RTD.i7_4_lut_LC_3_7_2  (
            .in0(N__19536),
            .in1(N__19374),
            .in2(N__19440),
            .in3(N__19410),
            .lcout(\RTD.adress_7_N_1339_7 ),
            .ltout(\RTD.adress_7_N_1339_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_LC_3_7_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_LC_3_7_3 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \RTD.i1_2_lut_3_lut_LC_3_7_3  (
            .in0(N__26258),
            .in1(_gnd_net_),
            .in2(N__19437),
            .in3(N__26544),
            .lcout(\RTD.n20832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i3_4_lut_LC_3_7_4 .C_ON=1'b0;
    defparam \RTD.i3_4_lut_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i3_4_lut_LC_3_7_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \RTD.i3_4_lut_LC_3_7_4  (
            .in0(N__19433),
            .in1(N__24691),
            .in2(N__21822),
            .in3(N__19421),
            .lcout(\RTD.n11_adj_1405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_4_lut_LC_3_7_5 .C_ON=1'b0;
    defparam \RTD.i2_4_lut_LC_3_7_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_4_lut_LC_3_7_5 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i2_4_lut_LC_3_7_5  (
            .in0(N__22777),
            .in1(N__19400),
            .in2(N__21881),
            .in3(N__19385),
            .lcout(\RTD.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i0_LC_3_7_6 .C_ON=1'b0;
    defparam \RTD.adress_i0_LC_3_7_6 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i0_LC_3_7_6 .LUT_INIT=16'b1100010111001111;
    LogicCell40 \RTD.adress_i0_LC_3_7_6  (
            .in0(N__19989),
            .in1(N__19368),
            .in2(N__26584),
            .in3(N__26259),
            .lcout(adress_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30517),
            .ce(N__19776),
            .sr(N__19658));
    defparam \RTD.adc_state_i2_LC_3_8_0 .C_ON=1'b0;
    defparam \RTD.adc_state_i2_LC_3_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i2_LC_3_8_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \RTD.adc_state_i2_LC_3_8_0  (
            .in0(N__26764),
            .in1(N__19850),
            .in2(N__26427),
            .in3(N__19503),
            .lcout(adc_state_2_adj_1481),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30525),
            .ce(N__19914),
            .sr(_gnd_net_));
    defparam \RTD.i4903_2_lut_LC_3_8_1 .C_ON=1'b0;
    defparam \RTD.i4903_2_lut_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i4903_2_lut_LC_3_8_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i4903_2_lut_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(N__26762),
            .in2(_gnd_net_),
            .in3(N__26534),
            .lcout(\RTD.n7318 ),
            .ltout(\RTD.n7318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i1_LC_3_8_2 .C_ON=1'b0;
    defparam \RTD.adc_state_i1_LC_3_8_2 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i1_LC_3_8_2 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \RTD.adc_state_i1_LC_3_8_2  (
            .in0(N__26381),
            .in1(N__19521),
            .in2(N__19347),
            .in3(N__26263),
            .lcout(\RTD.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30525),
            .ce(N__19914),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_LC_3_8_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_LC_3_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RTD.i1_2_lut_LC_3_8_3  (
            .in0(_gnd_net_),
            .in1(N__26535),
            .in2(_gnd_net_),
            .in3(N__20585),
            .lcout(),
            .ltout(\RTD.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i3_LC_3_8_4 .C_ON=1'b0;
    defparam \RTD.adc_state_i3_LC_3_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i3_LC_3_8_4 .LUT_INIT=16'b0101010111000000;
    LogicCell40 \RTD.adc_state_i3_LC_3_8_4  (
            .in0(N__26763),
            .in1(N__19527),
            .in2(N__19563),
            .in3(N__26385),
            .lcout(\RTD.adc_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30525),
            .ce(N__19914),
            .sr(_gnd_net_));
    defparam \RTD.i4_4_lut_LC_3_8_7 .C_ON=1'b0;
    defparam \RTD.i4_4_lut_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i4_4_lut_LC_3_8_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i4_4_lut_LC_3_8_7  (
            .in0(N__21179),
            .in1(N__19559),
            .in2(N__31300),
            .in3(N__19547),
            .lcout(\RTD.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i22_4_lut_LC_3_9_1 .C_ON=1'b0;
    defparam \RTD.i22_4_lut_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i22_4_lut_LC_3_9_1 .LUT_INIT=16'b0000000001000110;
    LogicCell40 \RTD.i22_4_lut_LC_3_9_1  (
            .in0(N__26261),
            .in1(N__26726),
            .in2(N__20072),
            .in3(N__20553),
            .lcout(\RTD.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i24_4_lut_4_lut_LC_3_9_2 .C_ON=1'b0;
    defparam \RTD.i24_4_lut_4_lut_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i24_4_lut_4_lut_LC_3_9_2 .LUT_INIT=16'b1010101011100110;
    LogicCell40 \RTD.i24_4_lut_4_lut_LC_3_9_2  (
            .in0(N__26725),
            .in1(N__26543),
            .in2(N__19515),
            .in3(N__26262),
            .lcout(\RTD.n11_adj_1403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_23_LC_3_9_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_23_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_23_LC_3_9_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \RTD.i1_2_lut_adj_23_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(N__20552),
            .in2(_gnd_net_),
            .in3(N__20586),
            .lcout(\RTD.n32 ),
            .ltout(\RTD.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19313_4_lut_LC_3_9_4 .C_ON=1'b0;
    defparam \RTD.i19313_4_lut_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i19313_4_lut_LC_3_9_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \RTD.i19313_4_lut_LC_3_9_4  (
            .in0(N__26380),
            .in1(N__19497),
            .in2(N__19506),
            .in3(N__20068),
            .lcout(\RTD.n21555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_31_LC_3_9_6 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_31_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_31_LC_3_9_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \RTD.i1_2_lut_adj_31_LC_3_9_6  (
            .in0(N__26251),
            .in1(N__26542),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RTD.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i0_LC_3_10_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i0_LC_3_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i0_LC_3_10_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.read_buf_i0_LC_3_10_0  (
            .in0(N__20261),
            .in1(N__20950),
            .in2(N__19491),
            .in3(N__20861),
            .lcout(read_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30526),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_adj_26_LC_3_10_2 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_adj_26_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_adj_26_LC_3_10_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \RTD.i2_3_lut_adj_26_LC_3_10_2  (
            .in0(N__26419),
            .in1(_gnd_net_),
            .in2(N__26837),
            .in3(N__26267),
            .lcout(n1_adj_1606),
            .ltout(n1_adj_1606_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i4_LC_3_10_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i4_LC_3_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i4_LC_3_10_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i4_LC_3_10_3  (
            .in0(N__20860),
            .in1(N__20092),
            .in2(N__19662),
            .in3(N__19635),
            .lcout(read_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30526),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_39_LC_3_10_4 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_39_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_39_LC_3_10_4 .LUT_INIT=16'b1011000010010001;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_39_LC_3_10_4  (
            .in0(N__26784),
            .in1(N__26580),
            .in2(N__26442),
            .in3(N__26266),
            .lcout(n13293),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_5 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_5  (
            .in0(N__26265),
            .in1(N__26785),
            .in2(N__26597),
            .in3(N__26420),
            .lcout(\RTD.n20160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i3_LC_3_11_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i3_LC_3_11_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i3_LC_3_11_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i3_LC_3_11_0  (
            .in0(N__19612),
            .in1(N__20952),
            .in2(N__19634),
            .in3(N__20863),
            .lcout(read_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30527),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i3_LC_3_11_2 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i3_LC_3_11_2 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i3_LC_3_11_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i3_LC_3_11_2  (
            .in0(N__19630),
            .in1(N__21670),
            .in2(N__50141),
            .in3(N__26815),
            .lcout(buf_readRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30527),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i2_LC_3_11_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i2_LC_3_11_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i2_LC_3_11_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i2_LC_3_11_4  (
            .in0(N__20250),
            .in1(N__20951),
            .in2(N__19614),
            .in3(N__20862),
            .lcout(read_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30527),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_main.i19883_1_lut_LC_5_1_5 .C_ON=1'b0;
    defparam \pll_main.i19883_1_lut_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \pll_main.i19883_1_lut_LC_5_1_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_main.i19883_1_lut_LC_5_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38765),
            .lcout(DDS_MCLK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.CS_52_LC_5_5_1 .C_ON=1'b0;
    defparam \RTD.CS_52_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \RTD.CS_52_LC_5_5_1 .LUT_INIT=16'b0000001101011111;
    LogicCell40 \RTD.CS_52_LC_5_5_1  (
            .in0(N__26593),
            .in1(N__19959),
            .in2(N__26447),
            .in3(N__26257),
            .lcout(RTD_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30416),
            .ce(N__19728),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i2_LC_5_6_2 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i2_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i2_LC_5_6_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \CLK_DDS.dds_state_i2_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__34750),
            .in2(_gnd_net_),
            .in3(N__34529),
            .lcout(dds_state_2_adj_1452),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54313),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19332_3_lut_3_lut_LC_5_6_4 .C_ON=1'b0;
    defparam \RTD.i19332_3_lut_3_lut_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i19332_3_lut_3_lut_LC_5_6_4 .LUT_INIT=16'b1000100010011001;
    LogicCell40 \RTD.i19332_3_lut_3_lut_LC_5_6_4  (
            .in0(N__26435),
            .in1(N__26829),
            .in2(_gnd_net_),
            .in3(N__26592),
            .lcout(\RTD.n11687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i4_LC_5_6_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i4_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i4_LC_5_6_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i4_LC_5_6_7  (
            .in0(N__33680),
            .in1(N__33388),
            .in2(N__28296),
            .in3(N__20429),
            .lcout(buf_adcdata_vac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54313),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i5_LC_5_7_0 .C_ON=1'b0;
    defparam \RTD.adress_i5_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i5_LC_5_7_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i5_LC_5_7_0  (
            .in0(N__19718),
            .in1(N__19812),
            .in2(N__19866),
            .in3(N__19767),
            .lcout(adress_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30467),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i6_LC_5_7_1 .C_ON=1'b0;
    defparam \RTD.adress_i6_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i6_LC_5_7_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.adress_i6_LC_5_7_1  (
            .in0(N__19768),
            .in1(N__19719),
            .in2(N__19818),
            .in3(N__19709),
            .lcout(adress_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30467),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i34_4_lut_4_lut_LC_5_7_2 .C_ON=1'b0;
    defparam \RTD.i34_4_lut_4_lut_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i34_4_lut_4_lut_LC_5_7_2 .LUT_INIT=16'b1101110110011101;
    LogicCell40 \RTD.i34_4_lut_4_lut_LC_5_7_2  (
            .in0(N__26594),
            .in1(N__26253),
            .in2(N__20042),
            .in3(N__19991),
            .lcout(),
            .ltout(\RTD.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i35_4_lut_4_lut_LC_5_7_3 .C_ON=1'b0;
    defparam \RTD.i35_4_lut_4_lut_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i35_4_lut_4_lut_LC_5_7_3 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \RTD.i35_4_lut_4_lut_LC_5_7_3  (
            .in0(N__26830),
            .in1(N__26436),
            .in2(N__19695),
            .in3(N__19843),
            .lcout(n13165),
            .ltout(n13165_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i1_LC_5_7_4 .C_ON=1'b0;
    defparam \RTD.adress_i1_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i1_LC_5_7_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \RTD.adress_i1_LC_5_7_4  (
            .in0(N__19692),
            .in1(N__19676),
            .in2(N__19680),
            .in3(N__19808),
            .lcout(adress_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30467),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12067_2_lut_LC_5_7_5 .C_ON=1'b0;
    defparam \RTD.i12067_2_lut_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i12067_2_lut_LC_5_7_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \RTD.i12067_2_lut_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(N__26437),
            .in2(_gnd_net_),
            .in3(N__26595),
            .lcout(n14479),
            .ltout(n14479_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i2_LC_5_7_6 .C_ON=1'b0;
    defparam \RTD.adress_i2_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i2_LC_5_7_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \RTD.adress_i2_LC_5_7_6  (
            .in0(N__19677),
            .in1(N__19787),
            .in2(N__19665),
            .in3(N__19765),
            .lcout(adress_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30467),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i4_LC_5_7_7 .C_ON=1'b0;
    defparam \RTD.adress_i4_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i4_LC_5_7_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.adress_i4_LC_5_7_7  (
            .in0(N__19766),
            .in1(N__19743),
            .in2(N__19817),
            .in3(N__19862),
            .lcout(adress_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30467),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_2_lut_3_lut_LC_5_8_0 .C_ON=1'b0;
    defparam \RTD.i2_2_lut_3_lut_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_2_lut_3_lut_LC_5_8_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \RTD.i2_2_lut_3_lut_LC_5_8_0  (
            .in0(N__26389),
            .in1(N__26760),
            .in2(_gnd_net_),
            .in3(N__26561),
            .lcout(\RTD.n20787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19242_3_lut_LC_5_8_1 .C_ON=1'b0;
    defparam \RTD.i19242_3_lut_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i19242_3_lut_LC_5_8_1 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \RTD.i19242_3_lut_LC_5_8_1  (
            .in0(N__26565),
            .in1(N__20551),
            .in2(_gnd_net_),
            .in3(N__20578),
            .lcout(),
            .ltout(\RTD.n21362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_5_8_2 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_5_8_2 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_5_8_2  (
            .in0(N__26766),
            .in1(N__19842),
            .in2(N__19854),
            .in3(N__26189),
            .lcout(\RTD.n17835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i7_LC_5_8_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i7_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i7_LC_5_8_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i7_LC_5_8_3  (
            .in0(N__21684),
            .in1(N__21039),
            .in2(N__50177),
            .in3(N__26767),
            .lcout(buf_readRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30507),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4933_2_lut_LC_5_8_4 .C_ON=1'b0;
    defparam \RTD.i4933_2_lut_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i4933_2_lut_LC_5_8_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i4933_2_lut_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__26560),
            .in2(_gnd_net_),
            .in3(N__26187),
            .lcout(\RTD.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19410_4_lut_4_lut_LC_5_8_5 .C_ON=1'b0;
    defparam \RTD.i19410_4_lut_4_lut_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i19410_4_lut_4_lut_LC_5_8_5 .LUT_INIT=16'b1100101101111000;
    LogicCell40 \RTD.i19410_4_lut_4_lut_LC_5_8_5  (
            .in0(N__26188),
            .in1(N__26765),
            .in2(N__26591),
            .in3(N__26390),
            .lcout(\RTD.n11740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i4_LC_5_8_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i4_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i4_LC_5_8_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i4_LC_5_8_6  (
            .in0(N__20109),
            .in1(N__21683),
            .in2(N__22700),
            .in3(N__26761),
            .lcout(buf_readRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30507),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i3_LC_5_8_7 .C_ON=1'b0;
    defparam \RTD.adress_i3_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i3_LC_5_8_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \RTD.adress_i3_LC_5_8_7  (
            .in0(N__19816),
            .in1(N__19739),
            .in2(N__19791),
            .in3(N__19769),
            .lcout(adress_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30507),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_9_0 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_9_0 .LUT_INIT=16'b0011000101010101;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_9_0  (
            .in0(N__26234),
            .in1(N__26820),
            .in2(N__20076),
            .in3(N__19896),
            .lcout(\RTD.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_38_LC_5_9_1 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_38_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_38_LC_5_9_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \RTD.i1_2_lut_adj_38_LC_5_9_1  (
            .in0(N__20043),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19995),
            .lcout(\RTD.n16638 ),
            .ltout(\RTD.n16638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_adj_24_LC_5_9_2 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_adj_24_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_adj_24_LC_5_9_2 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \RTD.i2_3_lut_adj_24_LC_5_9_2  (
            .in0(N__26233),
            .in1(_gnd_net_),
            .in2(N__19950),
            .in3(N__19937),
            .lcout(\RTD.n11726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i0_LC_5_9_3 .C_ON=1'b0;
    defparam \RTD.adc_state_i0_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i0_LC_5_9_3 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \RTD.adc_state_i0_LC_5_9_3  (
            .in0(N__19926),
            .in1(N__26434),
            .in2(_gnd_net_),
            .in3(N__19920),
            .lcout(\RTD.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30468),
            .ce(N__19907),
            .sr(_gnd_net_));
    defparam \RTD.i17182_3_lut_LC_5_9_4 .C_ON=1'b0;
    defparam \RTD.i17182_3_lut_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i17182_3_lut_LC_5_9_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \RTD.i17182_3_lut_LC_5_9_4  (
            .in0(N__20545),
            .in1(N__26590),
            .in2(_gnd_net_),
            .in3(N__20574),
            .lcout(\RTD.n19787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i31_3_lut_3_lut_LC_5_9_5 .C_ON=1'b0;
    defparam \RTD.i31_3_lut_3_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i31_3_lut_3_lut_LC_5_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RTD.i31_3_lut_3_lut_LC_5_9_5  (
            .in0(N__26589),
            .in1(N__26431),
            .in2(_gnd_net_),
            .in3(N__26232),
            .lcout(),
            .ltout(\RTD.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i30_4_lut_LC_5_9_6 .C_ON=1'b0;
    defparam \RTD.i30_4_lut_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i30_4_lut_LC_5_9_6 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \RTD.i30_4_lut_LC_5_9_6  (
            .in0(N__26432),
            .in1(N__26819),
            .in2(N__19890),
            .in3(N__19887),
            .lcout(\RTD.n11704 ),
            .ltout(\RTD.n11704_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12586_2_lut_LC_5_9_7 .C_ON=1'b0;
    defparam \RTD.i12586_2_lut_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i12586_2_lut_LC_5_9_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \RTD.i12586_2_lut_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19869),
            .in3(N__26433),
            .lcout(\RTD.n14999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_tmp_i1_LC_5_10_0 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i1_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i1_LC_5_10_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i1_LC_5_10_0  (
            .in0(N__26199),
            .in1(N__20133),
            .in2(N__21178),
            .in3(N__26847),
            .lcout(\RTD.cfg_tmp_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.cfg_tmp_i2_LC_5_10_1 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i2_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i2_LC_5_10_1 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.cfg_tmp_i2_LC_5_10_1  (
            .in0(N__26843),
            .in1(N__20190),
            .in2(N__21877),
            .in3(N__26206),
            .lcout(\RTD.cfg_tmp_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.cfg_tmp_i3_LC_5_10_2 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i3_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i3_LC_5_10_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i3_LC_5_10_2  (
            .in0(N__26200),
            .in1(N__20184),
            .in2(N__24696),
            .in3(N__26848),
            .lcout(\RTD.cfg_tmp_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.cfg_tmp_i4_LC_5_10_3 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i4_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i4_LC_5_10_3 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i4_LC_5_10_3  (
            .in0(N__26844),
            .in1(N__26204),
            .in2(N__22781),
            .in3(N__20178),
            .lcout(\RTD.cfg_tmp_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.cfg_tmp_i5_LC_5_10_4 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i5_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i5_LC_5_10_4 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \RTD.cfg_tmp_i5_LC_5_10_4  (
            .in0(N__26201),
            .in1(N__26846),
            .in2(N__21811),
            .in3(N__20172),
            .lcout(\RTD.cfg_tmp_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.cfg_tmp_i6_LC_5_10_5 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i6_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i6_LC_5_10_5 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i6_LC_5_10_5  (
            .in0(N__26845),
            .in1(N__26205),
            .in2(N__31385),
            .in3(N__20166),
            .lcout(\RTD.cfg_tmp_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.cfg_tmp_i7_LC_5_10_6 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i7_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i7_LC_5_10_6 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i7_LC_5_10_6  (
            .in0(N__26202),
            .in1(N__20160),
            .in2(N__31302),
            .in3(N__26849),
            .lcout(\RTD.cfg_tmp_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.cfg_tmp_i0_LC_5_10_7 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i0_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i0_LC_5_10_7 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i0_LC_5_10_7  (
            .in0(N__26842),
            .in1(N__26203),
            .in2(N__23257),
            .in3(N__20144),
            .lcout(\RTD.cfg_tmp_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30492),
            .ce(N__20127),
            .sr(N__20118));
    defparam \RTD.read_buf_i5_LC_5_11_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i5_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i5_LC_5_11_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.read_buf_i5_LC_5_11_0  (
            .in0(N__20893),
            .in1(N__20105),
            .in2(N__20229),
            .in3(N__20985),
            .lcout(read_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30506),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i0_LC_5_11_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i0_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i0_LC_5_11_1 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i0_LC_5_11_1  (
            .in0(N__26838),
            .in1(N__20273),
            .in2(N__43439),
            .in3(N__21701),
            .lcout(buf_readRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30506),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i1_LC_5_11_2 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i1_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i1_LC_5_11_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i1_LC_5_11_2  (
            .in0(N__21703),
            .in1(N__20245),
            .in2(N__37193),
            .in3(N__26840),
            .lcout(buf_readRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30506),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i1_LC_5_11_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i1_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i1_LC_5_11_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i1_LC_5_11_3  (
            .in0(N__20274),
            .in1(N__20984),
            .in2(N__20249),
            .in3(N__20895),
            .lcout(read_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30506),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i6_LC_5_11_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i6_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i6_LC_5_11_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i6_LC_5_11_4  (
            .in0(N__21704),
            .in1(N__20207),
            .in2(N__46304),
            .in3(N__26841),
            .lcout(buf_readRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30506),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i12_LC_5_11_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i12_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i12_LC_5_11_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i12_LC_5_11_6  (
            .in0(N__21702),
            .in1(N__20383),
            .in2(N__22727),
            .in3(N__26839),
            .lcout(buf_readRTD_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30506),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i12_LC_5_11_7 .C_ON=1'b0;
    defparam \RTD.read_buf_i12_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i12_LC_5_11_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i12_LC_5_11_7  (
            .in0(N__20801),
            .in1(N__20983),
            .in2(N__20385),
            .in3(N__20894),
            .lcout(read_buf_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30506),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i14_LC_5_12_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i14_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i14_LC_5_12_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.read_buf_i14_LC_5_12_1  (
            .in0(N__20896),
            .in1(N__20779),
            .in2(N__20366),
            .in3(N__20992),
            .lcout(read_buf_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30494),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i7_LC_5_12_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i7_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i7_LC_5_12_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \RTD.read_buf_i7_LC_5_12_2  (
            .in0(N__20206),
            .in1(N__20988),
            .in2(N__20911),
            .in3(N__21031),
            .lcout(read_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30494),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i5_LC_5_12_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i5_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i5_LC_5_12_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i5_LC_5_12_3  (
            .in0(N__20227),
            .in1(N__21710),
            .in2(N__51194),
            .in3(N__26833),
            .lcout(buf_readRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30494),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i6_LC_5_12_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i6_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i6_LC_5_12_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i6_LC_5_12_4  (
            .in0(N__20228),
            .in1(N__20987),
            .in2(N__20208),
            .in3(N__20899),
            .lcout(read_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30494),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i15_LC_5_12_5 .C_ON=1'b0;
    defparam \RTD.read_buf_i15_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i15_LC_5_12_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i15_LC_5_12_5  (
            .in0(N__20897),
            .in1(N__20660),
            .in2(N__20367),
            .in3(N__20993),
            .lcout(read_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30494),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i13_LC_5_12_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i13_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i13_LC_5_12_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i13_LC_5_12_6  (
            .in0(N__20384),
            .in1(N__20986),
            .in2(N__20781),
            .in3(N__20898),
            .lcout(read_buf_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30494),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i14_LC_5_12_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i14_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i14_LC_5_12_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i14_LC_5_12_7  (
            .in0(N__20362),
            .in1(N__21709),
            .in2(N__31403),
            .in3(N__26832),
            .lcout(buf_readRTD_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30494),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_0  (
            .in0(N__20327),
            .in1(N__33387),
            .in2(N__20349),
            .in3(N__31619),
            .lcout(cmd_rdadctmp_0_adj_1450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54408),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19764_LC_5_13_4.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19764_LC_5_13_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19764_LC_5_13_4.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19764_LC_5_13_4 (
            .in0(N__21793),
            .in1(N__55158),
            .in2(N__20763),
            .in3(N__57738),
            .lcout(n22405),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i5_LC_5_14_2.C_ON=1'b0;
    defparam buf_control_i5_LC_5_14_2.SEQ_MODE=4'b1000;
    defparam buf_control_i5_LC_5_14_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i5_LC_5_14_2 (
            .in0(N__56554),
            .in1(N__41891),
            .in2(N__43600),
            .in3(N__23047),
            .lcout(AMPV_POW),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54418),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_5_15_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_5_15_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i1_LC_5_15_5  (
            .in0(N__20331),
            .in1(N__33389),
            .in2(N__20316),
            .in3(N__31562),
            .lcout(cmd_rdadctmp_1_adj_1449),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54427),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_5_15_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_5_15_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i2_LC_5_15_7  (
            .in0(N__20315),
            .in1(N__33390),
            .in2(N__21068),
            .in3(N__31563),
            .lcout(cmd_rdadctmp_2_adj_1448),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54427),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.CS_28_LC_6_3_3 .C_ON=1'b0;
    defparam \CLK_DDS.CS_28_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.CS_28_LC_6_3_3 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \CLK_DDS.CS_28_LC_6_3_3  (
            .in0(N__34796),
            .in1(N__34567),
            .in2(_gnd_net_),
            .in3(N__34459),
            .lcout(DDS_CS1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54275),
            .ce(N__20286),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i23_4_lut_LC_6_4_1 .C_ON=1'b0;
    defparam \CLK_DDS.i23_4_lut_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i23_4_lut_LC_6_4_1 .LUT_INIT=16'b1100110110011001;
    LogicCell40 \CLK_DDS.i23_4_lut_LC_6_4_1  (
            .in0(N__34710),
            .in1(N__34548),
            .in2(N__44073),
            .in3(N__34458),
            .lcout(\CLK_DDS.n9_adj_1394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i5_LC_6_6_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i5_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i5_LC_6_6_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i5_LC_6_6_0  (
            .in0(N__35797),
            .in1(N__35625),
            .in2(N__20607),
            .in3(N__20456),
            .lcout(buf_adcdata_iac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54292),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i5_LC_6_6_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i5_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i5_LC_6_6_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i5_LC_6_6_2  (
            .in0(N__20477),
            .in1(N__33681),
            .in2(N__21612),
            .in3(N__33475),
            .lcout(buf_adcdata_vac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54292),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i19_3_lut_LC_6_6_3.C_ON=1'b0;
    defparam mux_130_Mux_5_i19_3_lut_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i19_3_lut_LC_6_6_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_5_i19_3_lut_LC_6_6_3 (
            .in0(N__21264),
            .in1(N__20476),
            .in2(_gnd_net_),
            .in3(N__57815),
            .lcout(),
            .ltout(n19_adj_1629_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i22_3_lut_LC_6_6_4.C_ON=1'b0;
    defparam mux_130_Mux_5_i22_3_lut_LC_6_6_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i22_3_lut_LC_6_6_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_5_i22_3_lut_LC_6_6_4 (
            .in0(_gnd_net_),
            .in1(N__20455),
            .in2(N__20442),
            .in3(N__53797),
            .lcout(n22_adj_1630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i6_LC_6_6_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i6_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i6_LC_6_6_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i6_LC_6_6_5  (
            .in0(N__35624),
            .in1(N__35798),
            .in2(N__21095),
            .in3(N__20648),
            .lcout(buf_adcdata_iac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54292),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i30_3_lut_LC_6_6_7.C_ON=1'b0;
    defparam mux_130_Mux_6_i30_3_lut_LC_6_6_7.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i30_3_lut_LC_6_6_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_6_i30_3_lut_LC_6_6_7 (
            .in0(N__20439),
            .in1(N__20628),
            .in2(_gnd_net_),
            .in3(N__54765),
            .lcout(n30_adj_1628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i19_3_lut_LC_6_7_0.C_ON=1'b0;
    defparam mux_130_Mux_4_i19_3_lut_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i19_3_lut_LC_6_7_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_4_i19_3_lut_LC_6_7_0 (
            .in0(N__24081),
            .in1(N__20425),
            .in2(_gnd_net_),
            .in3(N__57816),
            .lcout(),
            .ltout(n19_adj_1632_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i22_3_lut_LC_6_7_1.C_ON=1'b0;
    defparam mux_130_Mux_4_i22_3_lut_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i22_3_lut_LC_6_7_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_4_i22_3_lut_LC_6_7_1 (
            .in0(_gnd_net_),
            .in1(N__20398),
            .in2(N__20409),
            .in3(N__53799),
            .lcout(n22_adj_1633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i4_LC_6_7_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i4_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i4_LC_6_7_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i4_LC_6_7_3  (
            .in0(N__35802),
            .in1(N__35632),
            .in2(N__20622),
            .in3(N__20399),
            .lcout(buf_adcdata_iac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54301),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i22_3_lut_LC_6_7_4.C_ON=1'b0;
    defparam mux_130_Mux_6_i22_3_lut_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i22_3_lut_LC_6_7_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_130_Mux_6_i22_3_lut_LC_6_7_4 (
            .in0(N__53798),
            .in1(N__20644),
            .in2(_gnd_net_),
            .in3(N__21357),
            .lcout(n22_adj_1627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_6_7_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_6_7_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i12_LC_6_7_5  (
            .in0(N__20617),
            .in1(N__28103),
            .in2(N__28398),
            .in3(N__35633),
            .lcout(cmd_rdadctmp_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_6_7_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_6_7_6 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i13_LC_6_7_6  (
            .in0(N__35631),
            .in1(N__20618),
            .in2(N__28123),
            .in3(N__20599),
            .lcout(cmd_rdadctmp_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_6_7_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_6_7_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i14_LC_6_7_7  (
            .in0(N__21085),
            .in1(N__28104),
            .in2(N__20606),
            .in3(N__35634),
            .lcout(cmd_rdadctmp_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54301),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i10_LC_6_8_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i10_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i10_LC_6_8_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i10_LC_6_8_1  (
            .in0(N__20820),
            .in1(N__21708),
            .in2(N__21011),
            .in3(N__26831),
            .lcout(buf_readRTD_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30476),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i1_3_lut_LC_6_8_2 .C_ON=1'b0;
    defparam \CLK_DDS.i1_3_lut_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i1_3_lut_LC_6_8_2 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \CLK_DDS.i1_3_lut_LC_6_8_2  (
            .in0(N__34711),
            .in1(N__34536),
            .in2(_gnd_net_),
            .in3(N__34425),
            .lcout(\CLK_DDS.n16894 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_LC_6_8_6 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_LC_6_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \RTD.i2_3_lut_LC_6_8_6  (
            .in0(N__20699),
            .in1(N__20514),
            .in2(_gnd_net_),
            .in3(N__20497),
            .lcout(\RTD.n17799 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.bit_cnt_3771__i3_LC_6_9_0 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i3_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i3_LC_6_9_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \RTD.bit_cnt_3771__i3_LC_6_9_0  (
            .in0(N__20517),
            .in1(N__20544),
            .in2(N__20709),
            .in3(N__20499),
            .lcout(\RTD.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30449),
            .ce(N__20682),
            .sr(N__26088));
    defparam \RTD.bit_cnt_3771__i1_LC_6_9_1 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i1_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i1_LC_6_9_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RTD.bit_cnt_3771__i1_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__20701),
            .in2(_gnd_net_),
            .in3(N__20515),
            .lcout(\RTD.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30449),
            .ce(N__20682),
            .sr(N__26088));
    defparam \RTD.bit_cnt_3771__i2_LC_6_9_2 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i2_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i2_LC_6_9_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \RTD.bit_cnt_3771__i2_LC_6_9_2  (
            .in0(N__20516),
            .in1(_gnd_net_),
            .in2(N__20708),
            .in3(N__20498),
            .lcout(\RTD.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30449),
            .ce(N__20682),
            .sr(N__26088));
    defparam \RTD.bit_cnt_3771__i0_LC_6_9_3 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i0_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i0_LC_6_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \RTD.bit_cnt_3771__i0_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20700),
            .lcout(\RTD.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30449),
            .ce(N__20682),
            .sr(N__26088));
    defparam i15340_2_lut_3_lut_LC_6_9_6.C_ON=1'b0;
    defparam i15340_2_lut_3_lut_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam i15340_2_lut_3_lut_LC_6_9_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15340_2_lut_3_lut_LC_6_9_6 (
            .in0(N__40120),
            .in1(N__51726),
            .in2(_gnd_net_),
            .in3(N__55516),
            .lcout(n14_adj_1580),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15341_2_lut_3_lut_LC_6_9_7.C_ON=1'b0;
    defparam i15341_2_lut_3_lut_LC_6_9_7.SEQ_MODE=4'b0000;
    defparam i15341_2_lut_3_lut_LC_6_9_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15341_2_lut_3_lut_LC_6_9_7 (
            .in0(N__55517),
            .in1(N__50319),
            .in2(_gnd_net_),
            .in3(N__51727),
            .lcout(n14_adj_1551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i3_LC_6_10_0 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i3_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i3_LC_6_10_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \CLK_DDS.bit_cnt_i3_LC_6_10_0  (
            .in0(N__24777),
            .in1(N__21422),
            .in2(N__21402),
            .in3(N__21441),
            .lcout(bit_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54340),
            .ce(N__34751),
            .sr(N__20670));
    defparam \CLK_DDS.bit_cnt_i2_LC_6_10_1 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i2_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i2_LC_6_10_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \CLK_DDS.bit_cnt_i2_LC_6_10_1  (
            .in0(N__21421),
            .in1(N__21398),
            .in2(_gnd_net_),
            .in3(N__24776),
            .lcout(bit_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54340),
            .ce(N__34751),
            .sr(N__20670));
    defparam \CLK_DDS.bit_cnt_i1_LC_6_10_2 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i1_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i1_LC_6_10_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \CLK_DDS.bit_cnt_i1_LC_6_10_2  (
            .in0(N__24775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21420),
            .lcout(bit_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54340),
            .ce(N__34751),
            .sr(N__20670));
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_11_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_11_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i27_LC_6_11_1  (
            .in0(N__33450),
            .in1(N__24485),
            .in2(N__22637),
            .in3(N__31592),
            .lcout(cmd_rdadctmp_27_adj_1423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54354),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i11_LC_6_12_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i11_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i11_LC_6_12_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i11_LC_6_12_0  (
            .in0(N__20816),
            .in1(N__20990),
            .in2(N__20802),
            .in3(N__20904),
            .lcout(read_buf_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30493),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i15_LC_6_12_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i15_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i15_LC_6_12_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i15_LC_6_12_1  (
            .in0(N__20661),
            .in1(N__21712),
            .in2(N__31319),
            .in3(N__26835),
            .lcout(buf_readRTD_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30493),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i8_LC_6_12_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i8_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i8_LC_6_12_2 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \RTD.read_buf_i8_LC_6_12_2  (
            .in0(N__21733),
            .in1(N__20991),
            .in2(N__20913),
            .in3(N__21032),
            .lcout(read_buf_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30493),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i9_LC_6_12_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i9_LC_6_12_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i9_LC_6_12_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.read_buf_i9_LC_6_12_3  (
            .in0(N__20903),
            .in1(N__21734),
            .in2(N__20744),
            .in3(N__20994),
            .lcout(read_buf_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30493),
            .ce(),
            .sr(_gnd_net_));
    defparam i18472_3_lut_LC_6_12_5.C_ON=1'b0;
    defparam i18472_3_lut_LC_6_12_5.SEQ_MODE=4'b0000;
    defparam i18472_3_lut_LC_6_12_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18472_3_lut_LC_6_12_5 (
            .in0(N__21015),
            .in1(N__21843),
            .in2(_gnd_net_),
            .in3(N__57784),
            .lcout(n21082),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i10_LC_6_12_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i10_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i10_LC_6_12_6 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \RTD.read_buf_i10_LC_6_12_6  (
            .in0(N__20815),
            .in1(N__20989),
            .in2(N__20912),
            .in3(N__20740),
            .lcout(read_buf_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30493),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i11_LC_6_12_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i11_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i11_LC_6_12_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i11_LC_6_12_7  (
            .in0(N__20800),
            .in1(N__21711),
            .in2(N__24629),
            .in3(N__26834),
            .lcout(buf_readRTD_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30493),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i13_LC_6_13_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i13_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i13_LC_6_13_0 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i13_LC_6_13_0  (
            .in0(N__26851),
            .in1(N__20780),
            .in2(N__20762),
            .in3(N__21719),
            .lcout(buf_readRTD_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30459),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_LC_6_13_3.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_LC_6_13_3.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_LC_6_13_3 (
            .in0(N__21150),
            .in1(N__55159),
            .in2(N__20724),
            .in3(N__57740),
            .lcout(n22441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i9_LC_6_13_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i9_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i9_LC_6_13_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \RTD.READ_DATA_i9_LC_6_13_5  (
            .in0(N__21720),
            .in1(N__20720),
            .in2(N__20745),
            .in3(N__26852),
            .lcout(buf_readRTD_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30459),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_6_14_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_6_14_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i23_LC_6_14_0  (
            .in0(N__35535),
            .in1(N__22891),
            .in2(N__25127),
            .in3(N__28046),
            .lcout(cmd_rdadctmp_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54394),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_6_14_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_6_14_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i22_LC_6_14_1  (
            .in0(N__28045),
            .in1(N__35240),
            .in2(N__22895),
            .in3(N__35538),
            .lcout(cmd_rdadctmp_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54394),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i10_LC_6_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i10_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i10_LC_6_14_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i10_LC_6_14_3  (
            .in0(N__35742),
            .in1(N__35537),
            .in2(N__23346),
            .in3(N__46633),
            .lcout(buf_adcdata_iac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54394),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i1_LC_6_14_4.C_ON=1'b0;
    defparam buf_cfgRTD_i1_LC_6_14_4.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i1_LC_6_14_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i1_LC_6_14_4 (
            .in0(N__56555),
            .in1(N__27300),
            .in2(N__40161),
            .in3(N__21151),
            .lcout(buf_cfgRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54394),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_6  (
            .in0(N__35536),
            .in1(N__21299),
            .in2(N__22655),
            .in3(N__28047),
            .lcout(cmd_rdadctmp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54394),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_0  (
            .in0(N__31560),
            .in1(N__21050),
            .in2(N__21245),
            .in3(N__33273),
            .lcout(cmd_rdadctmp_4_adj_1446),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54409),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_6_15_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_6_15_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i16_LC_6_15_1  (
            .in0(N__35558),
            .in1(N__23143),
            .in2(N__28065),
            .in3(N__22946),
            .lcout(cmd_rdadctmp_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54409),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_192_LC_6_15_2.C_ON=1'b0;
    defparam i1_4_lut_adj_192_LC_6_15_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_192_LC_6_15_2.LUT_INIT=16'b0000111100000110;
    LogicCell40 i1_4_lut_adj_192_LC_6_15_2 (
            .in0(N__33264),
            .in1(N__30707),
            .in2(N__21116),
            .in3(N__27438),
            .lcout(),
            .ltout(n14_adj_1610_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.CS_37_LC_6_15_3 .C_ON=1'b0;
    defparam \ADC_VAC.CS_37_LC_6_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.CS_37_LC_6_15_3 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \ADC_VAC.CS_37_LC_6_15_3  (
            .in0(N__23099),
            .in1(N__21231),
            .in2(N__21129),
            .in3(N__33266),
            .lcout(VAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54409),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_6_15_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_6_15_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i15_LC_6_15_4  (
            .in0(N__22945),
            .in1(N__28005),
            .in2(N__21099),
            .in3(N__35559),
            .lcout(cmd_rdadctmp_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54409),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_6_15_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_6_15_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i3_LC_6_15_5  (
            .in0(N__21069),
            .in1(N__33265),
            .in2(N__21051),
            .in3(N__31559),
            .lcout(cmd_rdadctmp_3_adj_1447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54409),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_6  (
            .in0(N__31561),
            .in1(N__21926),
            .in2(N__21246),
            .in3(N__33274),
            .lcout(cmd_rdadctmp_5_adj_1445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54409),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i2_LC_6_16_1 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i2_LC_6_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i2_LC_6_16_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_VAC.adc_state_i2_LC_6_16_1  (
            .in0(N__33221),
            .in1(N__30702),
            .in2(_gnd_net_),
            .in3(N__27431),
            .lcout(DTRIG_N_918_adj_1451),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54419),
            .ce(N__21219),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i1_LC_6_16_3 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i1_LC_6_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i1_LC_6_16_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \ADC_VAC.adc_state_i1_LC_6_16_3  (
            .in0(N__33220),
            .in1(N__30701),
            .in2(_gnd_net_),
            .in3(N__27432),
            .lcout(adc_state_1_adj_1417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54419),
            .ce(N__21219),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_203_LC_6_16_5.C_ON=1'b0;
    defparam i1_2_lut_adj_203_LC_6_16_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_203_LC_6_16_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_203_LC_6_16_5 (
            .in0(_gnd_net_),
            .in1(N__30700),
            .in2(_gnd_net_),
            .in3(N__27430),
            .lcout(n20864),
            .ltout(n20864_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_3_lut_LC_6_16_6 .C_ON=1'b0;
    defparam \ADC_VAC.i1_3_lut_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_3_lut_LC_6_16_6 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \ADC_VAC.i1_3_lut_LC_6_16_6  (
            .in0(_gnd_net_),
            .in1(N__23100),
            .in2(N__21225),
            .in3(N__33219),
            .lcout(n12653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i30_4_lut_LC_6_17_2 .C_ON=1'b0;
    defparam \ADC_VAC.i30_4_lut_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i30_4_lut_LC_6_17_2 .LUT_INIT=16'b1110000001000101;
    LogicCell40 \ADC_VAC.i30_4_lut_LC_6_17_2  (
            .in0(N__30706),
            .in1(N__23101),
            .in2(N__27448),
            .in3(N__25404),
            .lcout(),
            .ltout(\ADC_VAC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19365_2_lut_LC_6_17_3 .C_ON=1'b0;
    defparam \ADC_VAC.i19365_2_lut_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19365_2_lut_LC_6_17_3 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \ADC_VAC.i19365_2_lut_LC_6_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21222),
            .in3(N__33259),
            .lcout(\ADC_VAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.CS_37_LC_6_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.CS_37_LC_6_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.CS_37_LC_6_18_0 .LUT_INIT=16'b0011001000110011;
    LogicCell40 \ADC_IAC.CS_37_LC_6_18_0  (
            .in0(N__35408),
            .in1(N__21186),
            .in2(N__25936),
            .in3(N__21351),
            .lcout(IAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54431),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_195_LC_6_18_1.C_ON=1'b0;
    defparam i1_4_lut_adj_195_LC_6_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_195_LC_6_18_1.LUT_INIT=16'b0000101100001110;
    LogicCell40 i1_4_lut_adj_195_LC_6_18_1 (
            .in0(N__29883),
            .in1(N__29973),
            .in2(N__21203),
            .in3(N__35407),
            .lcout(n14_adj_1612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_199_LC_6_18_2.C_ON=1'b0;
    defparam i1_2_lut_adj_199_LC_6_18_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_199_LC_6_18_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_199_LC_6_18_2 (
            .in0(_gnd_net_),
            .in1(N__29959),
            .in2(_gnd_net_),
            .in3(N__29882),
            .lcout(n20867),
            .ltout(n20867_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_3_lut_LC_6_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.i1_3_lut_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_3_lut_LC_6_18_3 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \ADC_IAC.i1_3_lut_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(N__25929),
            .in2(N__21345),
            .in3(N__35406),
            .lcout(n12498),
            .ltout(n12498_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_4  (
            .in0(N__35409),
            .in1(N__21342),
            .in2(N__21324),
            .in3(N__21320),
            .lcout(cmd_rdadctmp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54431),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_6_18_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_6_18_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_6_18_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i1_LC_6_18_6  (
            .in0(N__35410),
            .in1(N__21321),
            .in2(N__21312),
            .in3(N__28035),
            .lcout(cmd_rdadctmp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54431),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_6_18_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_6_18_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_6_18_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i2_LC_6_18_7  (
            .in0(N__28034),
            .in1(N__35411),
            .in2(N__21300),
            .in3(N__21311),
            .lcout(cmd_rdadctmp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54431),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_I_0_1_lut_LC_6_19_7.C_ON=1'b0;
    defparam acadc_rst_I_0_1_lut_LC_6_19_7.SEQ_MODE=4'b0000;
    defparam acadc_rst_I_0_1_lut_LC_6_19_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 acadc_rst_I_0_1_lut_LC_6_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40898),
            .lcout(AC_ADC_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i5_LC_7_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i5_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i5_LC_7_5_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i5_LC_7_5_4  (
            .in0(N__25701),
            .in1(N__48843),
            .in2(N__21263),
            .in3(N__22236),
            .lcout(buf_adcdata_vdc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53254),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i1_LC_7_6_0 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i1_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i1_LC_7_6_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLK_DDS.dds_state_i1_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__34547),
            .in2(_gnd_net_),
            .in3(N__34453),
            .lcout(dds_state_1_adj_1453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54287),
            .ce(N__21377),
            .sr(N__34772));
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_7_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_7_7_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i11_LC_7_7_0  (
            .in0(N__23988),
            .in1(N__22267),
            .in2(N__23888),
            .in3(N__48586),
            .lcout(cmd_rdadctmp_11_adj_1468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_1 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_1  (
            .in0(N__48583),
            .in1(N__24038),
            .in2(N__23630),
            .in3(N__23861),
            .lcout(cmd_rdadctmp_14_adj_1465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_7_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_7_7_2 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i22_LC_7_7_2  (
            .in0(N__22321),
            .in1(N__26047),
            .in2(N__23891),
            .in3(N__48589),
            .lcout(cmd_rdadctmp_22_adj_1457),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3  (
            .in0(N__48585),
            .in1(N__22322),
            .in2(N__22350),
            .in3(N__23869),
            .lcout(cmd_rdadctmp_21_adj_1458),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_4  (
            .in0(N__22345),
            .in1(N__23739),
            .in2(N__23890),
            .in3(N__48588),
            .lcout(cmd_rdadctmp_20_adj_1459),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_7_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_7_7_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i12_LC_7_7_5  (
            .in0(N__48582),
            .in1(N__23860),
            .in2(N__22272),
            .in3(N__24061),
            .lcout(cmd_rdadctmp_12_adj_1467),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_7_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_7_7_6 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i18_LC_7_7_6  (
            .in0(N__22376),
            .in1(N__23761),
            .in2(N__23889),
            .in3(N__48587),
            .lcout(cmd_rdadctmp_18_adj_1461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_7_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_7_7_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i17_LC_7_7_7  (
            .in0(N__48584),
            .in1(N__22375),
            .in2(N__23925),
            .in3(N__23862),
            .lcout(cmd_rdadctmp_17_adj_1462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53277),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i19_3_lut_LC_7_8_1.C_ON=1'b0;
    defparam mux_130_Mux_6_i19_3_lut_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i19_3_lut_LC_7_8_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_6_i19_3_lut_LC_7_8_1 (
            .in0(N__24339),
            .in1(N__21538),
            .in2(_gnd_net_),
            .in3(N__57747),
            .lcout(n19_adj_1626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_7_8_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_7_8_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i13_LC_7_8_2  (
            .in0(N__33490),
            .in1(N__21592),
            .in2(N__28292),
            .in3(N__31683),
            .lcout(cmd_rdadctmp_13_adj_1437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i7_LC_7_8_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i7_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i7_LC_7_8_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i7_LC_7_8_3  (
            .in0(N__33650),
            .in1(N__33492),
            .in2(N__21498),
            .in3(N__24292),
            .lcout(buf_adcdata_vac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_8_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_8_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i16_LC_7_8_4  (
            .in0(N__33491),
            .in1(N__21494),
            .in2(N__21473),
            .in3(N__31684),
            .lcout(cmd_rdadctmp_16_adj_1434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_8_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_8_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i17_LC_7_8_5  (
            .in0(N__31685),
            .in1(N__21469),
            .in2(N__31711),
            .in3(N__33493),
            .lcout(cmd_rdadctmp_17_adj_1433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i8_LC_7_8_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i8_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i8_LC_7_8_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i8_LC_7_8_6  (
            .in0(N__33489),
            .in1(N__33651),
            .in2(N__21474),
            .in3(N__21568),
            .lcout(buf_adcdata_vac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54302),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i30_3_lut_LC_7_8_7.C_ON=1'b0;
    defparam mux_130_Mux_4_i30_3_lut_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i30_3_lut_LC_7_8_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_4_i30_3_lut_LC_7_8_7 (
            .in0(N__21456),
            .in1(N__21447),
            .in2(_gnd_net_),
            .in3(N__54753),
            .lcout(n30_adj_1634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i0_LC_7_9_0 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i0_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i0_LC_7_9_0 .LUT_INIT=16'b1100010100000101;
    LogicCell40 \CLK_DDS.dds_state_i0_LC_7_9_0  (
            .in0(N__34437),
            .in1(N__21384),
            .in2(N__34752),
            .in3(N__21429),
            .lcout(dds_state_0_adj_1454),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54315),
            .ce(N__21378),
            .sr(_gnd_net_));
    defparam SecClk_292_LC_7_10_0.C_ON=1'b0;
    defparam SecClk_292_LC_7_10_0.SEQ_MODE=4'b1000;
    defparam SecClk_292_LC_7_10_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 SecClk_292_LC_7_10_0 (
            .in0(_gnd_net_),
            .in1(N__39168),
            .in2(_gnd_net_),
            .in3(N__31137),
            .lcout(TEST_LED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38751),
            .ce(),
            .sr(_gnd_net_));
    defparam i18974_2_lut_LC_7_10_2.C_ON=1'b0;
    defparam i18974_2_lut_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam i18974_2_lut_LC_7_10_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 i18974_2_lut_LC_7_10_2 (
            .in0(_gnd_net_),
            .in1(N__24774),
            .in2(_gnd_net_),
            .in3(N__21440),
            .lcout(n21456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_7_10_3 .C_ON=1'b0;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_7_10_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \CLK_DDS.i3_3_lut_4_lut_LC_7_10_3  (
            .in0(N__34595),
            .in1(N__34423),
            .in2(N__21423),
            .in3(N__21397),
            .lcout(n8_adj_1602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i19392_4_lut_LC_7_10_5 .C_ON=1'b0;
    defparam \CLK_DDS.i19392_4_lut_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19392_4_lut_LC_7_10_5 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \CLK_DDS.i19392_4_lut_LC_7_10_5  (
            .in0(N__34594),
            .in1(N__34424),
            .in2(N__44069),
            .in3(N__34706),
            .lcout(\CLK_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i19_LC_7_11_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i19_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i19_LC_7_11_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i19_LC_7_11_1  (
            .in0(N__33620),
            .in1(N__33307),
            .in2(N__25282),
            .in3(N__22636),
            .lcout(buf_adcdata_vac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54341),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_7_11_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_7_11_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i29_LC_7_11_2  (
            .in0(N__31670),
            .in1(N__22585),
            .in2(N__33375),
            .in3(N__22613),
            .lcout(cmd_rdadctmp_29_adj_1421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54341),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_7_11_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_7_11_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i14_LC_7_11_3  (
            .in0(N__21508),
            .in1(N__33308),
            .in2(N__21611),
            .in3(N__31668),
            .lcout(cmd_rdadctmp_14_adj_1436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54341),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_0_i19_3_lut_LC_7_11_4.C_ON=1'b0;
    defparam mux_129_Mux_0_i19_3_lut_LC_7_11_4.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i19_3_lut_LC_7_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_0_i19_3_lut_LC_7_11_4 (
            .in0(N__23679),
            .in1(N__21569),
            .in2(_gnd_net_),
            .in3(N__57572),
            .lcout(n19_adj_1486),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i6_LC_7_11_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i6_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i6_LC_7_11_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i6_LC_7_11_6  (
            .in0(N__33306),
            .in1(N__33621),
            .in2(N__21542),
            .in3(N__21512),
            .lcout(buf_adcdata_vac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54341),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_7  (
            .in0(N__21485),
            .in1(N__33309),
            .in2(N__21513),
            .in3(N__31669),
            .lcout(cmd_rdadctmp_15_adj_1435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54341),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i16_LC_7_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i16_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i16_LC_7_12_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i16_LC_7_12_0  (
            .in0(N__33603),
            .in1(N__33486),
            .in2(N__21764),
            .in3(N__22679),
            .lcout(buf_adcdata_vac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54355),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_7_12_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_7_12_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i23_LC_7_12_2  (
            .in0(N__24903),
            .in1(N__33487),
            .in2(N__24509),
            .in3(N__31628),
            .lcout(cmd_rdadctmp_23_adj_1427),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54355),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_7_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_7_12_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i24_LC_7_12_4  (
            .in0(N__24505),
            .in1(N__33488),
            .in2(N__21763),
            .in3(N__31629),
            .lcout(cmd_rdadctmp_24_adj_1426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54355),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_7_13_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_7_13_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i30_LC_7_13_1  (
            .in0(N__22596),
            .in1(N__33374),
            .in2(N__22857),
            .in3(N__31660),
            .lcout(cmd_rdadctmp_30_adj_1420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54367),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i3_LC_7_13_3.C_ON=1'b0;
    defparam buf_cfgRTD_i3_LC_7_13_3.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i3_LC_7_13_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i3_LC_7_13_3 (
            .in0(N__56558),
            .in1(N__27298),
            .in2(N__44229),
            .in3(N__24671),
            .lcout(buf_cfgRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54367),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i2_LC_7_13_4.C_ON=1'b0;
    defparam buf_cfgRTD_i2_LC_7_13_4.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i2_LC_7_13_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_cfgRTD_i2_LC_7_13_4 (
            .in0(N__27297),
            .in1(N__56559),
            .in2(N__44793),
            .in3(N__21844),
            .lcout(buf_cfgRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54367),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i5_LC_7_13_5.C_ON=1'b0;
    defparam buf_cfgRTD_i5_LC_7_13_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i5_LC_7_13_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i5_LC_7_13_5 (
            .in0(N__56557),
            .in1(N__27299),
            .in2(N__43605),
            .in3(N__21789),
            .lcout(buf_cfgRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54367),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_7_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_7_13_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i20_LC_7_13_6  (
            .in0(N__31994),
            .in1(N__28063),
            .in2(N__25036),
            .in3(N__35520),
            .lcout(cmd_rdadctmp_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54367),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_7_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_7_13_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i25_LC_7_13_7  (
            .in0(N__21765),
            .in1(N__33373),
            .in2(N__24416),
            .in3(N__31659),
            .lcout(cmd_rdadctmp_25_adj_1425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54367),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19694_LC_7_14_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19694_LC_7_14_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19694_LC_7_14_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19694_LC_7_14_2 (
            .in0(N__23025),
            .in1(N__54748),
            .in2(N__35196),
            .in3(N__53780),
            .lcout(),
            .ltout(n22321_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22321_bdd_4_lut_LC_7_14_3.C_ON=1'b0;
    defparam n22321_bdd_4_lut_LC_7_14_3.SEQ_MODE=4'b0000;
    defparam n22321_bdd_4_lut_LC_7_14_3.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22321_bdd_4_lut_LC_7_14_3 (
            .in0(N__54749),
            .in1(N__22788),
            .in2(N__21741),
            .in3(N__22908),
            .lcout(n22324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i8_LC_7_14_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i8_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i8_LC_7_14_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i8_LC_7_14_5  (
            .in0(N__21738),
            .in1(N__21718),
            .in2(N__23277),
            .in3(N__26856),
            .lcout(buf_readRTD_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30513),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_7_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_7_15_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i7_LC_7_15_2  (
            .in0(N__31565),
            .in1(N__21914),
            .in2(N__22562),
            .in3(N__33272),
            .lcout(cmd_rdadctmp_7_adj_1443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54395),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i15_LC_7_15_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i15_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i15_LC_7_15_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i15_LC_7_15_3  (
            .in0(N__35719),
            .in1(N__35459),
            .in2(N__52177),
            .in3(N__25126),
            .lcout(buf_adcdata_iac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54395),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.SCLK_35_LC_7_15_5 .C_ON=1'b0;
    defparam \ADC_VAC.SCLK_35_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.SCLK_35_LC_7_15_5 .LUT_INIT=16'b1111000101100000;
    LogicCell40 \ADC_VAC.SCLK_35_LC_7_15_5  (
            .in0(N__27439),
            .in1(N__33267),
            .in2(N__21947),
            .in3(N__30708),
            .lcout(VAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54395),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_7_15_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_7_15_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i6_LC_7_15_7  (
            .in0(N__21930),
            .in1(N__33268),
            .in2(N__21915),
            .in3(N__31564),
            .lcout(cmd_rdadctmp_6_adj_1444),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54395),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i0_LC_7_16_6 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i0_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i0_LC_7_16_6 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \ADC_VAC.adc_state_i0_LC_7_16_6  (
            .in0(N__30713),
            .in1(N__27440),
            .in2(N__33343),
            .in3(N__21903),
            .lcout(adc_state_0_adj_1418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54410),
            .ce(N__21894),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_7_17_0.C_ON=1'b0;
    defparam i1_2_lut_LC_7_17_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_7_17_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_LC_7_17_0 (
            .in0(_gnd_net_),
            .in1(N__29993),
            .in2(_gnd_net_),
            .in3(N__29902),
            .lcout(n20858),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i12393_2_lut_LC_7_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.i12393_2_lut_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i12393_2_lut_LC_7_17_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \ADC_IAC.i12393_2_lut_LC_7_17_1  (
            .in0(N__29994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25877),
            .lcout(\ADC_IAC.n14806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19093_4_lut_LC_7_17_4 .C_ON=1'b0;
    defparam \ADC_VAC.i19093_4_lut_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19093_4_lut_LC_7_17_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ADC_VAC.i19093_4_lut_LC_7_17_4  (
            .in0(N__33260),
            .in1(N__27434),
            .in2(N__25323),
            .in3(N__25446),
            .lcout(\ADC_VAC.n21312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_LC_7_17_5 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_LC_7_17_5 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \ADC_VAC.i1_4_lut_LC_7_17_5  (
            .in0(N__33245),
            .in1(N__23102),
            .in2(N__30720),
            .in3(N__25403),
            .lcout(),
            .ltout(\ADC_VAC.n20958_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_adj_4_LC_7_17_6 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_adj_4_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_adj_4_LC_7_17_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \ADC_VAC.i1_2_lut_adj_4_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21897),
            .in3(N__27433),
            .lcout(\ADC_VAC.n20959 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_7_18_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_7_18_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i17_LC_7_18_1  (
            .in0(N__23156),
            .in1(N__27975),
            .in2(N__23122),
            .in3(N__35405),
            .lcout(cmd_rdadctmp_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54428),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i2_LC_7_19_0 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i2_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i2_LC_7_19_0 .LUT_INIT=16'b0000111111000000;
    LogicCell40 \ADC_IAC.adc_state_i2_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__35403),
            .in2(N__29995),
            .in3(N__29901),
            .lcout(DTRIG_N_918),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54432),
            .ce(N__23505),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i1_LC_7_19_1 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i1_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i1_LC_7_19_1 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \ADC_IAC.adc_state_i1_LC_7_19_1  (
            .in0(N__29900),
            .in1(N__29974),
            .in2(_gnd_net_),
            .in3(N__35404),
            .lcout(adc_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54432),
            .ce(N__23505),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_3_lut_4_lut_4_lut_LC_8_2_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_3_lut_4_lut_4_lut_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_3_lut_4_lut_4_lut_LC_8_2_1 .LUT_INIT=16'b1101110110000000;
    LogicCell40 \ADC_VDC.i1_3_lut_3_lut_4_lut_4_lut_LC_8_2_1  (
            .in0(N__47385),
            .in1(N__48847),
            .in2(N__48357),
            .in3(N__48568),
            .lcout(\ADC_VDC.n13034 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7_4_lut_LC_8_2_2 .C_ON=1'b0;
    defparam \ADC_VDC.i7_4_lut_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7_4_lut_LC_8_2_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i7_4_lut_LC_8_2_2  (
            .in0(N__22014),
            .in1(N__21971),
            .in2(N__22035),
            .in3(N__22101),
            .lcout(),
            .ltout(\ADC_VDC.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i11_3_lut_LC_8_2_3 .C_ON=1'b0;
    defparam \ADC_VDC.i11_3_lut_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i11_3_lut_LC_8_2_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \ADC_VDC.i11_3_lut_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__23448),
            .in2(N__21996),
            .in3(N__23391),
            .lcout(\ADC_VDC.n18563 ),
            .ltout(\ADC_VDC.n18563_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16137_3_lut_LC_8_2_4 .C_ON=1'b0;
    defparam \ADC_VDC.i16137_3_lut_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16137_3_lut_LC_8_2_4 .LUT_INIT=16'b0011001111111100;
    LogicCell40 \ADC_VDC.i16137_3_lut_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(N__48350),
            .in2(N__21993),
            .in3(N__47384),
            .lcout(\ADC_VDC.n18566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19290_3_lut_LC_8_2_6 .C_ON=1'b0;
    defparam \ADC_VDC.i19290_3_lut_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19290_3_lut_LC_8_2_6 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \ADC_VDC.i19290_3_lut_LC_8_2_6  (
            .in0(N__24226),
            .in1(_gnd_net_),
            .in2(N__48871),
            .in3(N__21990),
            .lcout(),
            .ltout(\ADC_VDC.n21384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_8_2_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_8_2_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i34_LC_8_2_7  (
            .in0(N__48354),
            .in1(N__22386),
            .in2(N__21984),
            .in3(N__48569),
            .lcout(cmd_rdadcbuf_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53325),
            .ce(N__21981),
            .sr(_gnd_net_));
    defparam \ADC_VDC.avg_cnt_i0_LC_8_3_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i0_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i0_LC_8_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i0_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__21972),
            .in2(_gnd_net_),
            .in3(N__21960),
            .lcout(\ADC_VDC.avg_cnt_0 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\ADC_VDC.n19698 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i1_LC_8_3_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i1_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i1_LC_8_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i1_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__23417),
            .in2(_gnd_net_),
            .in3(N__22056),
            .lcout(\ADC_VDC.avg_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19698 ),
            .carryout(\ADC_VDC.n19699 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i2_LC_8_3_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i2_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i2_LC_8_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i2_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__23430),
            .in2(_gnd_net_),
            .in3(N__22053),
            .lcout(\ADC_VDC.avg_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19699 ),
            .carryout(\ADC_VDC.n19700 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i3_LC_8_3_3 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i3_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i3_LC_8_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i3_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__23474),
            .in2(_gnd_net_),
            .in3(N__22050),
            .lcout(\ADC_VDC.avg_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19700 ),
            .carryout(\ADC_VDC.n19701 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i4_LC_8_3_4 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i4_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i4_LC_8_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i4_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__23499),
            .in2(_gnd_net_),
            .in3(N__22047),
            .lcout(\ADC_VDC.avg_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19701 ),
            .carryout(\ADC_VDC.n19702 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i5_LC_8_3_5 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i5_LC_8_3_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i5_LC_8_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i5_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(N__23460),
            .in2(_gnd_net_),
            .in3(N__22044),
            .lcout(\ADC_VDC.avg_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19702 ),
            .carryout(\ADC_VDC.n19703 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i6_LC_8_3_6 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i6_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i6_LC_8_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i6_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(N__23403),
            .in2(_gnd_net_),
            .in3(N__22041),
            .lcout(\ADC_VDC.avg_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19703 ),
            .carryout(\ADC_VDC.n19704 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i7_LC_8_3_7 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i7_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i7_LC_8_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i7_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__23487),
            .in2(_gnd_net_),
            .in3(N__22038),
            .lcout(\ADC_VDC.avg_cnt_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19704 ),
            .carryout(\ADC_VDC.n19705 ),
            .clk(N__53319),
            .ce(N__22506),
            .sr(N__22443));
    defparam \ADC_VDC.avg_cnt_i8_LC_8_4_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i8_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i8_LC_8_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i8_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(N__22031),
            .in2(_gnd_net_),
            .in3(N__22017),
            .lcout(\ADC_VDC.avg_cnt_8 ),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\ADC_VDC.n19706 ),
            .clk(N__53320),
            .ce(N__22514),
            .sr(N__22452));
    defparam \ADC_VDC.avg_cnt_i9_LC_8_4_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i9_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i9_LC_8_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i9_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(N__22013),
            .in2(_gnd_net_),
            .in3(N__21999),
            .lcout(\ADC_VDC.avg_cnt_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19706 ),
            .carryout(\ADC_VDC.n19707 ),
            .clk(N__53320),
            .ce(N__22514),
            .sr(N__22452));
    defparam \ADC_VDC.avg_cnt_i10_LC_8_4_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i10_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i10_LC_8_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i10_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__22100),
            .in2(_gnd_net_),
            .in3(N__22086),
            .lcout(\ADC_VDC.avg_cnt_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19707 ),
            .carryout(\ADC_VDC.n19708 ),
            .clk(N__53320),
            .ce(N__22514),
            .sr(N__22452));
    defparam \ADC_VDC.avg_cnt_i11_LC_8_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.avg_cnt_i11_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i11_LC_8_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i11_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(N__23442),
            .in2(_gnd_net_),
            .in3(N__22083),
            .lcout(\ADC_VDC.avg_cnt_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53320),
            .ce(N__22514),
            .sr(N__22452));
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_0  (
            .in0(N__22184),
            .in1(N__23599),
            .in2(N__23838),
            .in3(N__48562),
            .lcout(cmd_rdadctmp_3_adj_1476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_8_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_8_5_1 .LUT_INIT=16'b1110000010101000;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_8_5_1  (
            .in0(N__48556),
            .in1(N__48347),
            .in2(N__48869),
            .in3(N__47364),
            .lcout(\ADC_VDC.n13010 ),
            .ltout(\ADC_VDC.n13010_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i12541_2_lut_LC_8_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.i12541_2_lut_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i12541_2_lut_LC_8_5_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ADC_VDC.i12541_2_lut_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22080),
            .in3(N__48557),
            .lcout(\ADC_VDC.n14915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3  (
            .in0(N__48558),
            .in1(N__48348),
            .in2(N__48870),
            .in3(N__47365),
            .lcout(n12871),
            .ltout(n12871_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_8_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_8_5_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i2_LC_8_5_4  (
            .in0(N__22183),
            .in1(N__22211),
            .in2(N__22077),
            .in3(N__48561),
            .lcout(cmd_rdadctmp_2_adj_1477),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_6 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_6  (
            .in0(N__22073),
            .in1(N__22210),
            .in2(N__23837),
            .in3(N__48560),
            .lcout(cmd_rdadctmp_1_adj_1478),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_7  (
            .in0(N__48559),
            .in1(N__23800),
            .in2(N__47426),
            .in3(N__22072),
            .lcout(cmd_rdadctmp_0_adj_1479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__22218),
            .in2(N__22074),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.cmd_rdadcbuf_0 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\ADC_VDC.n19663 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__22194),
            .in2(N__22212),
            .in3(N__22188),
            .lcout(\ADC_VDC.cmd_rdadcbuf_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19663 ),
            .carryout(\ADC_VDC.n19664 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__22167),
            .in2(N__22185),
            .in3(N__22161),
            .lcout(\ADC_VDC.cmd_rdadcbuf_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19664 ),
            .carryout(\ADC_VDC.n19665 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__22158),
            .in2(N__23601),
            .in3(N__22152),
            .lcout(\ADC_VDC.cmd_rdadcbuf_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19665 ),
            .carryout(\ADC_VDC.n19666 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__22149),
            .in2(N__23580),
            .in3(N__22143),
            .lcout(\ADC_VDC.cmd_rdadcbuf_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19666 ),
            .carryout(\ADC_VDC.n19667 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__22140),
            .in2(N__24160),
            .in3(N__22134),
            .lcout(\ADC_VDC.cmd_rdadcbuf_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19667 ),
            .carryout(\ADC_VDC.n19668 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__22131),
            .in2(N__24131),
            .in3(N__22125),
            .lcout(\ADC_VDC.cmd_rdadcbuf_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19668 ),
            .carryout(\ADC_VDC.n19669 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__24106),
            .in2(N__22122),
            .in3(N__22113),
            .lcout(\ADC_VDC.cmd_rdadcbuf_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19669 ),
            .carryout(\ADC_VDC.n19670 ),
            .clk(N__53256),
            .ce(N__22521),
            .sr(N__22453));
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__22110),
            .in2(N__23559),
            .in3(N__22104),
            .lcout(\ADC_VDC.cmd_rdadcbuf_8 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\ADC_VDC.n19671 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__22290),
            .in2(N__24011),
            .in3(N__22284),
            .lcout(\ADC_VDC.cmd_rdadcbuf_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19671 ),
            .carryout(\ADC_VDC.n19672 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__22281),
            .in2(N__23987),
            .in3(N__22275),
            .lcout(\ADC_VDC.cmd_rdadcbuf_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19672 ),
            .carryout(\ADC_VDC.n19673 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__25784),
            .in2(N__22271),
            .in3(N__22251),
            .lcout(cmd_rdadcbuf_11),
            .ltout(),
            .carryin(\ADC_VDC.n19673 ),
            .carryout(\ADC_VDC.n19674 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__23654),
            .in2(N__24062),
            .in3(N__22248),
            .lcout(cmd_rdadcbuf_12),
            .ltout(),
            .carryin(\ADC_VDC.n19674 ),
            .carryout(\ADC_VDC.n19675 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__23642),
            .in2(N__24037),
            .in3(N__22245),
            .lcout(cmd_rdadcbuf_13),
            .ltout(),
            .carryin(\ADC_VDC.n19675 ),
            .carryout(\ADC_VDC.n19676 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__23960),
            .in2(N__23626),
            .in3(N__22242),
            .lcout(cmd_rdadcbuf_14),
            .ltout(),
            .carryin(\ADC_VDC.n19676 ),
            .carryout(\ADC_VDC.n19677 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__24092),
            .in2(N__23948),
            .in3(N__22239),
            .lcout(cmd_rdadcbuf_15),
            .ltout(),
            .carryin(\ADC_VDC.n19677 ),
            .carryout(\ADC_VDC.n19678 ),
            .clk(N__53278),
            .ce(N__22513),
            .sr(N__22447));
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__22232),
            .in2(N__23917),
            .in3(N__22221),
            .lcout(cmd_rdadcbuf_16),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\ADC_VDC.n19679 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__24350),
            .in2(N__22377),
            .in3(N__22359),
            .lcout(cmd_rdadcbuf_17),
            .ltout(),
            .carryin(\ADC_VDC.n19679 ),
            .carryout(\ADC_VDC.n19680 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__23537),
            .in2(N__23762),
            .in3(N__22356),
            .lcout(cmd_rdadcbuf_18),
            .ltout(),
            .carryin(\ADC_VDC.n19680 ),
            .carryout(\ADC_VDC.n19681 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__23690),
            .in2(N__23734),
            .in3(N__22353),
            .lcout(cmd_rdadcbuf_19),
            .ltout(),
            .carryin(\ADC_VDC.n19681 ),
            .carryout(\ADC_VDC.n19682 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__24269),
            .in2(N__22349),
            .in3(N__22326),
            .lcout(cmd_rdadcbuf_20),
            .ltout(),
            .carryin(\ADC_VDC.n19682 ),
            .carryout(\ADC_VDC.n19683 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__25763),
            .in2(N__22323),
            .in3(N__22305),
            .lcout(cmd_rdadcbuf_21),
            .ltout(),
            .carryin(\ADC_VDC.n19683 ),
            .carryout(\ADC_VDC.n19684 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__24257),
            .in2(N__26051),
            .in3(N__22302),
            .lcout(cmd_rdadcbuf_22),
            .ltout(),
            .carryin(\ADC_VDC.n19684 ),
            .carryout(\ADC_VDC.n19685 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__24320),
            .in2(N__26028),
            .in3(N__22299),
            .lcout(cmd_rdadcbuf_23),
            .ltout(),
            .carryin(\ADC_VDC.n19685 ),
            .carryout(\ADC_VDC.n19686 ),
            .clk(N__53276),
            .ce(N__22519),
            .sr(N__22454));
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__24365),
            .in2(_gnd_net_),
            .in3(N__22296),
            .lcout(cmd_rdadcbuf_24),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\ADC_VDC.n19687 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__23705),
            .in2(_gnd_net_),
            .in3(N__22293),
            .lcout(cmd_rdadcbuf_25),
            .ltout(),
            .carryin(\ADC_VDC.n19687 ),
            .carryout(\ADC_VDC.n19688 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__26066),
            .in2(_gnd_net_),
            .in3(N__22545),
            .lcout(cmd_rdadcbuf_26),
            .ltout(),
            .carryin(\ADC_VDC.n19688 ),
            .carryout(\ADC_VDC.n19689 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__23378),
            .in2(_gnd_net_),
            .in3(N__22542),
            .lcout(cmd_rdadcbuf_27),
            .ltout(),
            .carryin(\ADC_VDC.n19689 ),
            .carryout(\ADC_VDC.n19690 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__24245),
            .in2(_gnd_net_),
            .in3(N__22539),
            .lcout(cmd_rdadcbuf_28),
            .ltout(),
            .carryin(\ADC_VDC.n19690 ),
            .carryout(\ADC_VDC.n19691 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__24527),
            .in2(_gnd_net_),
            .in3(N__22536),
            .lcout(cmd_rdadcbuf_29),
            .ltout(),
            .carryin(\ADC_VDC.n19691 ),
            .carryout(\ADC_VDC.n19692 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__24539),
            .in2(_gnd_net_),
            .in3(N__22533),
            .lcout(cmd_rdadcbuf_30),
            .ltout(),
            .carryin(\ADC_VDC.n19692 ),
            .carryout(\ADC_VDC.n19693 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__24551),
            .in2(_gnd_net_),
            .in3(N__22530),
            .lcout(cmd_rdadcbuf_31),
            .ltout(),
            .carryin(\ADC_VDC.n19693 ),
            .carryout(\ADC_VDC.n19694 ),
            .clk(N__53301),
            .ce(N__22515),
            .sr(N__22451));
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__24584),
            .in2(_gnd_net_),
            .in3(N__22527),
            .lcout(cmd_rdadcbuf_32),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\ADC_VDC.n19695 ),
            .clk(N__53318),
            .ce(N__22520),
            .sr(N__22455));
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__25802),
            .in2(_gnd_net_),
            .in3(N__22524),
            .lcout(cmd_rdadcbuf_33),
            .ltout(),
            .carryin(\ADC_VDC.n19695 ),
            .carryout(\ADC_VDC.n19696 ),
            .clk(N__53318),
            .ce(N__22520),
            .sr(N__22455));
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .C_ON=1'b0;
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.add_23_36_lut_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__24233),
            .in2(_gnd_net_),
            .in3(N__22389),
            .lcout(\ADC_VDC.cmd_rdadcbuf_35_N_1138_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18591_3_lut_LC_8_11_0.C_ON=1'b0;
    defparam i18591_3_lut_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam i18591_3_lut_LC_8_11_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18591_3_lut_LC_8_11_0 (
            .in0(N__23367),
            .in1(N__22675),
            .in2(_gnd_net_),
            .in3(N__57777),
            .lcout(n21201),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_8_11_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_8_11_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i4_LC_8_11_1  (
            .in0(N__22659),
            .in1(N__28097),
            .in2(N__35585),
            .in3(N__27026),
            .lcout(cmd_rdadctmp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54328),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i23_LC_8_11_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i23_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i23_LC_8_11_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i23_LC_8_11_2  (
            .in0(N__33377),
            .in1(N__33649),
            .in2(N__22875),
            .in3(N__24184),
            .lcout(buf_adcdata_vac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54328),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i20_LC_8_11_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i20_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i20_LC_8_11_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i20_LC_8_11_3  (
            .in0(N__33647),
            .in1(N__33379),
            .in2(N__25091),
            .in3(N__22612),
            .lcout(buf_adcdata_vac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54328),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_8_11_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_8_11_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i28_LC_8_11_4  (
            .in0(N__33378),
            .in1(N__31671),
            .in2(N__22614),
            .in3(N__22638),
            .lcout(cmd_rdadctmp_28_adj_1422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54328),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i21_LC_8_11_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i21_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i21_LC_8_11_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i21_LC_8_11_6  (
            .in0(N__33376),
            .in1(N__33648),
            .in2(N__22595),
            .in3(N__22810),
            .lcout(buf_adcdata_vac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54328),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_8_11_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_8_11_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i8_LC_8_11_7  (
            .in0(N__31672),
            .in1(N__26923),
            .in2(N__22569),
            .in3(N__33380),
            .lcout(cmd_rdadctmp_8_adj_1442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54328),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_8_12_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_8_12_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i22_LC_8_12_1  (
            .in0(N__31656),
            .in1(N__24946),
            .in2(N__24902),
            .in3(N__33484),
            .lcout(cmd_rdadctmp_22_adj_1428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54342),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_8_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_8_12_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i10_LC_8_12_4  (
            .in0(N__33481),
            .in1(N__33734),
            .in2(N__28333),
            .in3(N__31655),
            .lcout(cmd_rdadctmp_10_adj_1440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54342),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_8_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_8_12_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i31_LC_8_12_5  (
            .in0(N__31658),
            .in1(N__22855),
            .in2(N__22874),
            .in3(N__33485),
            .lcout(cmd_rdadctmp_31_adj_1419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54342),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_8_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_8_12_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i26_LC_8_12_6  (
            .in0(N__33482),
            .in1(N__24412),
            .in2(N__24484),
            .in3(N__31657),
            .lcout(cmd_rdadctmp_26_adj_1424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54342),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i22_LC_8_12_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i22_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i22_LC_8_12_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i22_LC_8_12_7  (
            .in0(N__33657),
            .in1(N__33483),
            .in2(N__40429),
            .in3(N__22856),
            .lcout(buf_adcdata_vac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54342),
            .ce(),
            .sr(_gnd_net_));
    defparam n22405_bdd_4_lut_LC_8_13_0.C_ON=1'b0;
    defparam n22405_bdd_4_lut_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam n22405_bdd_4_lut_LC_8_13_0.LUT_INIT=16'b1011101010011000;
    LogicCell40 n22405_bdd_4_lut_LC_8_13_0 (
            .in0(N__22839),
            .in1(N__55170),
            .in2(N__22820),
            .in3(N__24573),
            .lcout(n21097),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i4_LC_8_13_1.C_ON=1'b0;
    defparam buf_cfgRTD_i4_LC_8_13_1.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i4_LC_8_13_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i4_LC_8_13_1 (
            .in0(N__56560),
            .in1(N__27296),
            .in2(N__41496),
            .in3(N__22756),
            .lcout(buf_cfgRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54356),
            .ce(),
            .sr(_gnd_net_));
    defparam i18529_3_lut_LC_8_13_3.C_ON=1'b0;
    defparam i18529_3_lut_LC_8_13_3.SEQ_MODE=4'b0000;
    defparam i18529_3_lut_LC_8_13_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18529_3_lut_LC_8_13_3 (
            .in0(N__57794),
            .in1(N__27344),
            .in2(_gnd_net_),
            .in3(N__27629),
            .lcout(n21139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19778_LC_8_13_4.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19778_LC_8_13_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19778_LC_8_13_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19778_LC_8_13_4 (
            .in0(N__22755),
            .in1(N__57795),
            .in2(N__22737),
            .in3(N__55171),
            .lcout(n22417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i7_LC_8_13_5.C_ON=1'b0;
    defparam buf_device_acadc_i7_LC_8_13_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i7_LC_8_13_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i7_LC_8_13_5 (
            .in0(N__56561),
            .in1(N__44862),
            .in2(N__45362),
            .in3(N__31885),
            .lcout(VAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54356),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19621_LC_8_13_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19621_LC_8_13_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19621_LC_8_13_6.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19621_LC_8_13_6 (
            .in0(N__24591),
            .in1(N__55172),
            .in2(N__22710),
            .in3(N__53786),
            .lcout(n22231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_8_13_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_8_13_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i25_LC_8_13_7  (
            .in0(N__35551),
            .in1(N__27373),
            .in2(N__31964),
            .in3(N__28112),
            .lcout(cmd_rdadctmp_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54356),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_5_i23_3_lut_LC_8_14_0.C_ON=1'b0;
    defparam mux_128_Mux_5_i23_3_lut_LC_8_14_0.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_5_i23_3_lut_LC_8_14_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_5_i23_3_lut_LC_8_14_0 (
            .in0(N__23051),
            .in1(N__57786),
            .in2(_gnd_net_),
            .in3(N__32247),
            .lcout(),
            .ltout(n23_adj_1540_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18513_4_lut_LC_8_14_1.C_ON=1'b0;
    defparam i18513_4_lut_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam i18513_4_lut_LC_8_14_1.LUT_INIT=16'b0111010000110000;
    LogicCell40 i18513_4_lut_LC_8_14_1 (
            .in0(N__57787),
            .in1(N__55162),
            .in2(N__23028),
            .in3(N__33948),
            .lcout(n21123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam EIS_SYNCCLK_I_0_1_lut_LC_8_14_2.C_ON=1'b0;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_8_14_2.SEQ_MODE=4'b0000;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_8_14_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 EIS_SYNCCLK_I_0_1_lut_LC_8_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23019),
            .lcout(IAC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i7_LC_8_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i7_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i7_LC_8_14_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i7_LC_8_14_3  (
            .in0(N__35531),
            .in1(N__35756),
            .in2(N__22956),
            .in3(N__24826),
            .lcout(buf_adcdata_iac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54368),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19704_LC_8_14_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19704_LC_8_14_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19704_LC_8_14_4.LUT_INIT=16'b1101101011010000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19704_LC_8_14_4 (
            .in0(N__53779),
            .in1(N__22932),
            .in2(N__55213),
            .in3(N__27060),
            .lcout(n22327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19689_LC_8_14_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19689_LC_8_14_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19689_LC_8_14_5.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19689_LC_8_14_5 (
            .in0(N__22920),
            .in1(N__55164),
            .in2(N__23196),
            .in3(N__53778),
            .lcout(n22291),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19729_LC_8_14_6.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19729_LC_8_14_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19729_LC_8_14_6.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19729_LC_8_14_6 (
            .in0(N__55163),
            .in1(N__23173),
            .in2(N__24997),
            .in3(N__57788),
            .lcout(),
            .ltout(n22315_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22315_bdd_4_lut_LC_8_14_7.C_ON=1'b0;
    defparam n22315_bdd_4_lut_LC_8_14_7.SEQ_MODE=4'b0000;
    defparam n22315_bdd_4_lut_LC_8_14_7.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22315_bdd_4_lut_LC_8_14_7 (
            .in0(N__41630),
            .in1(N__27180),
            .in2(N__22911),
            .in3(N__55165),
            .lcout(n22318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_15_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_15_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i14_LC_8_15_0  (
            .in0(N__35806),
            .in1(N__35458),
            .in2(N__22902),
            .in3(N__47032),
            .lcout(buf_adcdata_iac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54382),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_80_LC_8_15_2.C_ON=1'b0;
    defparam i1_2_lut_adj_80_LC_8_15_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_80_LC_8_15_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_80_LC_8_15_2 (
            .in0(_gnd_net_),
            .in1(N__30721),
            .in2(_gnd_net_),
            .in3(N__27449),
            .lcout(n20853),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i6_LC_8_15_3.C_ON=1'b0;
    defparam buf_cfgRTD_i6_LC_8_15_3.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i6_LC_8_15_3.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_cfgRTD_i6_LC_8_15_3 (
            .in0(N__27295),
            .in1(N__45357),
            .in2(N__56568),
            .in3(N__31352),
            .lcout(buf_cfgRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54382),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i0_LC_8_15_4.C_ON=1'b0;
    defparam buf_cfgRTD_i0_LC_8_15_4.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i0_LC_8_15_4.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_cfgRTD_i0_LC_8_15_4 (
            .in0(N__23220),
            .in1(N__56563),
            .in2(N__43829),
            .in3(N__27294),
            .lcout(buf_cfgRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54382),
            .ce(),
            .sr(_gnd_net_));
    defparam i18592_3_lut_LC_8_15_5.C_ON=1'b0;
    defparam i18592_3_lut_LC_8_15_5.SEQ_MODE=4'b0000;
    defparam i18592_3_lut_LC_8_15_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18592_3_lut_LC_8_15_5 (
            .in0(N__57785),
            .in1(N__23276),
            .in2(_gnd_net_),
            .in3(N__23219),
            .lcout(n21202),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i6_LC_8_15_7.C_ON=1'b0;
    defparam buf_device_acadc_i6_LC_8_15_7.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i6_LC_8_15_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i6_LC_8_15_7 (
            .in0(N__56562),
            .in1(N__44861),
            .in2(N__43601),
            .in3(N__23174),
            .lcout(VAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54382),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i8_LC_8_16_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i8_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i8_LC_8_16_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i8_LC_8_16_0  (
            .in0(N__35492),
            .in1(N__35702),
            .in2(N__43504),
            .in3(N__23157),
            .lcout(buf_adcdata_iac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54396),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i9_LC_8_16_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i9_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i9_LC_8_16_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i9_LC_8_16_1  (
            .in0(N__35701),
            .in1(N__35495),
            .in2(N__23127),
            .in3(N__37159),
            .lcout(buf_adcdata_iac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54396),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_8_16_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_8_16_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i18_LC_8_16_2  (
            .in0(N__35493),
            .in1(N__23123),
            .in2(N__28118),
            .in3(N__23338),
            .lcout(cmd_rdadctmp_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54396),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_adj_5_LC_8_16_3 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_adj_5_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_adj_5_LC_8_16_3 .LUT_INIT=16'b0000000101000100;
    LogicCell40 \ADC_VAC.i1_4_lut_adj_5_LC_8_16_3  (
            .in0(N__33218),
            .in1(N__30709),
            .in2(N__23103),
            .in3(N__27441),
            .lcout(\ADC_VAC.n12594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_16_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i19_LC_8_16_4  (
            .in0(N__35494),
            .in1(N__23339),
            .in2(N__31993),
            .in3(N__28091),
            .lcout(cmd_rdadctmp_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54396),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.SCLK_35_LC_8_16_5 .C_ON=1'b0;
    defparam \ADC_IAC.SCLK_35_LC_8_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.SCLK_35_LC_8_16_5 .LUT_INIT=16'b1011111000000010;
    LogicCell40 \ADC_IAC.SCLK_35_LC_8_16_5  (
            .in0(N__30002),
            .in1(N__35496),
            .in2(N__29916),
            .in3(N__23306),
            .lcout(IAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54396),
            .ce(),
            .sr(_gnd_net_));
    defparam i15343_2_lut_3_lut_LC_8_16_6.C_ON=1'b0;
    defparam i15343_2_lut_3_lut_LC_8_16_6.SEQ_MODE=4'b0000;
    defparam i15343_2_lut_3_lut_LC_8_16_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15343_2_lut_3_lut_LC_8_16_6 (
            .in0(N__47794),
            .in1(N__51994),
            .in2(_gnd_net_),
            .in3(N__55560),
            .lcout(n14_adj_1553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.bit_cnt_i0_LC_8_17_0 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i0_LC_8_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i0_LC_8_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i0_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__25422),
            .in2(_gnd_net_),
            .in3(N__23295),
            .lcout(\ADC_IAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\ADC_IAC.n19649 ),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.bit_cnt_i1_LC_8_17_1 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i1_LC_8_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i1_LC_8_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i1_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__25571),
            .in2(_gnd_net_),
            .in3(N__23292),
            .lcout(\ADC_IAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_IAC.n19649 ),
            .carryout(\ADC_IAC.n19650 ),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.bit_cnt_i2_LC_8_17_2 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i2_LC_8_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i2_LC_8_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i2_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__25623),
            .in2(_gnd_net_),
            .in3(N__23289),
            .lcout(\ADC_IAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_IAC.n19650 ),
            .carryout(\ADC_IAC.n19651 ),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.bit_cnt_i3_LC_8_17_3 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i3_LC_8_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i3_LC_8_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i3_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__25598),
            .in2(_gnd_net_),
            .in3(N__23286),
            .lcout(\ADC_IAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_IAC.n19651 ),
            .carryout(\ADC_IAC.n19652 ),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.bit_cnt_i4_LC_8_17_4 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i4_LC_8_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i4_LC_8_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i4_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__25584),
            .in2(_gnd_net_),
            .in3(N__23283),
            .lcout(\ADC_IAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_IAC.n19652 ),
            .carryout(\ADC_IAC.n19653 ),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.bit_cnt_i5_LC_8_17_5 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i5_LC_8_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i5_LC_8_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i5_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__25611),
            .in2(_gnd_net_),
            .in3(N__23280),
            .lcout(\ADC_IAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_IAC.n19653 ),
            .carryout(\ADC_IAC.n19654 ),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.bit_cnt_i6_LC_8_17_6 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i6_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i6_LC_8_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i6_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__25436),
            .in2(_gnd_net_),
            .in3(N__23526),
            .lcout(\ADC_IAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_IAC.n19654 ),
            .carryout(\ADC_IAC.n19655 ),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.bit_cnt_i7_LC_8_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.bit_cnt_i7_LC_8_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i7_LC_8_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i7_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__25559),
            .in2(_gnd_net_),
            .in3(N__23523),
            .lcout(\ADC_IAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54411),
            .ce(N__25878),
            .sr(N__23520));
    defparam \ADC_IAC.adc_state_i0_LC_8_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i0_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i0_LC_8_18_3 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \ADC_IAC.adc_state_i0_LC_8_18_3  (
            .in0(N__35402),
            .in1(N__29890),
            .in2(N__29996),
            .in3(N__25542),
            .lcout(adc_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54420),
            .ce(N__25635),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i30_4_lut_LC_8_19_1 .C_ON=1'b0;
    defparam \ADC_IAC.i30_4_lut_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i30_4_lut_LC_8_19_1 .LUT_INIT=16'b1100100001010001;
    LogicCell40 \ADC_IAC.i30_4_lut_LC_8_19_1  (
            .in0(N__29967),
            .in1(N__29899),
            .in2(N__25922),
            .in3(N__25392),
            .lcout(),
            .ltout(\ADC_IAC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19367_2_lut_LC_8_19_2 .C_ON=1'b0;
    defparam \ADC_IAC.i19367_2_lut_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19367_2_lut_LC_8_19_2 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \ADC_IAC.i19367_2_lut_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23508),
            .in3(N__35401),
            .lcout(\ADC_IAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i8_4_lut_LC_9_3_2 .C_ON=1'b0;
    defparam \ADC_VDC.i8_4_lut_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i8_4_lut_LC_9_3_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i8_4_lut_LC_9_3_2  (
            .in0(N__23498),
            .in1(N__23486),
            .in2(N__23475),
            .in3(N__23459),
            .lcout(\ADC_VDC.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i9_4_lut_LC_9_3_6 .C_ON=1'b0;
    defparam \ADC_VDC.i9_4_lut_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i9_4_lut_LC_9_3_6 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \ADC_VDC.i9_4_lut_LC_9_3_6  (
            .in0(N__23441),
            .in1(N__23429),
            .in2(N__23418),
            .in3(N__23402),
            .lcout(\ADC_VDC.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_5_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i16_LC_9_5_0  (
            .in0(N__25685),
            .in1(N__48797),
            .in2(N__23363),
            .in3(N__23385),
            .lcout(buf_adcdata_vdc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53253),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_21_LC_9_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_21_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_21_LC_9_5_1 .LUT_INIT=16'b1011000011100000;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_21_LC_9_5_1  (
            .in0(N__48563),
            .in1(N__47367),
            .in2(N__48851),
            .in3(N__48349),
            .lcout(\ADC_VDC.n12899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i8_LC_9_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i8_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i8_LC_9_5_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i8_LC_9_5_5  (
            .in0(N__48796),
            .in1(N__25686),
            .in2(N__23672),
            .in3(N__23694),
            .lcout(buf_adcdata_vdc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53253),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7  (
            .in0(N__48564),
            .in1(N__23579),
            .in2(N__24161),
            .in3(N__23807),
            .lcout(cmd_rdadctmp_5_adj_1474),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53253),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i1_LC_9_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i1_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i1_LC_9_6_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i1_LC_9_6_0  (
            .in0(N__25687),
            .in1(N__48846),
            .in2(N__32864),
            .in3(N__23655),
            .lcout(buf_adcdata_vdc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53260),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_6_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i2_LC_9_6_1  (
            .in0(N__48845),
            .in1(N__25688),
            .in2(N__28226),
            .in3(N__23643),
            .lcout(buf_adcdata_vdc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53260),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2  (
            .in0(N__48565),
            .in1(N__23557),
            .in2(N__24012),
            .in3(N__23814),
            .lcout(cmd_rdadctmp_9_adj_1470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53260),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_3 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_3  (
            .in0(N__23944),
            .in1(N__23631),
            .in2(N__23839),
            .in3(N__48566),
            .lcout(cmd_rdadctmp_15_adj_1464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53260),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_9_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_9_6_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i4_LC_9_6_7  (
            .in0(N__23578),
            .in1(N__23600),
            .in2(N__23840),
            .in3(N__48567),
            .lcout(cmd_rdadctmp_4_adj_1475),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53260),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_0  (
            .in0(N__24107),
            .in1(N__23558),
            .in2(N__23894),
            .in3(N__48579),
            .lcout(cmd_rdadctmp_8_adj_1471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i7_LC_9_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i7_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i7_LC_9_7_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.ADC_DATA_i7_LC_9_7_1  (
            .in0(N__23538),
            .in1(N__24308),
            .in2(N__25752),
            .in3(N__48834),
            .lcout(buf_adcdata_vdc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_9_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_9_7_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i6_LC_9_7_2  (
            .in0(N__24127),
            .in1(N__24162),
            .in2(N__23893),
            .in3(N__48578),
            .lcout(cmd_rdadctmp_6_adj_1473),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_9_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_9_7_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i7_LC_9_7_3  (
            .in0(N__48576),
            .in1(N__24108),
            .in2(N__24135),
            .in3(N__23880),
            .lcout(cmd_rdadctmp_7_adj_1472),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i4_LC_9_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i4_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i4_LC_9_7_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i4_LC_9_7_4  (
            .in0(N__48832),
            .in1(N__25736),
            .in2(N__24080),
            .in3(N__24093),
            .lcout(buf_adcdata_vdc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_7_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i13_LC_9_7_5  (
            .in0(N__48575),
            .in1(N__24063),
            .in2(N__24039),
            .in3(N__23876),
            .lcout(cmd_rdadctmp_13_adj_1466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_7_6 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i10_LC_9_7_6  (
            .in0(N__23983),
            .in1(N__24010),
            .in2(N__23892),
            .in3(N__48577),
            .lcout(cmd_rdadctmp_10_adj_1469),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i3_LC_9_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i3_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i3_LC_9_7_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i3_LC_9_7_7  (
            .in0(N__25735),
            .in1(N__48833),
            .in2(N__27866),
            .in3(N__23964),
            .lcout(buf_adcdata_vdc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_9_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_9_8_0 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i16_LC_9_8_0  (
            .in0(N__23921),
            .in1(N__23949),
            .in2(N__23895),
            .in3(N__48591),
            .lcout(cmd_rdadctmp_16_adj_1463),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_9_8_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_9_8_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i19_LC_9_8_1  (
            .in0(N__48590),
            .in1(N__23887),
            .in2(N__23735),
            .in3(N__23766),
            .lcout(cmd_rdadctmp_19_adj_1460),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i14_LC_9_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i14_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i14_LC_9_8_2 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i14_LC_9_8_2  (
            .in0(N__23709),
            .in1(N__46364),
            .in2(N__48872),
            .in3(N__25742),
            .lcout(buf_adcdata_vdc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i13_LC_9_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i13_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i13_LC_9_8_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i13_LC_9_8_3  (
            .in0(N__25741),
            .in1(N__48854),
            .in2(N__24965),
            .in3(N__24366),
            .lcout(buf_adcdata_vdc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i6_LC_9_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i6_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i6_LC_9_8_4 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i6_LC_9_8_4  (
            .in0(N__24354),
            .in1(N__24332),
            .in2(N__48873),
            .in3(N__25743),
            .lcout(buf_adcdata_vdc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i12_LC_9_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i12_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i12_LC_9_8_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i12_LC_9_8_5  (
            .in0(N__25740),
            .in1(N__48853),
            .in2(N__24608),
            .in3(N__24321),
            .lcout(buf_adcdata_vdc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i19_3_lut_LC_9_8_6.C_ON=1'b0;
    defparam mux_130_Mux_7_i19_3_lut_LC_9_8_6.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i19_3_lut_LC_9_8_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_130_Mux_7_i19_3_lut_LC_9_8_6 (
            .in0(N__24309),
            .in1(N__57699),
            .in2(_gnd_net_),
            .in3(N__24293),
            .lcout(n19_adj_1623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i9_LC_9_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i9_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i9_LC_9_8_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i9_LC_9_8_7  (
            .in0(N__25744),
            .in1(N__48855),
            .in2(N__34958),
            .in3(N__24270),
            .lcout(buf_adcdata_vdc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_9_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_9_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i11_LC_9_9_0  (
            .in0(N__25745),
            .in1(N__48865),
            .in2(N__50939),
            .in3(N__24258),
            .lcout(buf_adcdata_vdc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i17_LC_9_9_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i17_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i17_LC_9_9_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i17_LC_9_9_1  (
            .in0(N__48862),
            .in1(N__25746),
            .in2(N__24453),
            .in3(N__24246),
            .lcout(buf_adcdata_vdc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i23_LC_9_9_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i23_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i23_LC_9_9_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i23_LC_9_9_2  (
            .in0(N__25751),
            .in1(N__48868),
            .in2(N__24207),
            .in3(N__24234),
            .lcout(buf_adcdata_vdc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16192_3_lut_LC_9_9_3 .C_ON=1'b0;
    defparam \ADC_VDC.i16192_3_lut_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16192_3_lut_LC_9_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ADC_VDC.i16192_3_lut_LC_9_9_3  (
            .in0(N__24206),
            .in1(N__24185),
            .in2(_gnd_net_),
            .in3(N__57776),
            .lcout(n19_adj_1527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i21_LC_9_9_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i21_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i21_LC_9_9_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i21_LC_9_9_4  (
            .in0(N__25750),
            .in1(N__48867),
            .in2(N__24569),
            .in3(N__24585),
            .lcout(buf_adcdata_vdc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i20_LC_9_9_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i20_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i20_LC_9_9_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i20_LC_9_9_5  (
            .in0(N__48864),
            .in1(N__25749),
            .in2(N__25058),
            .in3(N__24552),
            .lcout(buf_adcdata_vdc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i19_LC_9_9_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i19_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i19_LC_9_9_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i19_LC_9_9_6  (
            .in0(N__25748),
            .in1(N__48866),
            .in2(N__25235),
            .in3(N__24540),
            .lcout(buf_adcdata_vdc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i18_LC_9_9_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i18_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i18_LC_9_9_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i18_LC_9_9_7  (
            .in0(N__48863),
            .in1(N__25747),
            .in2(N__27101),
            .in3(N__24528),
            .lcout(buf_adcdata_vdc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i15_LC_9_10_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i15_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i15_LC_9_10_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i15_LC_9_10_0  (
            .in0(N__33345),
            .in1(N__33673),
            .in2(N__24516),
            .in3(N__50201),
            .lcout(buf_adcdata_vac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i18_LC_9_10_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i18_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i18_LC_9_10_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i18_LC_9_10_1  (
            .in0(N__33672),
            .in1(N__33347),
            .in2(N__24489),
            .in3(N__27080),
            .lcout(buf_adcdata_vac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(),
            .sr(_gnd_net_));
    defparam n22441_bdd_4_lut_LC_9_10_2.C_ON=1'b0;
    defparam n22441_bdd_4_lut_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam n22441_bdd_4_lut_LC_9_10_2.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22441_bdd_4_lut_LC_9_10_2 (
            .in0(N__24379),
            .in1(N__24452),
            .in2(N__24438),
            .in3(N__55175),
            .lcout(n22444),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i17_LC_9_10_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i17_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i17_LC_9_10_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i17_LC_9_10_3  (
            .in0(N__33671),
            .in1(N__33346),
            .in2(N__24423),
            .in3(N__24380),
            .lcout(buf_adcdata_vac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_9_10_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_9_10_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i7_LC_9_10_4  (
            .in0(N__28098),
            .in1(N__27045),
            .in2(N__24743),
            .in3(N__35579),
            .lcout(cmd_rdadctmp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54303),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i22_3_lut_LC_9_10_6.C_ON=1'b0;
    defparam mux_130_Mux_7_i22_3_lut_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i22_3_lut_LC_9_10_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_130_Mux_7_i22_3_lut_LC_9_10_6 (
            .in0(N__53777),
            .in1(N__24833),
            .in2(_gnd_net_),
            .in3(N__24804),
            .lcout(),
            .ltout(n22_adj_1624_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i30_3_lut_LC_9_10_7.C_ON=1'b0;
    defparam mux_130_Mux_7_i30_3_lut_LC_9_10_7.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i30_3_lut_LC_9_10_7.LUT_INIT=16'b1101100011011000;
    LogicCell40 mux_130_Mux_7_i30_3_lut_LC_9_10_7 (
            .in0(N__54706),
            .in1(N__24795),
            .in2(N__24780),
            .in3(_gnd_net_),
            .lcout(n30_adj_1625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i0_LC_9_11_0 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i0_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i0_LC_9_11_0 .LUT_INIT=16'b0000111101000000;
    LogicCell40 \CLK_DDS.bit_cnt_i0_LC_9_11_0  (
            .in0(N__34610),
            .in1(N__34463),
            .in2(N__34797),
            .in3(N__24763),
            .lcout(bit_cnt_0_adj_1456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54316),
            .ce(),
            .sr(_gnd_net_));
    defparam i15170_2_lut_LC_9_11_2.C_ON=1'b0;
    defparam i15170_2_lut_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam i15170_2_lut_LC_9_11_2.LUT_INIT=16'b1100110011111111;
    LogicCell40 i15170_2_lut_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(N__51905),
            .in2(_gnd_net_),
            .in3(N__49493),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3  (
            .in0(N__26867),
            .in1(N__28093),
            .in2(N__24747),
            .in3(N__35616),
            .lcout(cmd_rdadctmp_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54316),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.MOSI_31_LC_9_11_4 .C_ON=1'b0;
    defparam \CLK_DDS.MOSI_31_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.MOSI_31_LC_9_11_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \CLK_DDS.MOSI_31_LC_9_11_4  (
            .in0(N__34776),
            .in1(_gnd_net_),
            .in2(N__27228),
            .in3(N__24707),
            .lcout(DDS_MOSI1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54316),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19783_LC_9_11_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19783_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19783_LC_9_11_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19783_LC_9_11_5 (
            .in0(N__24678),
            .in1(N__55169),
            .in2(N__24636),
            .in3(N__57642),
            .lcout(n22435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i8_LC_9_11_6.C_ON=1'b0;
    defparam buf_dds1_i8_LC_9_11_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i8_LC_9_11_6.LUT_INIT=16'b1100000010001000;
    LogicCell40 buf_dds1_i8_LC_9_11_6 (
            .in0(N__27200),
            .in1(N__40669),
            .in2(N__43835),
            .in3(N__44975),
            .lcout(buf_dds1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54316),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i19_3_lut_LC_9_12_0.C_ON=1'b0;
    defparam mux_129_Mux_4_i19_3_lut_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i19_3_lut_LC_9_12_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_129_Mux_4_i19_3_lut_LC_9_12_0 (
            .in0(N__57668),
            .in1(N__24850),
            .in2(_gnd_net_),
            .in3(N__24612),
            .lcout(n19_adj_1511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_1  (
            .in0(N__33477),
            .in1(N__31515),
            .in2(N__24879),
            .in3(N__31686),
            .lcout(cmd_rdadctmp_20_adj_1430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54329),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i14_LC_9_12_2.C_ON=1'b0;
    defparam buf_dds1_i14_LC_9_12_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i14_LC_9_12_2.LUT_INIT=16'b1100000010001000;
    LogicCell40 buf_dds1_i14_LC_9_12_2 (
            .in0(N__28606),
            .in1(N__40670),
            .in2(N__45339),
            .in3(N__44976),
            .lcout(buf_dds1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54329),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i19_3_lut_LC_9_12_3.C_ON=1'b0;
    defparam mux_129_Mux_5_i19_3_lut_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i19_3_lut_LC_9_12_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_5_i19_3_lut_LC_9_12_3 (
            .in0(N__24969),
            .in1(N__24916),
            .in2(_gnd_net_),
            .in3(N__57667),
            .lcout(n19_adj_1497),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_9_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_9_12_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i21_LC_9_12_4  (
            .in0(N__31687),
            .in1(N__24877),
            .in2(N__24947),
            .in3(N__33480),
            .lcout(cmd_rdadctmp_21_adj_1429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54329),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_9_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_9_12_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i9_LC_9_12_5  (
            .in0(N__33478),
            .in1(N__33733),
            .in2(N__26930),
            .in3(N__31688),
            .lcout(cmd_rdadctmp_9_adj_1441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54329),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i13_LC_9_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i13_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i13_LC_9_12_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i13_LC_9_12_6  (
            .in0(N__24917),
            .in1(N__33658),
            .in2(N__24948),
            .in3(N__33479),
            .lcout(buf_adcdata_vac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54329),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i14_LC_9_12_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i14_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i14_LC_9_12_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i14_LC_9_12_7  (
            .in0(N__33476),
            .in1(N__24901),
            .in2(N__33679),
            .in3(N__46342),
            .lcout(buf_adcdata_vac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54329),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i12_LC_9_13_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i12_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i12_LC_9_13_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i12_LC_9_13_0  (
            .in0(N__35776),
            .in1(N__35557),
            .in2(N__25041),
            .in3(N__46255),
            .lcout(buf_adcdata_iac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54343),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i12_LC_9_13_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i12_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i12_LC_9_13_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i12_LC_9_13_1  (
            .in0(N__33456),
            .in1(N__24878),
            .in2(N__33674),
            .in3(N__24854),
            .lcout(buf_adcdata_vac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54343),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i7_LC_9_13_2.C_ON=1'b0;
    defparam buf_cfgRTD_i7_LC_9_13_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i7_LC_9_13_2.LUT_INIT=16'b0111010000110000;
    LogicCell40 buf_cfgRTD_i7_LC_9_13_2 (
            .in0(N__56552),
            .in1(N__27264),
            .in2(N__31280),
            .in3(N__42803),
            .lcout(buf_cfgRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54343),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_3  (
            .in0(N__35555),
            .in1(N__25131),
            .in2(N__27374),
            .in3(N__28114),
            .lcout(cmd_rdadctmp_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54343),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_9_13_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_9_13_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i27_LC_9_13_5  (
            .in0(N__35556),
            .in1(N__27321),
            .in2(N__27590),
            .in3(N__28115),
            .lcout(cmd_rdadctmp_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54343),
            .ce(),
            .sr(_gnd_net_));
    defparam n22417_bdd_4_lut_LC_9_13_6.C_ON=1'b0;
    defparam n22417_bdd_4_lut_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam n22417_bdd_4_lut_LC_9_13_6.LUT_INIT=16'b1010101011100100;
    LogicCell40 n22417_bdd_4_lut_LC_9_13_6 (
            .in0(N__25104),
            .in1(N__25090),
            .in2(N__25062),
            .in3(N__55173),
            .lcout(n22420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_9_13_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_9_13_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i21_LC_9_13_7  (
            .in0(N__35554),
            .in1(N__25037),
            .in2(N__35233),
            .in3(N__28113),
            .lcout(cmd_rdadctmp_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54343),
            .ce(),
            .sr(_gnd_net_));
    defparam i18528_3_lut_LC_9_14_0.C_ON=1'b0;
    defparam i18528_3_lut_LC_9_14_0.SEQ_MODE=4'b0000;
    defparam i18528_3_lut_LC_9_14_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18528_3_lut_LC_9_14_0 (
            .in0(N__27201),
            .in1(N__32036),
            .in2(_gnd_net_),
            .in3(N__57796),
            .lcout(),
            .ltout(n21138_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22291_bdd_4_lut_LC_9_14_1.C_ON=1'b0;
    defparam n22291_bdd_4_lut_LC_9_14_1.SEQ_MODE=4'b0000;
    defparam n22291_bdd_4_lut_LC_9_14_1.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22291_bdd_4_lut_LC_9_14_1 (
            .in0(N__25017),
            .in1(N__25011),
            .in2(N__25005),
            .in3(N__53781),
            .lcout(n22294),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i21_LC_9_14_2 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i21_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i21_LC_9_14_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i21_LC_9_14_2  (
            .in0(N__35757),
            .in1(N__35529),
            .in2(N__24998),
            .in3(N__25201),
            .lcout(buf_adcdata_iac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54357),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_9_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_9_14_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i29_LC_9_14_3  (
            .in0(N__35527),
            .in1(N__28116),
            .in2(N__25205),
            .in3(N__27551),
            .lcout(cmd_rdadctmp_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54357),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i22_LC_9_14_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i22_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i22_LC_9_14_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i22_LC_9_14_4  (
            .in0(N__35758),
            .in1(N__25183),
            .in2(N__31933),
            .in3(N__35530),
            .lcout(buf_adcdata_iac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54357),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_9_14_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_9_14_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i31_LC_9_14_5  (
            .in0(N__35528),
            .in1(N__28117),
            .in2(N__25185),
            .in3(N__25217),
            .lcout(cmd_rdadctmp_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54357),
            .ce(),
            .sr(_gnd_net_));
    defparam n22435_bdd_4_lut_LC_9_14_6.C_ON=1'b0;
    defparam n22435_bdd_4_lut_LC_9_14_6.SEQ_MODE=4'b0000;
    defparam n22435_bdd_4_lut_LC_9_14_6.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22435_bdd_4_lut_LC_9_14_6 (
            .in0(N__25286),
            .in1(N__25251),
            .in2(N__25242),
            .in3(N__55174),
            .lcout(n21076),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i23_LC_9_14_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i23_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i23_LC_9_14_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i23_LC_9_14_7  (
            .in0(N__35526),
            .in1(N__35759),
            .in2(N__25157),
            .in3(N__25218),
            .lcout(buf_adcdata_iac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54357),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_15_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_15_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i19_LC_9_15_0  (
            .in0(N__35805),
            .in1(N__35553),
            .in2(N__27591),
            .in3(N__43216),
            .lcout(buf_adcdata_iac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54369),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_9_15_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_9_15_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i30_LC_9_15_1  (
            .in0(N__35552),
            .in1(N__25206),
            .in2(N__25184),
            .in3(N__28092),
            .lcout(cmd_rdadctmp_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54369),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i15_LC_9_15_2.C_ON=1'b0;
    defparam buf_dds1_i15_LC_9_15_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i15_LC_9_15_2.LUT_INIT=16'b1110000000100000;
    LogicCell40 buf_dds1_i15_LC_9_15_2 (
            .in0(N__27479),
            .in1(N__44977),
            .in2(N__40674),
            .in3(N__42810),
            .lcout(buf_dds1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54369),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i17_3_lut_LC_9_15_3.C_ON=1'b0;
    defparam mux_128_Mux_7_i17_3_lut_LC_9_15_3.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i17_3_lut_LC_9_15_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_7_i17_3_lut_LC_9_15_3 (
            .in0(N__25150),
            .in1(N__25351),
            .in2(_gnd_net_),
            .in3(N__57792),
            .lcout(n17_adj_1526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_6_i16_3_lut_LC_9_15_5.C_ON=1'b0;
    defparam mux_128_Mux_6_i16_3_lut_LC_9_15_5.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_6_i16_3_lut_LC_9_15_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_6_i16_3_lut_LC_9_15_5 (
            .in0(N__28607),
            .in1(N__29428),
            .in2(_gnd_net_),
            .in3(N__57793),
            .lcout(n16_adj_1534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i14_LC_9_15_6.C_ON=1'b0;
    defparam buf_dds0_i14_LC_9_15_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i14_LC_9_15_6.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_dds0_i14_LC_9_15_6 (
            .in0(N__29429),
            .in1(N__56498),
            .in2(N__45363),
            .in3(N__47986),
            .lcout(buf_dds0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54369),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i8_LC_9_15_7.C_ON=1'b0;
    defparam buf_device_acadc_i8_LC_9_15_7.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i8_LC_9_15_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i8_LC_9_15_7 (
            .in0(N__56497),
            .in1(N__44860),
            .in2(N__42815),
            .in3(N__25352),
            .lcout(VAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54369),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.bit_cnt_i0_LC_9_16_0 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i0_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i0_LC_9_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i0_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__25485),
            .in2(_gnd_net_),
            .in3(N__25338),
            .lcout(\ADC_VAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\ADC_VAC.n19656 ),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_VAC.bit_cnt_i1_LC_9_16_1 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i1_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i1_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i1_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__25511),
            .in2(_gnd_net_),
            .in3(N__25335),
            .lcout(\ADC_VAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC.n19656 ),
            .carryout(\ADC_VAC.n19657 ),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_VAC.bit_cnt_i2_LC_9_16_2 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i2_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i2_LC_9_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i2_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__25497),
            .in2(_gnd_net_),
            .in3(N__25332),
            .lcout(\ADC_VAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC.n19657 ),
            .carryout(\ADC_VAC.n19658 ),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_VAC.bit_cnt_i3_LC_9_16_3 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i3_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i3_LC_9_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i3_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__25524),
            .in2(_gnd_net_),
            .in3(N__25329),
            .lcout(\ADC_VAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC.n19658 ),
            .carryout(\ADC_VAC.n19659 ),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_VAC.bit_cnt_i4_LC_9_16_4 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i4_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i4_LC_9_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i4_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__25536),
            .in2(_gnd_net_),
            .in3(N__25326),
            .lcout(\ADC_VAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC.n19659 ),
            .carryout(\ADC_VAC.n19660 ),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_VAC.bit_cnt_i5_LC_9_16_5 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i5_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i5_LC_9_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i5_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__25316),
            .in2(_gnd_net_),
            .in3(N__25299),
            .lcout(\ADC_VAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC.n19660 ),
            .carryout(\ADC_VAC.n19661 ),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_VAC.bit_cnt_i6_LC_9_16_6 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i6_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i6_LC_9_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i6_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__25473),
            .in2(_gnd_net_),
            .in3(N__25296),
            .lcout(\ADC_VAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC.n19661 ),
            .carryout(\ADC_VAC.n19662 ),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_VAC.bit_cnt_i7_LC_9_16_7 .C_ON=1'b0;
    defparam \ADC_VAC.bit_cnt_i7_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i7_LC_9_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i7_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__25458),
            .in2(_gnd_net_),
            .in3(N__25293),
            .lcout(\ADC_VAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54383),
            .ce(N__30749),
            .sr(N__30639));
    defparam \ADC_IAC.i1_4_lut_LC_9_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_LC_9_17_0 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_IAC.i1_4_lut_LC_9_17_0  (
            .in0(N__30001),
            .in1(N__35394),
            .in2(N__25941),
            .in3(N__25391),
            .lcout(),
            .ltout(\ADC_IAC.n20960_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_2_lut_LC_9_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.i1_2_lut_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_2_lut_LC_9_17_1 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \ADC_IAC.i1_2_lut_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25638),
            .in3(N__29911),
            .lcout(\ADC_IAC.n20961 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19262_4_lut_LC_9_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.i19262_4_lut_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19262_4_lut_LC_9_17_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \ADC_IAC.i19262_4_lut_LC_9_17_3  (
            .in0(N__25622),
            .in1(N__25610),
            .in2(N__25599),
            .in3(N__25583),
            .lcout(),
            .ltout(\ADC_IAC.n21295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19068_4_lut_LC_9_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.i19068_4_lut_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19068_4_lut_LC_9_17_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ADC_IAC.i19068_4_lut_LC_9_17_4  (
            .in0(N__25572),
            .in1(N__25560),
            .in2(N__25545),
            .in3(N__25410),
            .lcout(\ADC_IAC.n21294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i18419_4_lut_LC_9_17_5 .C_ON=1'b0;
    defparam \ADC_VAC.i18419_4_lut_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i18419_4_lut_LC_9_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i18419_4_lut_LC_9_17_5  (
            .in0(N__25535),
            .in1(N__25523),
            .in2(N__25512),
            .in3(N__25496),
            .lcout(),
            .ltout(\ADC_VAC.n21029_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i18433_4_lut_LC_9_17_6 .C_ON=1'b0;
    defparam \ADC_VAC.i18433_4_lut_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i18433_4_lut_LC_9_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i18433_4_lut_LC_9_17_6  (
            .in0(N__25484),
            .in1(N__25472),
            .in2(N__25461),
            .in3(N__25457),
            .lcout(\ADC_VAC.n21043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i6_4_lut_LC_9_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.i6_4_lut_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i6_4_lut_LC_9_18_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \ADC_IAC.i6_4_lut_LC_9_18_0  (
            .in0(N__35325),
            .in1(N__29910),
            .in2(N__25437),
            .in3(N__25421),
            .lcout(\ADC_IAC.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_trig_300_LC_9_18_5.C_ON=1'b0;
    defparam acadc_trig_300_LC_9_18_5.SEQ_MODE=4'b1000;
    defparam acadc_trig_300_LC_9_18_5.LUT_INIT=16'b1101000111000000;
    LogicCell40 acadc_trig_300_LC_9_18_5 (
            .in0(N__30308),
            .in1(N__30180),
            .in2(N__25402),
            .in3(N__37297),
            .lcout(acadc_trig),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_trig_300C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_adj_3_LC_9_18_6 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_adj_3_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_adj_3_LC_9_18_6 .LUT_INIT=16'b0000000101000100;
    LogicCell40 \ADC_IAC.i1_4_lut_adj_3_LC_9_18_6  (
            .in0(N__35324),
            .in1(N__30000),
            .in2(N__25940),
            .in3(N__29909),
            .lcout(\ADC_IAC.n12473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_10_3_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_10_3_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_91_2_lut_LC_10_3_2  (
            .in0(_gnd_net_),
            .in1(N__27810),
            .in2(_gnd_net_),
            .in3(N__55831),
            .lcout(\comm_spi.iclk_N_763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19333_4_lut_4_lut_LC_10_3_5 .C_ON=1'b0;
    defparam \ADC_VDC.i19333_4_lut_4_lut_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19333_4_lut_4_lut_LC_10_3_5 .LUT_INIT=16'b1111101011101011;
    LogicCell40 \ADC_VDC.i19333_4_lut_4_lut_LC_10_3_5  (
            .in0(N__48528),
            .in1(N__48338),
            .in2(N__48836),
            .in3(N__47383),
            .lcout(),
            .ltout(\ADC_VDC.n11676_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.SCLK_46_LC_10_3_6 .C_ON=1'b0;
    defparam \ADC_VDC.SCLK_46_LC_10_3_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.SCLK_46_LC_10_3_6 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.SCLK_46_LC_10_3_6  (
            .in0(N__48339),
            .in1(N__25835),
            .in2(N__25854),
            .in3(N__27849),
            .lcout(VDC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53294),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_12178_12179_reset_LC_10_4_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12178_12179_reset_LC_10_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.iclk_40_12178_12179_reset_LC_10_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12178_12179_reset_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27822),
            .lcout(\comm_spi.n14597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54270),
            .ce(),
            .sr(N__25824));
    defparam \ADC_VDC.ADC_DATA_i22_LC_10_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i22_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i22_LC_10_5_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \ADC_VDC.ADC_DATA_i22_LC_10_5_1  (
            .in0(N__25684),
            .in1(N__25812),
            .in2(N__40451),
            .in3(N__48800),
            .lcout(buf_adcdata_vdc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53293),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i0_LC_10_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i0_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i0_LC_10_5_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i0_LC_10_5_3  (
            .in0(N__25682),
            .in1(N__48799),
            .in2(N__25964),
            .in3(N__25791),
            .lcout(buf_adcdata_vdc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53293),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i10_LC_10_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i10_LC_10_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i10_LC_10_5_4 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \ADC_VDC.ADC_DATA_i10_LC_10_5_4  (
            .in0(N__35972),
            .in1(N__48804),
            .in2(N__25773),
            .in3(N__25683),
            .lcout(buf_adcdata_vdc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53293),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_20_LC_10_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_20_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_20_LC_10_5_5 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_adj_20_LC_10_5_5  (
            .in0(N__48538),
            .in1(N__48345),
            .in2(N__48852),
            .in3(N__47366),
            .lcout(n13087),
            .ltout(n13087_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i15_LC_10_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i15_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i15_LC_10_5_6 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \ADC_VDC.ADC_DATA_i15_LC_10_5_6  (
            .in0(N__50231),
            .in1(N__48805),
            .in2(N__26076),
            .in3(N__26073),
            .lcout(buf_adcdata_vdc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53293),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_19_LC_10_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_19_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_19_LC_10_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_19_LC_10_5_7  (
            .in0(_gnd_net_),
            .in1(N__48537),
            .in2(_gnd_net_),
            .in3(N__48798),
            .lcout(\ADC_VDC.n20656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_0 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_0  (
            .in0(N__26055),
            .in1(N__48346),
            .in2(N__26024),
            .in3(N__32733),
            .lcout(\ADC_VDC.cmd_rdadctmp_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53255),
            .ce(N__26004),
            .sr(N__25992));
    defparam \comm_spi.i19415_4_lut_3_lut_LC_10_6_3 .C_ON=1'b0;
    defparam \comm_spi.i19415_4_lut_3_lut_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19415_4_lut_3_lut_LC_10_6_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \comm_spi.i19415_4_lut_3_lut_LC_10_6_3  (
            .in0(N__55833),
            .in1(_gnd_net_),
            .in2(N__27828),
            .in3(N__25983),
            .lcout(\comm_spi.n22860 ),
            .ltout(\comm_spi.n22860_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12180_3_lut_LC_10_6_4 .C_ON=1'b0;
    defparam \comm_spi.i12180_3_lut_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12180_3_lut_LC_10_6_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.i12180_3_lut_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__27780),
            .in2(N__25977),
            .in3(N__25974),
            .lcout(\comm_spi.iclk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_10_6_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_10_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_90_2_lut_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__27824),
            .in2(_gnd_net_),
            .in3(N__55832),
            .lcout(\comm_spi.iclk_N_762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i19_3_lut_LC_10_7_0.C_ON=1'b0;
    defparam mux_130_Mux_0_i19_3_lut_LC_10_7_0.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i19_3_lut_LC_10_7_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_0_i19_3_lut_LC_10_7_0 (
            .in0(N__25965),
            .in1(N__26893),
            .in2(_gnd_net_),
            .in3(N__57756),
            .lcout(),
            .ltout(n19_adj_1484_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i22_3_lut_LC_10_7_1.C_ON=1'b0;
    defparam mux_130_Mux_0_i22_3_lut_LC_10_7_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i22_3_lut_LC_10_7_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_0_i22_3_lut_LC_10_7_1 (
            .in0(_gnd_net_),
            .in1(N__26959),
            .in2(N__25947),
            .in3(N__53771),
            .lcout(),
            .ltout(n22_adj_1483_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i30_3_lut_LC_10_7_2.C_ON=1'b0;
    defparam mux_130_Mux_0_i30_3_lut_LC_10_7_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i30_3_lut_LC_10_7_2.LUT_INIT=16'b1111110000110000;
    LogicCell40 mux_130_Mux_0_i30_3_lut_LC_10_7_2 (
            .in0(_gnd_net_),
            .in1(N__54754),
            .in2(N__25944),
            .in3(N__26991),
            .lcout(n30_adj_1482),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i0_LC_10_7_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i0_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i0_LC_10_7_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i0_LC_10_7_3  (
            .in0(N__35815),
            .in1(N__26879),
            .in2(N__26966),
            .in3(N__35636),
            .lcout(buf_adcdata_iac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i0_LC_10_7_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i0_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i0_LC_10_7_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i0_LC_10_7_4  (
            .in0(N__33675),
            .in1(N__33501),
            .in2(N__26940),
            .in3(N__26894),
            .lcout(buf_adcdata_vac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_10_7_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_10_7_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i9_LC_10_7_6  (
            .in0(N__35635),
            .in1(N__28153),
            .in2(N__26880),
            .in3(N__28125),
            .lcout(cmd_rdadctmp_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54276),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.bit_cnt_3767__i3_LC_10_8_0 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i3_LC_10_8_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i3_LC_10_8_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \comm_spi.bit_cnt_3767__i3_LC_10_8_0  (
            .in0(N__28438),
            .in1(N__35884),
            .in2(N__28422),
            .in3(N__28458),
            .lcout(\comm_spi.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__55870));
    defparam \comm_spi.bit_cnt_3767__i2_LC_10_8_1 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i2_LC_10_8_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i2_LC_10_8_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \comm_spi.bit_cnt_3767__i2_LC_10_8_1  (
            .in0(N__28457),
            .in1(N__28418),
            .in2(_gnd_net_),
            .in3(N__28439),
            .lcout(\comm_spi.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__55870));
    defparam \comm_spi.bit_cnt_3767__i1_LC_10_8_2 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i1_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i1_LC_10_8_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \comm_spi.bit_cnt_3767__i1_LC_10_8_2  (
            .in0(N__28417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28456),
            .lcout(\comm_spi.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__55870));
    defparam \comm_spi.bit_cnt_3767__i0_LC_10_8_3 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i0_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i0_LC_10_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \comm_spi.bit_cnt_3767__i0_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28416),
            .lcout(\comm_spi.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__55870));
    defparam \RTD.i1_3_lut_4_lut_LC_10_9_0 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_4_lut_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_4_lut_LC_10_9_0 .LUT_INIT=16'b1010001010010100;
    LogicCell40 \RTD.i1_3_lut_4_lut_LC_10_9_0  (
            .in0(N__26850),
            .in1(N__26598),
            .in2(N__26448),
            .in3(N__26264),
            .lcout(\RTD.n15065 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i12467_3_lut_LC_10_9_4 .C_ON=1'b0;
    defparam \SIG_DDS.i12467_3_lut_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i12467_3_lut_LC_10_9_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \SIG_DDS.i12467_3_lut_LC_10_9_4  (
            .in0(N__42288),
            .in1(N__41334),
            .in2(_gnd_net_),
            .in3(N__43070),
            .lcout(n14884),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.SCLK_27_LC_10_9_5 .C_ON=1'b0;
    defparam \CLK_DDS.SCLK_27_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.SCLK_27_LC_10_9_5 .LUT_INIT=16'b0111001000110001;
    LogicCell40 \CLK_DDS.SCLK_27_LC_10_9_5  (
            .in0(N__34749),
            .in1(N__34609),
            .in2(N__27119),
            .in3(N__34457),
            .lcout(DDS_SCK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54288),
            .ce(),
            .sr(_gnd_net_));
    defparam i18471_3_lut_LC_10_9_7.C_ON=1'b0;
    defparam i18471_3_lut_LC_10_9_7.SEQ_MODE=4'b0000;
    defparam i18471_3_lut_LC_10_9_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18471_3_lut_LC_10_9_7 (
            .in0(N__27102),
            .in1(N__27076),
            .in2(_gnd_net_),
            .in3(N__57737),
            .lcout(n21081),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_10_10_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_10_10_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i6_LC_10_10_0  (
            .in0(N__27015),
            .in1(N__35570),
            .in2(N__28122),
            .in3(N__27044),
            .lcout(cmd_rdadctmp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54293),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_10_10_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_10_10_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i5_LC_10_10_1  (
            .in0(N__27033),
            .in1(N__28099),
            .in2(N__35621),
            .in3(N__27014),
            .lcout(cmd_rdadctmp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54293),
            .ce(),
            .sr(_gnd_net_));
    defparam i19404_2_lut_3_lut_LC_10_10_4.C_ON=1'b0;
    defparam i19404_2_lut_3_lut_LC_10_10_4.SEQ_MODE=4'b0000;
    defparam i19404_2_lut_3_lut_LC_10_10_4.LUT_INIT=16'b0000000000010001;
    LogicCell40 i19404_2_lut_3_lut_LC_10_10_4 (
            .in0(N__37317),
            .in1(N__30309),
            .in2(_gnd_net_),
            .in3(N__40890),
            .lcout(n21037),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i4_LC_10_10_5.C_ON=1'b0;
    defparam comm_buf_6__i4_LC_10_10_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i4_LC_10_10_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_buf_6__i4_LC_10_10_5 (
            .in0(N__35004),
            .in1(N__46762),
            .in2(N__57004),
            .in3(N__39530),
            .lcout(comm_buf_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54293),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i2_LC_10_10_6.C_ON=1'b0;
    defparam comm_buf_6__i2_LC_10_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i2_LC_10_10_6.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i2_LC_10_10_6 (
            .in0(N__39686),
            .in1(N__56868),
            .in2(N__47223),
            .in3(N__35003),
            .lcout(comm_buf_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54293),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i11_LC_10_10_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i11_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i11_LC_10_10_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i11_LC_10_10_7  (
            .in0(N__33670),
            .in1(N__33344),
            .in2(N__50920),
            .in3(N__31514),
            .lcout(buf_adcdata_vac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54293),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i7_LC_10_11_0.C_ON=1'b0;
    defparam buf_control_i7_LC_10_11_0.SEQ_MODE=4'b1000;
    defparam buf_control_i7_LC_10_11_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 buf_control_i7_LC_10_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27006),
            .lcout(buf_control_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54304),
            .ce(N__27153),
            .sr(N__39573));
    defparam i1_2_lut_adj_225_LC_10_11_1.C_ON=1'b0;
    defparam i1_2_lut_adj_225_LC_10_11_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_225_LC_10_11_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_adj_225_LC_10_11_1 (
            .in0(N__49491),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55515),
            .lcout(),
            .ltout(n11347_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_262_LC_10_11_2.C_ON=1'b0;
    defparam i1_4_lut_adj_262_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_262_LC_10_11_2.LUT_INIT=16'b1000110010001000;
    LogicCell40 i1_4_lut_adj_262_LC_10_11_2 (
            .in0(N__57064),
            .in1(N__49601),
            .in2(N__27156),
            .in3(N__52011),
            .lcout(n11919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i23_3_lut_LC_10_11_3.C_ON=1'b0;
    defparam mux_128_Mux_7_i23_3_lut_LC_10_11_3.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i23_3_lut_LC_10_11_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_7_i23_3_lut_LC_10_11_3 (
            .in0(N__27147),
            .in1(N__57641),
            .in2(_gnd_net_),
            .in3(N__32370),
            .lcout(n23_adj_1529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15166_2_lut_LC_10_11_4.C_ON=1'b0;
    defparam i15166_2_lut_LC_10_11_4.SEQ_MODE=4'b0000;
    defparam i15166_2_lut_LC_10_11_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 i15166_2_lut_LC_10_11_4 (
            .in0(N__57062),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49490),
            .lcout(n17564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_309_LC_10_11_5.C_ON=1'b0;
    defparam i1_2_lut_adj_309_LC_10_11_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_309_LC_10_11_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_309_LC_10_11_5 (
            .in0(_gnd_net_),
            .in1(N__55513),
            .in2(_gnd_net_),
            .in3(N__57061),
            .lcout(n12219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12096_2_lut_LC_10_11_6.C_ON=1'b0;
    defparam i12096_2_lut_LC_10_11_6.SEQ_MODE=4'b0000;
    defparam i12096_2_lut_LC_10_11_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 i12096_2_lut_LC_10_11_6 (
            .in0(N__57063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52010),
            .lcout(n14506),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15336_2_lut_3_lut_LC_10_11_7.C_ON=1'b0;
    defparam i15336_2_lut_3_lut_LC_10_11_7.SEQ_MODE=4'b0000;
    defparam i15336_2_lut_3_lut_LC_10_11_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15336_2_lut_3_lut_LC_10_11_7 (
            .in0(N__52009),
            .in1(N__45340),
            .in2(_gnd_net_),
            .in3(N__55514),
            .lcout(n14_adj_1576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i10_LC_10_12_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i10_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i10_LC_10_12_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i10_LC_10_12_0  (
            .in0(N__34612),
            .in1(N__34785),
            .in2(N__29385),
            .in3(N__31806),
            .lcout(\CLK_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i11_LC_10_12_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i11_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i11_LC_10_12_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i11_LC_10_12_1  (
            .in0(N__34780),
            .in1(N__34615),
            .in2(N__27141),
            .in3(N__43971),
            .lcout(\CLK_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i12_LC_10_12_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i12_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i12_LC_10_12_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i12_LC_10_12_2  (
            .in0(N__34613),
            .in1(N__34786),
            .in2(N__27246),
            .in3(N__40317),
            .lcout(\CLK_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i13_LC_10_12_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i13_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i13_LC_10_12_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i13_LC_10_12_3  (
            .in0(N__34781),
            .in1(N__34616),
            .in2(N__27237),
            .in3(N__27175),
            .lcout(\CLK_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i0_LC_10_12_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i0_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i0_LC_10_12_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i0_LC_10_12_4  (
            .in0(N__34611),
            .in1(N__34784),
            .in2(N__27227),
            .in3(N__33924),
            .lcout(\CLK_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i15_LC_10_12_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i15_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i15_LC_10_12_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i15_LC_10_12_5  (
            .in0(N__34782),
            .in1(N__34617),
            .in2(N__28578),
            .in3(N__27480),
            .lcout(tmp_buf_15_adj_1455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i7_LC_10_12_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i7_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i7_LC_10_12_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \CLK_DDS.tmp_buf_i7_LC_10_12_6  (
            .in0(N__34614),
            .in1(N__34787),
            .in2(N__33855),
            .in3(N__28518),
            .lcout(\CLK_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i8_LC_10_12_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i8_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i8_LC_10_12_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i8_LC_10_12_7  (
            .in0(N__34783),
            .in1(N__34618),
            .in2(N__27210),
            .in3(N__27199),
            .lcout(\CLK_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54317),
            .ce(N__34386),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_13_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_13_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i20_LC_10_13_0  (
            .in0(N__35617),
            .in1(N__35779),
            .in2(N__27558),
            .in3(N__40369),
            .lcout(buf_adcdata_iac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i13_LC_10_13_1.C_ON=1'b0;
    defparam buf_dds1_i13_LC_10_13_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i13_LC_10_13_1.LUT_INIT=16'b1100111110101010;
    LogicCell40 buf_dds1_i13_LC_10_13_1 (
            .in0(N__27176),
            .in1(N__37728),
            .in2(N__57132),
            .in3(N__44978),
            .lcout(buf_dds1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i12_LC_10_13_2.C_ON=1'b0;
    defparam buf_dds0_i12_LC_10_13_2.SEQ_MODE=4'b1000;
    defparam buf_dds0_i12_LC_10_13_2.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i12_LC_10_13_2 (
            .in0(N__56550),
            .in1(N__40339),
            .in2(N__41493),
            .in3(N__48009),
            .lcout(buf_dds0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i18_LC_10_13_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i18_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i18_LC_10_13_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i18_LC_10_13_3  (
            .in0(N__35778),
            .in1(N__35620),
            .in2(N__27320),
            .in3(N__40696),
            .lcout(buf_adcdata_iac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i7_LC_10_13_4.C_ON=1'b0;
    defparam buf_dds0_i7_LC_10_13_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i7_LC_10_13_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i7_LC_10_13_4 (
            .in0(N__56551),
            .in1(N__32321),
            .in2(N__50320),
            .in3(N__48010),
            .lcout(buf_dds0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i16_LC_10_13_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i16_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i16_LC_10_13_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i16_LC_10_13_5  (
            .in0(N__35777),
            .in1(N__35619),
            .in2(N__27375),
            .in3(N__27343),
            .lcout(buf_adcdata_iac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_13_6 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i26_LC_10_13_6  (
            .in0(N__35618),
            .in1(N__27313),
            .in2(N__28124),
            .in3(N__31963),
            .lcout(cmd_rdadctmp_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54330),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i16_3_lut_LC_10_13_7.C_ON=1'b0;
    defparam mux_129_Mux_7_i16_3_lut_LC_10_13_7.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i16_3_lut_LC_10_13_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_7_i16_3_lut_LC_10_13_7 (
            .in0(N__33848),
            .in1(N__32317),
            .in2(_gnd_net_),
            .in3(N__57739),
            .lcout(n16_adj_1504),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i16_3_lut_LC_10_14_0.C_ON=1'b0;
    defparam mux_129_Mux_5_i16_3_lut_LC_10_14_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i16_3_lut_LC_10_14_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_5_i16_3_lut_LC_10_14_0 (
            .in0(N__33884),
            .in1(N__29449),
            .in2(_gnd_net_),
            .in3(N__57665),
            .lcout(n16_adj_1496),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_252_LC_10_14_1.C_ON=1'b0;
    defparam i1_4_lut_adj_252_LC_10_14_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_252_LC_10_14_1.LUT_INIT=16'b1010000010100010;
    LogicCell40 i1_4_lut_adj_252_LC_10_14_1 (
            .in0(N__57098),
            .in1(N__41533),
            .in2(N__56549),
            .in3(N__34116),
            .lcout(n12395),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19058_2_lut_LC_10_14_2.C_ON=1'b0;
    defparam i19058_2_lut_LC_10_14_2.SEQ_MODE=4'b0000;
    defparam i19058_2_lut_LC_10_14_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19058_2_lut_LC_10_14_2 (
            .in0(_gnd_net_),
            .in1(N__57666),
            .in2(_gnd_net_),
            .in3(N__36231),
            .lcout(n21285),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i11_LC_10_14_4.C_ON=1'b0;
    defparam buf_dds0_i11_LC_10_14_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i11_LC_10_14_4.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_dds0_i11_LC_10_14_4 (
            .in0(N__43993),
            .in1(N__56488),
            .in2(N__44227),
            .in3(N__47995),
            .lcout(buf_dds0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54344),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i5_LC_10_14_5.C_ON=1'b0;
    defparam buf_dds0_i5_LC_10_14_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i5_LC_10_14_5.LUT_INIT=16'b0111001001010000;
    LogicCell40 buf_dds0_i5_LC_10_14_5 (
            .in0(N__47996),
            .in1(N__56499),
            .in2(N__29454),
            .in3(N__51437),
            .lcout(buf_dds0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54344),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_10_14_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_10_14_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i28_LC_10_14_6  (
            .in0(N__27586),
            .in1(N__28064),
            .in2(N__35598),
            .in3(N__27550),
            .lcout(cmd_rdadctmp_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54344),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i2_LC_10_14_7.C_ON=1'b0;
    defparam buf_device_acadc_i2_LC_10_14_7.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i2_LC_10_14_7.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_device_acadc_i2_LC_10_14_7 (
            .in0(N__44849),
            .in1(N__56500),
            .in2(N__40156),
            .in3(N__39787),
            .lcout(IAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54344),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19654_LC_10_15_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19654_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19654_LC_10_15_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19654_LC_10_15_0 (
            .in0(N__27534),
            .in1(N__55057),
            .in2(N__31242),
            .in3(N__53680),
            .lcout(),
            .ltout(n22279_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22279_bdd_4_lut_LC_10_15_1.C_ON=1'b0;
    defparam n22279_bdd_4_lut_LC_10_15_1.SEQ_MODE=4'b0000;
    defparam n22279_bdd_4_lut_LC_10_15_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22279_bdd_4_lut_LC_10_15_1 (
            .in0(N__53681),
            .in1(N__27459),
            .in2(N__27519),
            .in3(N__27516),
            .lcout(n22282),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19749_LC_10_15_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19749_LC_10_15_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19749_LC_10_15_2.LUT_INIT=16'b1110011010100010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19749_LC_10_15_2 (
            .in0(N__55058),
            .in1(N__53682),
            .in2(N__52671),
            .in3(N__30042),
            .lcout(),
            .ltout(n22363_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22363_bdd_4_lut_LC_10_15_3.C_ON=1'b0;
    defparam n22363_bdd_4_lut_LC_10_15_3.SEQ_MODE=4'b0000;
    defparam n22363_bdd_4_lut_LC_10_15_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22363_bdd_4_lut_LC_10_15_3 (
            .in0(N__53683),
            .in1(N__27510),
            .in2(N__27501),
            .in3(N__27498),
            .lcout(),
            .ltout(n22366_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1553158_i1_3_lut_LC_10_15_4.C_ON=1'b0;
    defparam i1553158_i1_3_lut_LC_10_15_4.SEQ_MODE=4'b0000;
    defparam i1553158_i1_3_lut_LC_10_15_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1553158_i1_3_lut_LC_10_15_4 (
            .in0(_gnd_net_),
            .in1(N__27489),
            .in2(N__27483),
            .in3(N__54719),
            .lcout(n30_adj_1531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i16_3_lut_LC_10_15_5.C_ON=1'b0;
    defparam mux_128_Mux_7_i16_3_lut_LC_10_15_5.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i16_3_lut_LC_10_15_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_7_i16_3_lut_LC_10_15_5 (
            .in0(N__27475),
            .in1(N__32074),
            .in2(_gnd_net_),
            .in3(N__57783),
            .lcout(n16_adj_1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.DTRIG_39_LC_10_15_6 .C_ON=1'b0;
    defparam \ADC_VAC.DTRIG_39_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.DTRIG_39_LC_10_15_6 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \ADC_VAC.DTRIG_39_LC_10_15_6  (
            .in0(N__30729),
            .in1(N__27453),
            .in2(N__33457),
            .in3(N__32211),
            .lcout(acadc_dtrig_v),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54358),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i9_LC_10_16_0.C_ON=1'b0;
    defparam buf_dds0_i9_LC_10_16_0.SEQ_MODE=4'b1000;
    defparam buf_dds0_i9_LC_10_16_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i9_LC_10_16_0 (
            .in0(N__56480),
            .in1(N__39727),
            .in2(N__40160),
            .in3(N__47969),
            .lcout(buf_dds0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54370),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i1_LC_10_16_1.C_ON=1'b0;
    defparam buf_device_acadc_i1_LC_10_16_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i1_LC_10_16_1.LUT_INIT=16'b0011000010111000;
    LogicCell40 buf_device_acadc_i1_LC_10_16_1 (
            .in0(N__43831),
            .in1(N__44856),
            .in2(N__27625),
            .in3(N__56484),
            .lcout(IAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54370),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i15_LC_10_16_2.C_ON=1'b0;
    defparam buf_dds0_i15_LC_10_16_2.SEQ_MODE=4'b1000;
    defparam buf_dds0_i15_LC_10_16_2.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i15_LC_10_16_2 (
            .in0(N__56479),
            .in1(N__32078),
            .in2(N__42814),
            .in3(N__47967),
            .lcout(buf_dds0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54370),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i8_LC_10_16_3.C_ON=1'b0;
    defparam buf_dds0_i8_LC_10_16_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i8_LC_10_16_3.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i8_LC_10_16_3 (
            .in0(N__47968),
            .in1(N__56482),
            .in2(N__43836),
            .in3(N__32035),
            .lcout(buf_dds0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54370),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_327_LC_10_16_4.C_ON=1'b0;
    defparam acadc_rst_327_LC_10_16_4.SEQ_MODE=4'b1000;
    defparam acadc_rst_327_LC_10_16_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_rst_327_LC_10_16_4 (
            .in0(N__44787),
            .in1(N__36254),
            .in2(_gnd_net_),
            .in3(N__40884),
            .lcout(acadc_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54370),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i4_LC_10_16_5.C_ON=1'b0;
    defparam buf_control_i4_LC_10_16_5.SEQ_MODE=4'b1000;
    defparam buf_control_i4_LC_10_16_5.LUT_INIT=16'b0011000010111000;
    LogicCell40 buf_control_i4_LC_10_16_5 (
            .in0(N__41494),
            .in1(N__41861),
            .in2(N__31849),
            .in3(N__56483),
            .lcout(VDC_RNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54370),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_247_LC_10_16_6.C_ON=1'b0;
    defparam i1_3_lut_adj_247_LC_10_16_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_247_LC_10_16_6.LUT_INIT=16'b1011101100000000;
    LogicCell40 i1_3_lut_adj_247_LC_10_16_6 (
            .in0(N__56478),
            .in1(N__30195),
            .in2(_gnd_net_),
            .in3(N__57096),
            .lcout(n12367),
            .ltout(n12367_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i1_LC_10_16_7.C_ON=1'b0;
    defparam buf_dds0_i1_LC_10_16_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i1_LC_10_16_7.LUT_INIT=16'b0010111100100000;
    LogicCell40 buf_dds0_i1_LC_10_16_7 (
            .in0(N__37448),
            .in1(N__56481),
            .in2(N__27597),
            .in3(N__32134),
            .lcout(buf_dds0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54370),
            .ce(),
            .sr(_gnd_net_));
    defparam i14145_4_lut_LC_10_17_0.C_ON=1'b0;
    defparam i14145_4_lut_LC_10_17_0.SEQ_MODE=4'b0000;
    defparam i14145_4_lut_LC_10_17_0.LUT_INIT=16'b1111000001110111;
    LogicCell40 i14145_4_lut_LC_10_17_0 (
            .in0(N__43910),
            .in1(N__30018),
            .in2(N__34041),
            .in3(N__30285),
            .lcout(),
            .ltout(n16563_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i0_LC_10_17_1.C_ON=1'b0;
    defparam eis_state_i0_LC_10_17_1.SEQ_MODE=4'b1010;
    defparam eis_state_i0_LC_10_17_1.LUT_INIT=16'b1111110000010001;
    LogicCell40 eis_state_i0_LC_10_17_1 (
            .in0(N__30286),
            .in1(N__30118),
            .in2(N__27594),
            .in3(N__27765),
            .lcout(eis_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__30075),
            .sr(N__40891));
    defparam eis_state_1__bdd_4_lut_4_lut_LC_10_17_2.C_ON=1'b0;
    defparam eis_state_1__bdd_4_lut_4_lut_LC_10_17_2.SEQ_MODE=4'b0000;
    defparam eis_state_1__bdd_4_lut_4_lut_LC_10_17_2.LUT_INIT=16'b0101100011111000;
    LogicCell40 eis_state_1__bdd_4_lut_4_lut_LC_10_17_2 (
            .in0(N__30116),
            .in1(N__30036),
            .in2(N__37300),
            .in3(N__29798),
            .lcout(n22255),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3787_3_lut_3_lut_4_lut_LC_10_17_4.C_ON=1'b0;
    defparam i3787_3_lut_3_lut_4_lut_LC_10_17_4.SEQ_MODE=4'b0000;
    defparam i3787_3_lut_3_lut_4_lut_LC_10_17_4.LUT_INIT=16'b0010000000000000;
    LogicCell40 i3787_3_lut_3_lut_4_lut_LC_10_17_4 (
            .in0(N__30117),
            .in1(N__40864),
            .in2(N__37299),
            .in3(N__29799),
            .lcout(iac_raw_buf_N_734),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19371_4_lut_LC_10_17_5.C_ON=1'b0;
    defparam i19371_4_lut_LC_10_17_5.SEQ_MODE=4'b0000;
    defparam i19371_4_lut_LC_10_17_5.LUT_INIT=16'b0000000100010001;
    LogicCell40 i19371_4_lut_LC_10_17_5 (
            .in0(N__40863),
            .in1(N__37272),
            .in2(N__30302),
            .in3(N__30114),
            .lcout(n11654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_260_LC_10_17_6.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_260_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_260_LC_10_17_6.LUT_INIT=16'b0000000000100011;
    LogicCell40 i1_3_lut_4_lut_adj_260_LC_10_17_6 (
            .in0(N__30115),
            .in1(N__30281),
            .in2(N__37298),
            .in3(N__40862),
            .lcout(n13457),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i1_LC_10_17_7.C_ON=1'b0;
    defparam eis_state_i1_LC_10_17_7.SEQ_MODE=4'b1010;
    defparam eis_state_i1_LC_10_17_7.LUT_INIT=16'b1100110011011100;
    LogicCell40 eis_state_i1_LC_10_17_7 (
            .in0(N__30127),
            .in1(N__29787),
            .in2(N__37309),
            .in3(N__30171),
            .lcout(eis_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__30075),
            .sr(N__40891));
    defparam data_index_i4_LC_10_18_0.C_ON=1'b0;
    defparam data_index_i4_LC_10_18_0.SEQ_MODE=4'b1000;
    defparam data_index_i4_LC_10_18_0.LUT_INIT=16'b0010111100100000;
    LogicCell40 data_index_i4_LC_10_18_0 (
            .in0(N__47640),
            .in1(N__56504),
            .in2(N__57144),
            .in3(N__47622),
            .lcout(data_index_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54397),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_start_329_LC_10_18_3.C_ON=1'b0;
    defparam eis_start_329_LC_10_18_3.SEQ_MODE=4'b1000;
    defparam eis_start_329_LC_10_18_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_start_329_LC_10_18_3 (
            .in0(N__43830),
            .in1(N__36258),
            .in2(_gnd_net_),
            .in3(N__43905),
            .lcout(eis_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54397),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i1_LC_10_18_4.C_ON=1'b0;
    defparam acadc_skipCount_i1_LC_10_18_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i1_LC_10_18_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i1_LC_10_18_4 (
            .in0(N__56505),
            .in1(N__44328),
            .in2(N__37455),
            .in3(N__37115),
            .lcout(acadc_skipCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54397),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_280_LC_10_18_5.C_ON=1'b0;
    defparam i1_4_lut_adj_280_LC_10_18_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_280_LC_10_18_5.LUT_INIT=16'b1011101100001011;
    LogicCell40 i1_4_lut_adj_280_LC_10_18_5 (
            .in0(N__49602),
            .in1(N__30191),
            .in2(N__56553),
            .in3(N__57139),
            .lcout(n11396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_200_LC_10_18_7.C_ON=1'b0;
    defparam i1_2_lut_adj_200_LC_10_18_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_200_LC_10_18_7.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_200_LC_10_18_7 (
            .in0(_gnd_net_),
            .in1(N__43904),
            .in2(_gnd_net_),
            .in3(N__30017),
            .lcout(n16571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19342_2_lut_LC_11_3_5 .C_ON=1'b0;
    defparam \ADC_VDC.i19342_2_lut_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19342_2_lut_LC_11_3_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ADC_VDC.i19342_2_lut_LC_11_3_5  (
            .in0(_gnd_net_),
            .in1(N__48759),
            .in2(_gnd_net_),
            .in3(N__48457),
            .lcout(\ADC_VDC.n21952 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.MISO_48_12186_12187_reset_LC_11_4_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12186_12187_reset_LC_11_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.MISO_48_12186_12187_reset_LC_11_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.MISO_48_12186_12187_reset_LC_11_4_0  (
            .in0(N__31422),
            .in1(N__30765),
            .in2(_gnd_net_),
            .in3(N__35176),
            .lcout(\comm_spi.n14605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12186_12187_resetC_net ),
            .ce(),
            .sr(N__35107));
    defparam clk_cnt_3761_3762__i1_LC_11_5_0.C_ON=1'b1;
    defparam clk_cnt_3761_3762__i1_LC_11_5_0.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i1_LC_11_5_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3761_3762__i1_LC_11_5_0 (
            .in0(_gnd_net_),
            .in1(N__30606),
            .in2(_gnd_net_),
            .in3(N__27843),
            .lcout(clk_cnt_0),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(n19746),
            .clk(N__38741),
            .ce(),
            .sr(N__30543));
    defparam clk_cnt_3761_3762__i2_LC_11_5_1.C_ON=1'b1;
    defparam clk_cnt_3761_3762__i2_LC_11_5_1.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i2_LC_11_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3761_3762__i2_LC_11_5_1 (
            .in0(_gnd_net_),
            .in1(N__30569),
            .in2(_gnd_net_),
            .in3(N__27840),
            .lcout(clk_cnt_1),
            .ltout(),
            .carryin(n19746),
            .carryout(n19747),
            .clk(N__38741),
            .ce(),
            .sr(N__30543));
    defparam clk_cnt_3761_3762__i3_LC_11_5_2.C_ON=1'b1;
    defparam clk_cnt_3761_3762__i3_LC_11_5_2.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i3_LC_11_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3761_3762__i3_LC_11_5_2 (
            .in0(_gnd_net_),
            .in1(N__30582),
            .in2(_gnd_net_),
            .in3(N__27837),
            .lcout(clk_cnt_2),
            .ltout(),
            .carryin(n19747),
            .carryout(n19748),
            .clk(N__38741),
            .ce(),
            .sr(N__30543));
    defparam clk_cnt_3761_3762__i4_LC_11_5_3.C_ON=1'b1;
    defparam clk_cnt_3761_3762__i4_LC_11_5_3.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i4_LC_11_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3761_3762__i4_LC_11_5_3 (
            .in0(_gnd_net_),
            .in1(N__30555),
            .in2(_gnd_net_),
            .in3(N__27834),
            .lcout(clk_cnt_3),
            .ltout(),
            .carryin(n19748),
            .carryout(n19749),
            .clk(N__38741),
            .ce(),
            .sr(N__30543));
    defparam clk_cnt_3761_3762__i5_LC_11_5_4.C_ON=1'b0;
    defparam clk_cnt_3761_3762__i5_LC_11_5_4.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i5_LC_11_5_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3761_3762__i5_LC_11_5_4 (
            .in0(_gnd_net_),
            .in1(N__30594),
            .in2(_gnd_net_),
            .in3(N__27831),
            .lcout(clk_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38741),
            .ce(),
            .sr(N__30543));
    defparam \comm_spi.iclk_40_12178_12179_set_LC_11_6_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12178_12179_set_LC_11_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.iclk_40_12178_12179_set_LC_11_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.iclk_40_12178_12179_set_LC_11_6_0  (
            .in0(N__27823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54272),
            .ce(),
            .sr(N__27774));
    defparam \ADC_IAC.ADC_DATA_i1_LC_11_7_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i1_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i1_LC_11_7_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_IAC.ADC_DATA_i1_LC_11_7_0  (
            .in0(N__35626),
            .in1(N__32842),
            .in2(N__35816),
            .in3(N__28155),
            .lcout(buf_adcdata_iac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i19_3_lut_LC_11_7_1.C_ON=1'b0;
    defparam mux_130_Mux_2_i19_3_lut_LC_11_7_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i19_3_lut_LC_11_7_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_2_i19_3_lut_LC_11_7_1 (
            .in0(N__28230),
            .in1(N__27886),
            .in2(_gnd_net_),
            .in3(N__57755),
            .lcout(),
            .ltout(n19_adj_1639_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i22_3_lut_LC_11_7_2.C_ON=1'b0;
    defparam mux_130_Mux_2_i22_3_lut_LC_11_7_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i22_3_lut_LC_11_7_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_2_i22_3_lut_LC_11_7_2 (
            .in0(_gnd_net_),
            .in1(N__28171),
            .in2(N__28209),
            .in3(N__53722),
            .lcout(n22_adj_1640),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i30_3_lut_LC_11_7_3.C_ON=1'b0;
    defparam mux_130_Mux_5_i30_3_lut_LC_11_7_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i30_3_lut_LC_11_7_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_5_i30_3_lut_LC_11_7_3 (
            .in0(N__28206),
            .in1(N__28194),
            .in2(_gnd_net_),
            .in3(N__54755),
            .lcout(n30_adj_1631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i2_LC_11_7_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i2_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i2_LC_11_7_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_IAC.ADC_DATA_i2_LC_11_7_4  (
            .in0(N__35627),
            .in1(N__28172),
            .in2(N__35817),
            .in3(N__28139),
            .lcout(buf_adcdata_iac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_5  (
            .in0(N__28154),
            .in1(N__28066),
            .in2(N__28140),
            .in3(N__35629),
            .lcout(cmd_rdadctmp_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_11_7_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_11_7_6 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i11_LC_11_7_6  (
            .in0(N__35628),
            .in1(N__28138),
            .in2(N__28108),
            .in3(N__28387),
            .lcout(cmd_rdadctmp_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i2_LC_11_7_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i2_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i2_LC_11_7_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_VAC.ADC_DATA_i2_LC_11_7_7  (
            .in0(N__33676),
            .in1(N__27887),
            .in2(N__33507),
            .in3(N__28347),
            .lcout(buf_adcdata_vac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54273),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i19_3_lut_LC_11_8_0.C_ON=1'b0;
    defparam mux_130_Mux_3_i19_3_lut_LC_11_8_0.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i19_3_lut_LC_11_8_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_3_i19_3_lut_LC_11_8_0 (
            .in0(N__27870),
            .in1(N__28360),
            .in2(_gnd_net_),
            .in3(N__57698),
            .lcout(n19_adj_1636),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i9_LC_11_8_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i9_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i9_LC_11_8_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i9_LC_11_8_1  (
            .in0(N__33502),
            .in1(N__33663),
            .in2(N__34933),
            .in3(N__31721),
            .lcout(buf_adcdata_vac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i2_3_lut_LC_11_8_2 .C_ON=1'b0;
    defparam \comm_spi.i2_3_lut_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i2_3_lut_LC_11_8_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \comm_spi.i2_3_lut_LC_11_8_2  (
            .in0(N__28455),
            .in1(_gnd_net_),
            .in2(N__28440),
            .in3(N__28415),
            .lcout(\comm_spi.n17036 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_8_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_8_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i3_LC_11_8_3  (
            .in0(N__35808),
            .in1(N__35630),
            .in2(N__28397),
            .in3(N__31039),
            .lcout(buf_adcdata_iac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_8_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_8_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i3_LC_11_8_4  (
            .in0(N__33662),
            .in1(N__33504),
            .in2(N__28314),
            .in3(N__28361),
            .lcout(buf_adcdata_vac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_11_8_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_11_8_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i11_LC_11_8_5  (
            .in0(N__33503),
            .in1(N__28306),
            .in2(N__28346),
            .in3(N__31691),
            .lcout(cmd_rdadctmp_11_adj_1439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_11_8_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_11_8_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i12_LC_11_8_6  (
            .in0(N__31692),
            .in1(N__28282),
            .in2(N__28313),
            .in3(N__33505),
            .lcout(cmd_rdadctmp_12_adj_1438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54277),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i30_3_lut_LC_11_8_7.C_ON=1'b0;
    defparam mux_130_Mux_2_i30_3_lut_LC_11_8_7.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i30_3_lut_LC_11_8_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_130_Mux_2_i30_3_lut_LC_11_8_7 (
            .in0(N__28260),
            .in1(N__28254),
            .in2(_gnd_net_),
            .in3(N__54756),
            .lcout(n30_adj_1641),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secclk_cnt_3765_3766__i1_LC_11_9_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i1_LC_11_9_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i1_LC_11_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i1_LC_11_9_0 (
            .in0(_gnd_net_),
            .in1(N__31107),
            .in2(_gnd_net_),
            .in3(N__28239),
            .lcout(secclk_cnt_0),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(n19750),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i2_LC_11_9_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i2_LC_11_9_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i2_LC_11_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i2_LC_11_9_1 (
            .in0(_gnd_net_),
            .in1(N__30878),
            .in2(_gnd_net_),
            .in3(N__28236),
            .lcout(secclk_cnt_1),
            .ltout(),
            .carryin(n19750),
            .carryout(n19751),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i3_LC_11_9_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i3_LC_11_9_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i3_LC_11_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i3_LC_11_9_2 (
            .in0(_gnd_net_),
            .in1(N__31214),
            .in2(_gnd_net_),
            .in3(N__28233),
            .lcout(secclk_cnt_2),
            .ltout(),
            .carryin(n19751),
            .carryout(n19752),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i4_LC_11_9_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i4_LC_11_9_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i4_LC_11_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i4_LC_11_9_3 (
            .in0(_gnd_net_),
            .in1(N__30915),
            .in2(_gnd_net_),
            .in3(N__28485),
            .lcout(secclk_cnt_3),
            .ltout(),
            .carryin(n19752),
            .carryout(n19753),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i5_LC_11_9_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i5_LC_11_9_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i5_LC_11_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i5_LC_11_9_4 (
            .in0(_gnd_net_),
            .in1(N__31068),
            .in2(_gnd_net_),
            .in3(N__28482),
            .lcout(secclk_cnt_4),
            .ltout(),
            .carryin(n19753),
            .carryout(n19754),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i6_LC_11_9_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i6_LC_11_9_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i6_LC_11_9_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i6_LC_11_9_5 (
            .in0(_gnd_net_),
            .in1(N__30864),
            .in2(_gnd_net_),
            .in3(N__28479),
            .lcout(secclk_cnt_5),
            .ltout(),
            .carryin(n19754),
            .carryout(n19755),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i7_LC_11_9_6.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i7_LC_11_9_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i7_LC_11_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i7_LC_11_9_6 (
            .in0(_gnd_net_),
            .in1(N__30954),
            .in2(_gnd_net_),
            .in3(N__28476),
            .lcout(secclk_cnt_6),
            .ltout(),
            .carryin(n19755),
            .carryout(n19756),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i8_LC_11_9_7.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i8_LC_11_9_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i8_LC_11_9_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i8_LC_11_9_7 (
            .in0(_gnd_net_),
            .in1(N__31199),
            .in2(_gnd_net_),
            .in3(N__28473),
            .lcout(secclk_cnt_7),
            .ltout(),
            .carryin(n19756),
            .carryout(n19757),
            .clk(N__38746),
            .ce(),
            .sr(N__31145));
    defparam secclk_cnt_3765_3766__i9_LC_11_10_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i9_LC_11_10_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i9_LC_11_10_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i9_LC_11_10_0 (
            .in0(_gnd_net_),
            .in1(N__30891),
            .in2(_gnd_net_),
            .in3(N__28470),
            .lcout(secclk_cnt_8),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(n19758),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i10_LC_11_10_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i10_LC_11_10_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i10_LC_11_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i10_LC_11_10_1 (
            .in0(_gnd_net_),
            .in1(N__30996),
            .in2(_gnd_net_),
            .in3(N__28467),
            .lcout(secclk_cnt_9),
            .ltout(),
            .carryin(n19758),
            .carryout(n19759),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i11_LC_11_10_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i11_LC_11_10_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i11_LC_11_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i11_LC_11_10_2 (
            .in0(_gnd_net_),
            .in1(N__30929),
            .in2(_gnd_net_),
            .in3(N__28464),
            .lcout(secclk_cnt_10),
            .ltout(),
            .carryin(n19759),
            .carryout(n19760),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i12_LC_11_10_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i12_LC_11_10_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i12_LC_11_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i12_LC_11_10_3 (
            .in0(_gnd_net_),
            .in1(N__31082),
            .in2(_gnd_net_),
            .in3(N__28461),
            .lcout(secclk_cnt_11),
            .ltout(),
            .carryin(n19760),
            .carryout(n19761),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i13_LC_11_10_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i13_LC_11_10_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i13_LC_11_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i13_LC_11_10_4 (
            .in0(_gnd_net_),
            .in1(N__31457),
            .in2(_gnd_net_),
            .in3(N__28512),
            .lcout(secclk_cnt_12),
            .ltout(),
            .carryin(n19761),
            .carryout(n19762),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i14_LC_11_10_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i14_LC_11_10_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i14_LC_11_10_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i14_LC_11_10_5 (
            .in0(_gnd_net_),
            .in1(N__31188),
            .in2(_gnd_net_),
            .in3(N__28509),
            .lcout(secclk_cnt_13),
            .ltout(),
            .carryin(n19762),
            .carryout(n19763),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i15_LC_11_10_6.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i15_LC_11_10_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i15_LC_11_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i15_LC_11_10_6 (
            .in0(_gnd_net_),
            .in1(N__30942),
            .in2(_gnd_net_),
            .in3(N__28506),
            .lcout(secclk_cnt_14),
            .ltout(),
            .carryin(n19763),
            .carryout(n19764),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i16_LC_11_10_7.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i16_LC_11_10_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i16_LC_11_10_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i16_LC_11_10_7 (
            .in0(_gnd_net_),
            .in1(N__30903),
            .in2(_gnd_net_),
            .in3(N__28503),
            .lcout(secclk_cnt_15),
            .ltout(),
            .carryin(n19764),
            .carryout(n19765),
            .clk(N__38747),
            .ce(),
            .sr(N__31138));
    defparam secclk_cnt_3765_3766__i17_LC_11_11_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i17_LC_11_11_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i17_LC_11_11_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i17_LC_11_11_0 (
            .in0(_gnd_net_),
            .in1(N__31227),
            .in2(_gnd_net_),
            .in3(N__28500),
            .lcout(secclk_cnt_16),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(n19766),
            .clk(N__38748),
            .ce(),
            .sr(N__31146));
    defparam secclk_cnt_3765_3766__i18_LC_11_11_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i18_LC_11_11_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i18_LC_11_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i18_LC_11_11_1 (
            .in0(_gnd_net_),
            .in1(N__31008),
            .in2(_gnd_net_),
            .in3(N__28497),
            .lcout(secclk_cnt_17),
            .ltout(),
            .carryin(n19766),
            .carryout(n19767),
            .clk(N__38748),
            .ce(),
            .sr(N__31146));
    defparam secclk_cnt_3765_3766__i19_LC_11_11_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i19_LC_11_11_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i19_LC_11_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i19_LC_11_11_2 (
            .in0(_gnd_net_),
            .in1(N__31095),
            .in2(_gnd_net_),
            .in3(N__28494),
            .lcout(secclk_cnt_18),
            .ltout(),
            .carryin(n19767),
            .carryout(n19768),
            .clk(N__38748),
            .ce(),
            .sr(N__31146));
    defparam secclk_cnt_3765_3766__i20_LC_11_11_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i20_LC_11_11_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i20_LC_11_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i20_LC_11_11_3 (
            .in0(_gnd_net_),
            .in1(N__31470),
            .in2(_gnd_net_),
            .in3(N__28491),
            .lcout(secclk_cnt_19),
            .ltout(),
            .carryin(n19768),
            .carryout(n19769),
            .clk(N__38748),
            .ce(),
            .sr(N__31146));
    defparam secclk_cnt_3765_3766__i21_LC_11_11_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i21_LC_11_11_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i21_LC_11_11_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i21_LC_11_11_4 (
            .in0(_gnd_net_),
            .in1(N__31158),
            .in2(_gnd_net_),
            .in3(N__28488),
            .lcout(secclk_cnt_20),
            .ltout(),
            .carryin(n19769),
            .carryout(n19770),
            .clk(N__38748),
            .ce(),
            .sr(N__31146));
    defparam secclk_cnt_3765_3766__i22_LC_11_11_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i22_LC_11_11_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i22_LC_11_11_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i22_LC_11_11_5 (
            .in0(_gnd_net_),
            .in1(N__31482),
            .in2(_gnd_net_),
            .in3(N__28620),
            .lcout(secclk_cnt_21),
            .ltout(),
            .carryin(n19770),
            .carryout(n19771),
            .clk(N__38748),
            .ce(),
            .sr(N__31146));
    defparam secclk_cnt_3765_3766__i23_LC_11_11_6.C_ON=1'b0;
    defparam secclk_cnt_3765_3766__i23_LC_11_11_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i23_LC_11_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i23_LC_11_11_6 (
            .in0(_gnd_net_),
            .in1(N__31443),
            .in2(_gnd_net_),
            .in3(N__28617),
            .lcout(secclk_cnt_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38748),
            .ce(),
            .sr(N__31146));
    defparam \CLK_DDS.tmp_buf_i14_LC_11_12_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i14_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i14_LC_11_12_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \CLK_DDS.tmp_buf_i14_LC_11_12_0  (
            .in0(N__34596),
            .in1(N__34791),
            .in2(N__28614),
            .in3(N__28584),
            .lcout(\CLK_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i1_LC_11_12_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i1_LC_11_12_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \CLK_DDS.tmp_buf_i1_LC_11_12_1  (
            .in0(N__34788),
            .in1(N__34601),
            .in2(N__33762),
            .in3(N__28569),
            .lcout(\CLK_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i2_LC_11_12_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i2_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i2_LC_11_12_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i2_LC_11_12_2  (
            .in0(N__34597),
            .in1(N__34792),
            .in2(N__28563),
            .in3(N__46893),
            .lcout(\CLK_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i3_LC_11_12_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i3_LC_11_12_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \CLK_DDS.tmp_buf_i3_LC_11_12_3  (
            .in0(N__46956),
            .in1(N__34795),
            .in2(N__28554),
            .in3(N__34602),
            .lcout(\CLK_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i4_LC_11_12_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i4_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i4_LC_11_12_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i4_LC_11_12_4  (
            .in0(N__34598),
            .in1(N__34793),
            .in2(N__28545),
            .in3(N__33999),
            .lcout(\CLK_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i5_LC_11_12_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i5_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i5_LC_11_12_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i5_LC_11_12_5  (
            .in0(N__34789),
            .in1(N__34600),
            .in2(N__28536),
            .in3(N__33885),
            .lcout(\CLK_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i6_LC_11_12_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i6_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i6_LC_11_12_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i6_LC_11_12_6  (
            .in0(N__34599),
            .in1(N__34794),
            .in2(N__28527),
            .in3(N__40761),
            .lcout(\CLK_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i9_LC_11_12_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i9_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i9_LC_11_12_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \CLK_DDS.tmp_buf_i9_LC_11_12_7  (
            .in0(N__34790),
            .in1(N__40241),
            .in2(N__34619),
            .in3(N__29391),
            .lcout(\CLK_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54305),
            .ce(N__34382),
            .sr(_gnd_net_));
    defparam data_count_i0_i0_LC_11_13_0.C_ON=1'b1;
    defparam data_count_i0_i0_LC_11_13_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i0_LC_11_13_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i0_LC_11_13_0 (
            .in0(_gnd_net_),
            .in1(N__37953),
            .in2(N__29293),
            .in3(_gnd_net_),
            .lcout(data_count_0),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(n19586),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i1_LC_11_13_1.C_ON=1'b1;
    defparam data_count_i0_i1_LC_11_13_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i1_LC_11_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i1_LC_11_13_1 (
            .in0(_gnd_net_),
            .in1(N__29179),
            .in2(_gnd_net_),
            .in3(N__29160),
            .lcout(data_count_1),
            .ltout(),
            .carryin(n19586),
            .carryout(n19587),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i2_LC_11_13_2.C_ON=1'b1;
    defparam data_count_i0_i2_LC_11_13_2.SEQ_MODE=4'b1000;
    defparam data_count_i0_i2_LC_11_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i2_LC_11_13_2 (
            .in0(_gnd_net_),
            .in1(N__29074),
            .in2(_gnd_net_),
            .in3(N__29052),
            .lcout(data_count_2),
            .ltout(),
            .carryin(n19587),
            .carryout(n19588),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i3_LC_11_13_3.C_ON=1'b1;
    defparam data_count_i0_i3_LC_11_13_3.SEQ_MODE=4'b1000;
    defparam data_count_i0_i3_LC_11_13_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i3_LC_11_13_3 (
            .in0(_gnd_net_),
            .in1(N__28969),
            .in2(_gnd_net_),
            .in3(N__28947),
            .lcout(data_count_3),
            .ltout(),
            .carryin(n19588),
            .carryout(n19589),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i4_LC_11_13_4.C_ON=1'b1;
    defparam data_count_i0_i4_LC_11_13_4.SEQ_MODE=4'b1000;
    defparam data_count_i0_i4_LC_11_13_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i4_LC_11_13_4 (
            .in0(_gnd_net_),
            .in1(N__28858),
            .in2(_gnd_net_),
            .in3(N__28836),
            .lcout(data_count_4),
            .ltout(),
            .carryin(n19589),
            .carryout(n19590),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i5_LC_11_13_5.C_ON=1'b1;
    defparam data_count_i0_i5_LC_11_13_5.SEQ_MODE=4'b1000;
    defparam data_count_i0_i5_LC_11_13_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i5_LC_11_13_5 (
            .in0(_gnd_net_),
            .in1(N__28753),
            .in2(_gnd_net_),
            .in3(N__28728),
            .lcout(data_count_5),
            .ltout(),
            .carryin(n19590),
            .carryout(n19591),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i6_LC_11_13_6.C_ON=1'b1;
    defparam data_count_i0_i6_LC_11_13_6.SEQ_MODE=4'b1000;
    defparam data_count_i0_i6_LC_11_13_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i6_LC_11_13_6 (
            .in0(_gnd_net_),
            .in1(N__28645),
            .in2(_gnd_net_),
            .in3(N__28623),
            .lcout(data_count_6),
            .ltout(),
            .carryin(n19591),
            .carryout(n19592),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i7_LC_11_13_7.C_ON=1'b1;
    defparam data_count_i0_i7_LC_11_13_7.SEQ_MODE=4'b1000;
    defparam data_count_i0_i7_LC_11_13_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i7_LC_11_13_7 (
            .in0(_gnd_net_),
            .in1(N__29701),
            .in2(_gnd_net_),
            .in3(N__29682),
            .lcout(data_count_7),
            .ltout(),
            .carryin(n19592),
            .carryout(n19593),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38558),
            .sr(N__38482));
    defparam data_count_i0_i8_LC_11_14_0.C_ON=1'b1;
    defparam data_count_i0_i8_LC_11_14_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i8_LC_11_14_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i8_LC_11_14_0 (
            .in0(_gnd_net_),
            .in1(N__29593),
            .in2(_gnd_net_),
            .in3(N__29574),
            .lcout(data_count_8),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(n19594),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__38552),
            .sr(N__38496));
    defparam data_count_i0_i9_LC_11_14_1.C_ON=1'b0;
    defparam data_count_i0_i9_LC_11_14_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i9_LC_11_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i9_LC_11_14_1 (
            .in0(_gnd_net_),
            .in1(N__29482),
            .in2(_gnd_net_),
            .in3(N__29571),
            .lcout(data_count_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__38552),
            .sr(N__38496));
    defparam \SIG_DDS.tmp_buf_i10_LC_11_15_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i10_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i10_LC_11_15_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i10_LC_11_15_0  (
            .in0(N__42268),
            .in1(N__43066),
            .in2(N__29817),
            .in3(N__40980),
            .lcout(\SIG_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i11_LC_11_15_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i11_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i11_LC_11_15_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i11_LC_11_15_1  (
            .in0(N__43062),
            .in1(N__42272),
            .in2(N__29463),
            .in3(N__44000),
            .lcout(\SIG_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i5_LC_11_15_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i5_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i5_LC_11_15_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i5_LC_11_15_2  (
            .in0(N__42270),
            .in1(N__43068),
            .in2(N__32052),
            .in3(N__29453),
            .lcout(\SIG_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i13_LC_11_15_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i13_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i13_LC_11_15_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i13_LC_11_15_3  (
            .in0(N__43064),
            .in1(N__42274),
            .in2(N__29400),
            .in3(N__41631),
            .lcout(\SIG_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i14_LC_11_15_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i14_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i14_LC_11_15_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \SIG_DDS.tmp_buf_i14_LC_11_15_4  (
            .in0(N__42269),
            .in1(N__43067),
            .in2(N__29436),
            .in3(N__29415),
            .lcout(\SIG_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i12_LC_11_15_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i12_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i12_LC_11_15_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i12_LC_11_15_5  (
            .in0(N__43063),
            .in1(N__42273),
            .in2(N__29409),
            .in3(N__40346),
            .lcout(\SIG_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i9_LC_11_15_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i9_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i9_LC_11_15_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i9_LC_11_15_6  (
            .in0(N__42271),
            .in1(N__43069),
            .in2(N__32013),
            .in3(N__39728),
            .lcout(\SIG_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i6_LC_11_15_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i6_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i6_LC_11_15_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i6_LC_11_15_7  (
            .in0(N__43065),
            .in1(N__42275),
            .in2(N__29808),
            .in3(N__40734),
            .lcout(\SIG_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54345),
            .ce(N__42090),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_217_LC_11_16_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_217_LC_11_16_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_217_LC_11_16_0.LUT_INIT=16'b0010001000000000;
    LogicCell40 i1_2_lut_3_lut_adj_217_LC_11_16_0 (
            .in0(N__32177),
            .in1(N__30296),
            .in2(_gnd_net_),
            .in3(N__32207),
            .lcout(n16554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_168_LC_11_16_1.C_ON=1'b0;
    defparam i5_4_lut_adj_168_LC_11_16_1.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_168_LC_11_16_1.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_adj_168_LC_11_16_1 (
            .in0(N__32439),
            .in1(N__32478),
            .in2(N__32274),
            .in3(N__32290),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_238_LC_11_16_2.C_ON=1'b0;
    defparam i1_4_lut_adj_238_LC_11_16_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_238_LC_11_16_2.LUT_INIT=16'b1000100010001100;
    LogicCell40 i1_4_lut_adj_238_LC_11_16_2 (
            .in0(N__56519),
            .in1(N__57097),
            .in2(N__33111),
            .in3(N__41778),
            .lcout(n11915),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_LC_11_16_3 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_LC_11_16_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ADC_VAC.i1_2_lut_LC_11_16_3  (
            .in0(N__32206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32176),
            .lcout(iac_raw_buf_N_736),
            .ltout(iac_raw_buf_N_736_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_11_16_4.C_ON=1'b0;
    defparam i24_4_lut_LC_11_16_4.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_11_16_4.LUT_INIT=16'b0110011011100100;
    LogicCell40 i24_4_lut_LC_11_16_4 (
            .in0(N__30306),
            .in1(N__30122),
            .in2(N__29790),
            .in3(N__37292),
            .lcout(n17_adj_1622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19331_4_lut_LC_11_16_5.C_ON=1'b0;
    defparam i19331_4_lut_LC_11_16_5.SEQ_MODE=4'b0000;
    defparam i19331_4_lut_LC_11_16_5.LUT_INIT=16'b0001101100010011;
    LogicCell40 i19331_4_lut_LC_11_16_5 (
            .in0(N__37293),
            .in1(N__30307),
            .in2(N__30135),
            .in3(N__32151),
            .lcout(),
            .ltout(n20826_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_end_299_LC_11_16_6.C_ON=1'b0;
    defparam eis_end_299_LC_11_16_6.SEQ_MODE=4'b1000;
    defparam eis_end_299_LC_11_16_6.LUT_INIT=16'b1010101011001010;
    LogicCell40 eis_end_299_LC_11_16_6 (
            .in0(N__30051),
            .in1(N__30297),
            .in2(N__29781),
            .in3(N__40877),
            .lcout(eis_end),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_end_299C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i26_3_lut_LC_11_16_7.C_ON=1'b0;
    defparam mux_128_Mux_7_i26_3_lut_LC_11_16_7.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i26_3_lut_LC_11_16_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_128_Mux_7_i26_3_lut_LC_11_16_7 (
            .in0(N__38004),
            .in1(N__57823),
            .in2(_gnd_net_),
            .in3(N__30050),
            .lcout(n26_adj_1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18989_2_lut_3_lut_LC_11_17_0.C_ON=1'b0;
    defparam i18989_2_lut_3_lut_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam i18989_2_lut_3_lut_LC_11_17_0.LUT_INIT=16'b0010001010101010;
    LogicCell40 i18989_2_lut_3_lut_LC_11_17_0 (
            .in0(N__30295),
            .in1(N__32213),
            .in2(_gnd_net_),
            .in3(N__32174),
            .lcout(n21234),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_11_17_1.C_ON=1'b0;
    defparam i14_4_lut_LC_11_17_1.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_11_17_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_LC_11_17_1 (
            .in0(N__32376),
            .in1(N__41565),
            .in2(N__30030),
            .in3(N__32382),
            .lcout(),
            .ltout(n30_adj_1604_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_LC_11_17_2.C_ON=1'b0;
    defparam i15_4_lut_LC_11_17_2.SEQ_MODE=4'b0000;
    defparam i15_4_lut_LC_11_17_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_LC_11_17_2 (
            .in0(N__29823),
            .in1(N__38412),
            .in2(N__30021),
            .in3(N__29829),
            .lcout(n31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.DTRIG_39_LC_11_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.DTRIG_39_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.DTRIG_39_LC_11_17_3 .LUT_INIT=16'b1011101010101000;
    LogicCell40 \ADC_IAC.DTRIG_39_LC_11_17_3  (
            .in0(N__32175),
            .in1(N__35569),
            .in2(N__30006),
            .in3(N__29912),
            .lcout(acadc_dtrig_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54371),
            .ce(),
            .sr(_gnd_net_));
    defparam i15109_2_lut_LC_11_17_4.C_ON=1'b0;
    defparam i15109_2_lut_LC_11_17_4.SEQ_MODE=4'b0000;
    defparam i15109_2_lut_LC_11_17_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i15109_2_lut_LC_11_17_4 (
            .in0(_gnd_net_),
            .in1(N__32212),
            .in2(_gnd_net_),
            .in3(N__32173),
            .lcout(n17507),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_61_i14_2_lut_LC_11_17_5.C_ON=1'b0;
    defparam equal_61_i14_2_lut_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam equal_61_i14_2_lut_LC_11_17_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 equal_61_i14_2_lut_LC_11_17_5 (
            .in0(_gnd_net_),
            .in1(N__32715),
            .in2(_gnd_net_),
            .in3(N__32239),
            .lcout(),
            .ltout(n14_adj_1509_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_11_17_6.C_ON=1'b0;
    defparam i10_4_lut_LC_11_17_6.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_11_17_6.LUT_INIT=16'b1111111111110110;
    LogicCell40 i10_4_lut_LC_11_17_6 (
            .in0(N__32514),
            .in1(N__43639),
            .in2(N__29832),
            .in3(N__32223),
            .lcout(n26_adj_1508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_170_LC_11_18_0.C_ON=1'b0;
    defparam i2_4_lut_adj_170_LC_11_18_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_170_LC_11_18_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_170_LC_11_18_0 (
            .in0(N__32417),
            .in1(N__46837),
            .in2(N__32556),
            .in3(N__37111),
            .lcout(n18_adj_1609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i4_LC_11_18_2.C_ON=1'b0;
    defparam acadc_skipCount_i4_LC_11_18_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i4_LC_11_18_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i4_LC_11_18_2 (
            .in0(N__56546),
            .in1(N__44327),
            .in2(N__47801),
            .in3(N__46838),
            .lcout(acadc_skipCount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54385),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_11_18_3.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_11_18_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_11_18_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_4_lut_LC_11_18_3 (
            .in0(N__55208),
            .in1(N__57782),
            .in2(N__41540),
            .in3(N__53721),
            .lcout(n20915),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18376_4_lut_LC_11_18_5.C_ON=1'b0;
    defparam i18376_4_lut_LC_11_18_5.SEQ_MODE=4'b0000;
    defparam i18376_4_lut_LC_11_18_5.LUT_INIT=16'b1111111110111000;
    LogicCell40 i18376_4_lut_LC_11_18_5 (
            .in0(N__30126),
            .in1(N__37291),
            .in2(N__30298),
            .in3(N__40885),
            .lcout(n20985),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i11_LC_11_18_6.C_ON=1'b0;
    defparam acadc_skipCount_i11_LC_11_18_6.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i11_LC_11_18_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i11_LC_11_18_6 (
            .in0(N__56545),
            .in1(N__44326),
            .in2(N__44226),
            .in3(N__41926),
            .lcout(acadc_skipCount_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54385),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i2_LC_11_18_7.C_ON=1'b0;
    defparam buf_control_i2_LC_11_18_7.SEQ_MODE=4'b1000;
    defparam buf_control_i2_LC_11_18_7.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_control_i2_LC_11_18_7 (
            .in0(N__41874),
            .in1(N__56547),
            .in2(N__44788),
            .in3(N__31765),
            .lcout(SELIRNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54385),
            .ce(),
            .sr(_gnd_net_));
    defparam i19109_2_lut_LC_11_19_0.C_ON=1'b0;
    defparam i19109_2_lut_LC_11_19_0.SEQ_MODE=4'b0000;
    defparam i19109_2_lut_LC_11_19_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19109_2_lut_LC_11_19_0 (
            .in0(_gnd_net_),
            .in1(N__30139),
            .in2(_gnd_net_),
            .in3(N__34037),
            .lcout(n21337),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i34_3_lut_LC_11_19_1.C_ON=1'b0;
    defparam i34_3_lut_LC_11_19_1.SEQ_MODE=4'b0000;
    defparam i34_3_lut_LC_11_19_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i34_3_lut_LC_11_19_1 (
            .in0(N__30140),
            .in1(N__37958),
            .in2(_gnd_net_),
            .in3(N__30170),
            .lcout(),
            .ltout(n13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i2_LC_11_19_2.C_ON=1'b0;
    defparam eis_state_i2_LC_11_19_2.SEQ_MODE=4'b1010;
    defparam eis_state_i2_LC_11_19_2.LUT_INIT=16'b1110110001100100;
    LogicCell40 eis_state_i2_LC_11_19_2 (
            .in0(N__37308),
            .in1(N__30274),
            .in2(N__30159),
            .in3(N__30156),
            .lcout(eis_end_N_724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i2C_net),
            .ce(N__30074),
            .sr(N__40889));
    defparam i24_4_lut_adj_188_LC_11_19_3.C_ON=1'b0;
    defparam i24_4_lut_adj_188_LC_11_19_3.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_188_LC_11_19_3.LUT_INIT=16'b1111110010101100;
    LogicCell40 i24_4_lut_adj_188_LC_11_19_3 (
            .in0(N__43906),
            .in1(N__30150),
            .in2(N__30141),
            .in3(N__34296),
            .lcout(),
            .ltout(n11_adj_1621_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19384_3_lut_LC_11_19_4.C_ON=1'b0;
    defparam i19384_3_lut_LC_11_19_4.SEQ_MODE=4'b0000;
    defparam i19384_3_lut_LC_11_19_4.LUT_INIT=16'b0011111111111111;
    LogicCell40 i19384_3_lut_LC_11_19_4 (
            .in0(_gnd_net_),
            .in1(N__37307),
            .in2(N__30078),
            .in3(N__30273),
            .lcout(n11744),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19350_2_lut_LC_11_20_7.C_ON=1'b0;
    defparam i19350_2_lut_LC_11_20_7.SEQ_MODE=4'b0000;
    defparam i19350_2_lut_LC_11_20_7.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19350_2_lut_LC_11_20_7 (
            .in0(_gnd_net_),
            .in1(N__30272),
            .in2(_gnd_net_),
            .in3(N__32646),
            .lcout(n14671),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7704_3_lut_4_lut_LC_12_3_1 .C_ON=1'b0;
    defparam \ADC_VDC.i7704_3_lut_4_lut_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7704_3_lut_4_lut_LC_12_3_1 .LUT_INIT=16'b0011010010111100;
    LogicCell40 \ADC_VDC.i7704_3_lut_4_lut_LC_12_3_1  (
            .in0(N__48299),
            .in1(N__47361),
            .in2(N__47490),
            .in3(N__34830),
            .lcout(),
            .ltout(\ADC_VDC.n10119_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_12_3_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_12_3_2 .LUT_INIT=16'b1011101011111110;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_LC_12_3_2  (
            .in0(N__48760),
            .in1(N__48465),
            .in2(N__30213),
            .in3(N__32568),
            .lcout(\ADC_VDC.n12807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i3_LC_12_3_3 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i3_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i3_LC_12_3_3 .LUT_INIT=16'b0100001000001010;
    LogicCell40 \ADC_VDC.adc_state_i3_LC_12_3_3  (
            .in0(N__48466),
            .in1(N__48279),
            .in2(N__48772),
            .in3(N__47362),
            .lcout(adc_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53298),
            .ce(N__30210),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16150_3_lut_LC_12_3_5 .C_ON=1'b0;
    defparam \ADC_VDC.i16150_3_lut_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16150_3_lut_LC_12_3_5 .LUT_INIT=16'b1101110110101010;
    LogicCell40 \ADC_VDC.i16150_3_lut_LC_12_3_5  (
            .in0(N__47473),
            .in1(N__48278),
            .in2(_gnd_net_),
            .in3(N__47360),
            .lcout(\ADC_VDC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_10_LC_12_3_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_10_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_10_LC_12_3_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_10_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__48689),
            .in2(_gnd_net_),
            .in3(N__48464),
            .lcout(\ADC_VDC.n20899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i0_LC_12_4_0.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i0_LC_12_4_0.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i0_LC_12_4_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i0_LC_12_4_0 (
            .in0(_gnd_net_),
            .in1(N__30801),
            .in2(_gnd_net_),
            .in3(N__30204),
            .lcout(dds0_mclkcnt_0),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(n19739),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i1_LC_12_4_1.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i1_LC_12_4_1.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i1_LC_12_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i1_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(N__30839),
            .in2(_gnd_net_),
            .in3(N__30201),
            .lcout(dds0_mclkcnt_1),
            .ltout(),
            .carryin(n19739),
            .carryout(n19740),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i2_LC_12_4_2.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i2_LC_12_4_2.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i2_LC_12_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i2_LC_12_4_2 (
            .in0(_gnd_net_),
            .in1(N__30813),
            .in2(_gnd_net_),
            .in3(N__30198),
            .lcout(dds0_mclkcnt_2),
            .ltout(),
            .carryin(n19740),
            .carryout(n19741),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i3_LC_12_4_3.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i3_LC_12_4_3.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i3_LC_12_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i3_LC_12_4_3 (
            .in0(_gnd_net_),
            .in1(N__30321),
            .in2(_gnd_net_),
            .in3(N__30621),
            .lcout(dds0_mclkcnt_3),
            .ltout(),
            .carryin(n19741),
            .carryout(n19742),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i4_LC_12_4_4.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i4_LC_12_4_4.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i4_LC_12_4_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i4_LC_12_4_4 (
            .in0(_gnd_net_),
            .in1(N__30825),
            .in2(_gnd_net_),
            .in3(N__30618),
            .lcout(dds0_mclkcnt_4),
            .ltout(),
            .carryin(n19742),
            .carryout(n19743),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i5_LC_12_4_5.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i5_LC_12_4_5.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i5_LC_12_4_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i5_LC_12_4_5 (
            .in0(_gnd_net_),
            .in1(N__30852),
            .in2(_gnd_net_),
            .in3(N__30615),
            .lcout(dds0_mclkcnt_5),
            .ltout(),
            .carryin(n19743),
            .carryout(n19744),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i6_LC_12_4_6.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i6_LC_12_4_6.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i6_LC_12_4_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i6_LC_12_4_6 (
            .in0(_gnd_net_),
            .in1(N__30771),
            .in2(_gnd_net_),
            .in3(N__30612),
            .lcout(dds0_mclkcnt_6),
            .ltout(),
            .carryin(n19744),
            .carryout(n19745),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i7_LC_12_4_7.C_ON=1'b0;
    defparam dds0_mclkcnt_i7_3772__i7_LC_12_4_7.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i7_LC_12_4_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i7_LC_12_4_7 (
            .in0(_gnd_net_),
            .in1(N__30786),
            .in2(_gnd_net_),
            .in3(N__30609),
            .lcout(dds0_mclkcnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_250_LC_12_5_0.C_ON=1'b0;
    defparam i1_2_lut_adj_250_LC_12_5_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_250_LC_12_5_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_adj_250_LC_12_5_0 (
            .in0(N__30605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30593),
            .lcout(),
            .ltout(n6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_253_LC_12_5_1.C_ON=1'b0;
    defparam i4_4_lut_adj_253_LC_12_5_1.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_253_LC_12_5_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i4_4_lut_adj_253_LC_12_5_1 (
            .in0(N__30581),
            .in1(N__30570),
            .in2(N__30558),
            .in3(N__30554),
            .lcout(n14714),
            .ltout(n14714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_RTD_287_LC_12_5_2.C_ON=1'b0;
    defparam clk_RTD_287_LC_12_5_2.SEQ_MODE=4'b1000;
    defparam clk_RTD_287_LC_12_5_2.LUT_INIT=16'b0000111111110000;
    LogicCell40 clk_RTD_287_LC_12_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30531),
            .in3(N__30346),
            .lcout(clk_RTD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38740),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_12_5_3.C_ON=1'b0;
    defparam i5_4_lut_LC_12_5_3.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_12_5_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_LC_12_5_3 (
            .in0(N__30320),
            .in1(N__30851),
            .in2(N__30840),
            .in3(N__30824),
            .lcout(),
            .ltout(n12_adj_1480_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_12_5_4.C_ON=1'b0;
    defparam i6_4_lut_LC_12_5_4.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_12_5_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_12_5_4 (
            .in0(N__30812),
            .in1(N__30800),
            .in2(N__30789),
            .in3(N__30785),
            .lcout(n20799),
            .ltout(n20799_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15251_2_lut_LC_12_5_5.C_ON=1'b0;
    defparam i15251_2_lut_LC_12_5_5.SEQ_MODE=4'b0000;
    defparam i15251_2_lut_LC_12_5_5.LUT_INIT=16'b1111000000000000;
    LogicCell40 i15251_2_lut_LC_12_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30774),
            .in3(N__30974),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imiso_83_12192_12193_reset_LC_12_6_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12192_12193_reset_LC_12_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imiso_83_12192_12193_reset_LC_12_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.imiso_83_12192_12193_reset_LC_12_6_0  (
            .in0(N__35178),
            .in1(N__34352),
            .in2(_gnd_net_),
            .in3(N__32882),
            .lcout(\comm_spi.n14611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12192_12193_resetC_net ),
            .ce(),
            .sr(N__35109));
    defparam \comm_spi.MISO_48_12186_12187_set_LC_12_7_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12186_12187_set_LC_12_7_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.MISO_48_12186_12187_set_LC_12_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.MISO_48_12186_12187_set_LC_12_7_0  (
            .in0(N__31418),
            .in1(N__30761),
            .in2(_gnd_net_),
            .in3(N__35172),
            .lcout(\comm_spi.n14604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12186_12187_setC_net ),
            .ce(),
            .sr(N__35045));
    defparam \ADC_VAC.i12431_2_lut_LC_12_7_5 .C_ON=1'b0;
    defparam \ADC_VAC.i12431_2_lut_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i12431_2_lut_LC_12_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ADC_VAC.i12431_2_lut_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__30750),
            .in2(_gnd_net_),
            .in3(N__30728),
            .lcout(\ADC_VAC.n14844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_12_7_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_12_7_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_89_2_lut_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__55637),
            .in2(_gnd_net_),
            .in3(N__55777),
            .lcout(\comm_spi.imosi_N_753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i7_LC_12_8_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i7_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i7_LC_12_8_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i7_LC_12_8_0  (
            .in0(N__35894),
            .in1(N__46404),
            .in2(_gnd_net_),
            .in3(N__35846),
            .lcout(comm_rx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(),
            .sr(N__55869));
    defparam \comm_spi.data_rx_i6_LC_12_8_1 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i6_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i6_LC_12_8_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i6_LC_12_8_1  (
            .in0(N__35845),
            .in1(N__52058),
            .in2(_gnd_net_),
            .in3(N__35893),
            .lcout(comm_rx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(),
            .sr(N__55869));
    defparam \comm_spi.data_rx_i5_LC_12_8_2 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i5_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i5_LC_12_8_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i5_LC_12_8_2  (
            .in0(N__35892),
            .in1(N__46715),
            .in2(_gnd_net_),
            .in3(N__35844),
            .lcout(comm_rx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(),
            .sr(N__55869));
    defparam \comm_spi.data_rx_i4_LC_12_8_3 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i4_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i4_LC_12_8_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i4_LC_12_8_3  (
            .in0(N__35843),
            .in1(N__51054),
            .in2(_gnd_net_),
            .in3(N__35891),
            .lcout(comm_rx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(),
            .sr(N__55869));
    defparam \comm_spi.data_rx_i3_LC_12_8_4 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i3_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i3_LC_12_8_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i3_LC_12_8_4  (
            .in0(N__35890),
            .in1(N__47174),
            .in2(_gnd_net_),
            .in3(N__35842),
            .lcout(comm_rx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(),
            .sr(N__55869));
    defparam \comm_spi.data_rx_i2_LC_12_8_5 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i2_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i2_LC_12_8_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i2_LC_12_8_5  (
            .in0(N__35841),
            .in1(N__45724),
            .in2(_gnd_net_),
            .in3(N__35889),
            .lcout(comm_rx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(),
            .sr(N__55869));
    defparam \comm_spi.data_rx_i1_LC_12_8_6 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i1_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i1_LC_12_8_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \comm_spi.data_rx_i1_LC_12_8_6  (
            .in0(N__35888),
            .in1(N__35840),
            .in2(_gnd_net_),
            .in3(N__53050),
            .lcout(comm_rx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(),
            .sr(N__55869));
    defparam dds0_mclk_294_LC_12_9_0.C_ON=1'b0;
    defparam dds0_mclk_294_LC_12_9_0.SEQ_MODE=4'b1000;
    defparam dds0_mclk_294_LC_12_9_0.LUT_INIT=16'b1010101001100110;
    LogicCell40 dds0_mclk_294_LC_12_9_0 (
            .in0(N__38690),
            .in1(N__30978),
            .in2(_gnd_net_),
            .in3(N__30963),
            .lcout(dds0_mclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclk_294C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i4_4_lut_LC_12_9_1 .C_ON=1'b0;
    defparam \SIG_DDS.i4_4_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i4_4_lut_LC_12_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \SIG_DDS.i4_4_lut_LC_12_9_1  (
            .in0(N__43134),
            .in1(N__43150),
            .in2(N__43098),
            .in3(N__41301),
            .lcout(\SIG_DDS.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_196_LC_12_9_4.C_ON=1'b0;
    defparam i11_4_lut_adj_196_LC_12_9_4.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_196_LC_12_9_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_196_LC_12_9_4 (
            .in0(N__30953),
            .in1(N__30941),
            .in2(N__30930),
            .in3(N__30914),
            .lcout(n27_adj_1597),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_12_9_5.C_ON=1'b0;
    defparam i9_4_lut_LC_12_9_5.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_12_9_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_12_9_5 (
            .in0(N__30902),
            .in1(N__30890),
            .in2(N__30879),
            .in3(N__30863),
            .lcout(n25_adj_1574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_193_LC_12_10_0.C_ON=1'b0;
    defparam i10_4_lut_adj_193_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_193_LC_12_10_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_193_LC_12_10_0 (
            .in0(N__31226),
            .in1(N__31215),
            .in2(N__31203),
            .in3(N__31187),
            .lcout(),
            .ltout(n26_adj_1575_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_205_LC_12_10_1.C_ON=1'b0;
    defparam i15_4_lut_adj_205_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_205_LC_12_10_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_205_LC_12_10_1 (
            .in0(N__31056),
            .in1(N__31176),
            .in2(N__31170),
            .in3(N__31167),
            .lcout(),
            .ltout(n19856_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_206_LC_12_10_2.C_ON=1'b0;
    defparam i7_4_lut_adj_206_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_206_LC_12_10_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 i7_4_lut_adj_206_LC_12_10_2 (
            .in0(N__31431),
            .in1(N__30984),
            .in2(N__31161),
            .in3(N__31157),
            .lcout(n14715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_189_LC_12_10_3.C_ON=1'b0;
    defparam i12_4_lut_adj_189_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_189_LC_12_10_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_189_LC_12_10_3 (
            .in0(N__31106),
            .in1(N__31094),
            .in2(N__31083),
            .in3(N__31067),
            .lcout(n28_adj_1505),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i0_LC_12_10_4 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i0_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i0_LC_12_10_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \SIG_DDS.bit_cnt_i0_LC_12_10_4  (
            .in0(N__43157),
            .in1(N__43061),
            .in2(_gnd_net_),
            .in3(N__42881),
            .lcout(bit_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54280),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i22_3_lut_LC_12_10_6.C_ON=1'b0;
    defparam mux_130_Mux_3_i22_3_lut_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i22_3_lut_LC_12_10_6.LUT_INIT=16'b1100101011001010;
    LogicCell40 mux_130_Mux_3_i22_3_lut_LC_12_10_6 (
            .in0(N__31040),
            .in1(N__31017),
            .in2(N__53795),
            .in3(_gnd_net_),
            .lcout(n22_adj_1637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_12_11_0.C_ON=1'b0;
    defparam i2_2_lut_LC_12_11_0.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_12_11_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2_2_lut_LC_12_11_0 (
            .in0(_gnd_net_),
            .in1(N__31007),
            .in2(_gnd_net_),
            .in3(N__30995),
            .lcout(n10_adj_1601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_11_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_96_2_lut_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__34902),
            .in2(_gnd_net_),
            .in3(N__55866),
            .lcout(\comm_spi.data_tx_7__N_770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i30_3_lut_LC_12_11_2.C_ON=1'b0;
    defparam mux_130_Mux_3_i30_3_lut_LC_12_11_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i30_3_lut_LC_12_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_3_i30_3_lut_LC_12_11_2 (
            .in0(N__31746),
            .in1(N__31728),
            .in2(_gnd_net_),
            .in3(N__54644),
            .lcout(n30_adj_1638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_12_11_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_12_11_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i18_LC_12_11_4  (
            .in0(N__31722),
            .in1(N__33494),
            .in2(N__33129),
            .in3(N__31689),
            .lcout(cmd_rdadctmp_18_adj_1432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54286),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_12_11_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_12_11_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i19_LC_12_11_5  (
            .in0(N__31690),
            .in1(N__31498),
            .in2(N__33506),
            .in3(N__33127),
            .lcout(cmd_rdadctmp_19_adj_1431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54286),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_197_LC_12_11_7.C_ON=1'b0;
    defparam i6_4_lut_adj_197_LC_12_11_7.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_197_LC_12_11_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_adj_197_LC_12_11_7 (
            .in0(N__31481),
            .in1(N__31469),
            .in2(N__31458),
            .in3(N__31442),
            .lcout(n14_adj_1599),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imiso_83_12192_12193_set_LC_12_12_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12192_12193_set_LC_12_12_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imiso_83_12192_12193_set_LC_12_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.imiso_83_12192_12193_set_LC_12_12_0  (
            .in0(N__35177),
            .in1(N__34359),
            .in2(_gnd_net_),
            .in3(N__32889),
            .lcout(\comm_spi.n14610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12192_12193_setC_net ),
            .ce(),
            .sr(N__35049));
    defparam mux_128_Mux_6_i20_3_lut_LC_12_12_2.C_ON=1'b0;
    defparam mux_128_Mux_6_i20_3_lut_LC_12_12_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_6_i20_3_lut_LC_12_12_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_6_i20_3_lut_LC_12_12_2 (
            .in0(N__31404),
            .in1(N__31371),
            .in2(_gnd_net_),
            .in3(N__57383),
            .lcout(n20_adj_1537),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i20_3_lut_LC_12_12_4.C_ON=1'b0;
    defparam mux_128_Mux_7_i20_3_lut_LC_12_12_4.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i20_3_lut_LC_12_12_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_7_i20_3_lut_LC_12_12_4 (
            .in0(N__31323),
            .in1(N__31287),
            .in2(_gnd_net_),
            .in3(N__57381),
            .lcout(n20_adj_1528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_0_i16_3_lut_LC_12_12_5.C_ON=1'b0;
    defparam mux_129_Mux_0_i16_3_lut_LC_12_12_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i16_3_lut_LC_12_12_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_0_i16_3_lut_LC_12_12_5 (
            .in0(N__57382),
            .in1(N__33919),
            .in2(_gnd_net_),
            .in3(N__33968),
            .lcout(n16_adj_1487),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i16_3_lut_LC_12_12_6.C_ON=1'b0;
    defparam mux_129_Mux_1_i16_3_lut_LC_12_12_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i16_3_lut_LC_12_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_1_i16_3_lut_LC_12_12_6 (
            .in0(N__33754),
            .in1(N__32145),
            .in2(_gnd_net_),
            .in3(N__57384),
            .lcout(n16_adj_1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i11_LC_12_13_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i11_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i11_LC_12_13_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_IAC.ADC_DATA_i11_LC_12_13_0  (
            .in0(N__35803),
            .in1(N__52774),
            .in2(N__32001),
            .in3(N__35623),
            .lcout(buf_adcdata_iac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i17_LC_12_13_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i17_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i17_LC_12_13_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i17_LC_12_13_1  (
            .in0(N__35622),
            .in1(N__35804),
            .in2(N__31968),
            .in3(N__39754),
            .lcout(buf_adcdata_iac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i13_LC_12_13_2.C_ON=1'b0;
    defparam req_data_cnt_i13_LC_12_13_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i13_LC_12_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i13_LC_12_13_2 (
            .in0(N__37717),
            .in1(N__41742),
            .in2(_gnd_net_),
            .in3(N__33944),
            .lcout(req_data_cnt_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_6_i17_3_lut_LC_12_13_4.C_ON=1'b0;
    defparam mux_128_Mux_6_i17_3_lut_LC_12_13_4.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_6_i17_3_lut_LC_12_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_6_i17_3_lut_LC_12_13_4 (
            .in0(N__57591),
            .in1(N__31937),
            .in2(_gnd_net_),
            .in3(N__31895),
            .lcout(n17_adj_1535),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i10_LC_12_13_5.C_ON=1'b0;
    defparam buf_dds1_i10_LC_12_13_5.SEQ_MODE=4'b1000;
    defparam buf_dds1_i10_LC_12_13_5.LUT_INIT=16'b1100000010001000;
    LogicCell40 buf_dds1_i10_LC_12_13_5 (
            .in0(N__31802),
            .in1(N__40667),
            .in2(N__44792),
            .in3(N__44957),
            .lcout(buf_dds1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54300),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_4_i23_3_lut_LC_12_13_6.C_ON=1'b0;
    defparam mux_128_Mux_4_i23_3_lut_LC_12_13_6.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_4_i23_3_lut_LC_12_13_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_128_Mux_4_i23_3_lut_LC_12_13_6 (
            .in0(N__57590),
            .in1(_gnd_net_),
            .in2(N__31859),
            .in3(N__32295),
            .lcout(n23_adj_1541),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i0_LC_12_14_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i0_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i0_LC_12_14_0 .LUT_INIT=16'b1010000000110011;
    LogicCell40 \SIG_DDS.dds_state_i0_LC_12_14_0  (
            .in0(N__35997),
            .in1(N__41284),
            .in2(N__31821),
            .in3(N__43044),
            .lcout(dds_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54314),
            .ce(N__36092),
            .sr(_gnd_net_));
    defparam i18462_3_lut_LC_12_14_1.C_ON=1'b0;
    defparam i18462_3_lut_LC_12_14_1.SEQ_MODE=4'b0000;
    defparam i18462_3_lut_LC_12_14_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18462_3_lut_LC_12_14_1 (
            .in0(N__31798),
            .in1(N__40976),
            .in2(_gnd_net_),
            .in3(N__57592),
            .lcout(n21072),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18477_3_lut_LC_12_14_3.C_ON=1'b0;
    defparam i18477_3_lut_LC_12_14_3.SEQ_MODE=4'b0000;
    defparam i18477_3_lut_LC_12_14_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 i18477_3_lut_LC_12_14_3 (
            .in0(N__31775),
            .in1(N__57593),
            .in2(_gnd_net_),
            .in3(N__32272),
            .lcout(n21087),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_12_14_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_12_14_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_12_14_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i1_2_lut_3_lut_LC_12_14_6 (
            .in0(N__43568),
            .in1(N__51879),
            .in2(_gnd_net_),
            .in3(N__55547),
            .lcout(n14_adj_1583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_256_LC_12_14_7.C_ON=1'b0;
    defparam i1_2_lut_adj_256_LC_12_14_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_256_LC_12_14_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_256_LC_12_14_7 (
            .in0(_gnd_net_),
            .in1(N__55545),
            .in2(_gnd_net_),
            .in3(N__50052),
            .lcout(n20856),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i0_LC_12_15_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i0_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i0_LC_12_15_0 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i0_LC_12_15_0  (
            .in0(N__36773),
            .in1(N__43047),
            .in2(N__42287),
            .in3(N__33967),
            .lcout(\SIG_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i1_LC_12_15_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i1_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i1_LC_12_15_1 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \SIG_DDS.tmp_buf_i1_LC_12_15_1  (
            .in0(N__32144),
            .in1(N__32112),
            .in2(N__42282),
            .in3(N__43052),
            .lcout(\SIG_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i2_LC_12_15_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i2_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i2_LC_12_15_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \SIG_DDS.tmp_buf_i2_LC_12_15_2  (
            .in0(N__32106),
            .in1(N__42248),
            .in2(N__47928),
            .in3(N__43049),
            .lcout(\SIG_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i3_LC_12_15_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i3_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i3_LC_12_15_3 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i3_LC_12_15_3  (
            .in0(N__43045),
            .in1(N__32100),
            .in2(N__42283),
            .in3(N__46923),
            .lcout(\SIG_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i15_LC_12_15_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i15_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i15_LC_12_15_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \SIG_DDS.tmp_buf_i15_LC_12_15_4  (
            .in0(N__32094),
            .in1(N__43048),
            .in2(N__32088),
            .in3(N__42262),
            .lcout(tmp_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i4_LC_12_15_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i4_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i4_LC_12_15_5 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \SIG_DDS.tmp_buf_i4_LC_12_15_5  (
            .in0(N__33806),
            .in1(N__43051),
            .in2(N__42284),
            .in3(N__32058),
            .lcout(\SIG_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i8_LC_12_15_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i8_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i8_LC_12_15_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \SIG_DDS.tmp_buf_i8_LC_12_15_6  (
            .in0(N__32301),
            .in1(N__42249),
            .in2(N__32043),
            .in3(N__43050),
            .lcout(\SIG_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i7_LC_12_15_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i7_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i7_LC_12_15_7 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i7_LC_12_15_7  (
            .in0(N__43046),
            .in1(N__32331),
            .in2(N__42285),
            .in3(N__32325),
            .lcout(\SIG_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54327),
            .ce(N__42089),
            .sr(_gnd_net_));
    defparam buf_dds0_i4_LC_12_16_0.C_ON=1'b0;
    defparam buf_dds0_i4_LC_12_16_0.SEQ_MODE=4'b1000;
    defparam buf_dds0_i4_LC_12_16_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i4_LC_12_16_0 (
            .in0(N__56446),
            .in1(N__33802),
            .in2(N__47805),
            .in3(N__47997),
            .lcout(buf_dds0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54339),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i12_LC_12_16_1.C_ON=1'b0;
    defparam acadc_skipCount_i12_LC_12_16_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i12_LC_12_16_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i12_LC_12_16_1 (
            .in0(N__56441),
            .in1(N__44323),
            .in2(N__41495),
            .in3(N__32294),
            .lcout(acadc_skipCount_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54339),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i6_LC_12_16_2.C_ON=1'b0;
    defparam buf_control_i6_LC_12_16_2.SEQ_MODE=4'b1000;
    defparam buf_control_i6_LC_12_16_2.LUT_INIT=16'b0111010000110000;
    LogicCell40 buf_control_i6_LC_12_16_2 (
            .in0(N__56445),
            .in1(N__41862),
            .in2(N__38675),
            .in3(N__45353),
            .lcout(buf_control_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54339),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i10_LC_12_16_3.C_ON=1'b0;
    defparam acadc_skipCount_i10_LC_12_16_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i10_LC_12_16_3.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i10_LC_12_16_3 (
            .in0(N__56440),
            .in1(N__44322),
            .in2(N__32273),
            .in3(N__44779),
            .lcout(acadc_skipCount_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54339),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i13_LC_12_16_4.C_ON=1'b0;
    defparam acadc_skipCount_i13_LC_12_16_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i13_LC_12_16_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i13_LC_12_16_4 (
            .in0(N__44321),
            .in1(N__43589),
            .in2(N__56540),
            .in3(N__32243),
            .lcout(acadc_skipCount_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54339),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i5_LC_12_16_5.C_ON=1'b0;
    defparam acadc_skipCount_i5_LC_12_16_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i5_LC_12_16_5.LUT_INIT=16'b0000110010101010;
    LogicCell40 acadc_skipCount_i5_LC_12_16_5 (
            .in0(N__52811),
            .in1(N__51438),
            .in2(N__56539),
            .in3(N__44324),
            .lcout(acadc_skipCount_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54339),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_12_16_6.C_ON=1'b0;
    defparam i4_4_lut_LC_12_16_6.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_12_16_6.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_LC_12_16_6 (
            .in0(N__32538),
            .in1(N__32400),
            .in2(N__50087),
            .in3(N__52810),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_232_LC_12_16_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_232_LC_12_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_232_LC_12_16_7.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_adj_232_LC_12_16_7 (
            .in0(N__32217),
            .in1(N__32178),
            .in2(_gnd_net_),
            .in3(N__34030),
            .lcout(n4_adj_1546),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_12_17_0.C_ON=1'b0;
    defparam i7_4_lut_LC_12_17_0.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_12_17_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i7_4_lut_LC_12_17_0 (
            .in0(N__32694),
            .in1(N__32457),
            .in2(N__41927),
            .in3(N__33820),
            .lcout(n23_adj_1501),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_12_17_2.C_ON=1'b0;
    defparam i8_4_lut_LC_12_17_2.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_12_17_2.LUT_INIT=16'b0111101111011110;
    LogicCell40 i8_4_lut_LC_12_17_2 (
            .in0(N__32496),
            .in1(N__32673),
            .in2(N__34074),
            .in3(N__32359),
            .lcout(n24_adj_1642),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i8_LC_12_17_3.C_ON=1'b0;
    defparam acadc_skipCount_i8_LC_12_17_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i8_LC_12_17_3.LUT_INIT=16'b0000101011001010;
    LogicCell40 acadc_skipCount_i8_LC_12_17_3 (
            .in0(N__43649),
            .in1(N__43824),
            .in2(N__44331),
            .in3(N__56471),
            .lcout(acadc_skipCount_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54353),
            .ce(),
            .sr(_gnd_net_));
    defparam i15345_2_lut_3_lut_LC_12_17_4.C_ON=1'b0;
    defparam i15345_2_lut_3_lut_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam i15345_2_lut_3_lut_LC_12_17_4.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15345_2_lut_3_lut_LC_12_17_4 (
            .in0(N__51878),
            .in1(N__37431),
            .in2(_gnd_net_),
            .in3(N__55546),
            .lcout(n14_adj_1556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i15_LC_12_17_5.C_ON=1'b0;
    defparam acadc_skipCount_i15_LC_12_17_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i15_LC_12_17_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i15_LC_12_17_5 (
            .in0(N__32360),
            .in1(N__56467),
            .in2(N__42816),
            .in3(N__44299),
            .lcout(acadc_skipCount_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54353),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i9_LC_12_17_6.C_ON=1'b0;
    defparam acadc_skipCount_i9_LC_12_17_6.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i9_LC_12_17_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i9_LC_12_17_6 (
            .in0(N__44297),
            .in1(N__40121),
            .in2(N__56548),
            .in3(N__34073),
            .lcout(acadc_skipCount_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54353),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i14_LC_12_17_7.C_ON=1'b0;
    defparam acadc_skipCount_i14_LC_12_17_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i14_LC_12_17_7.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i14_LC_12_17_7 (
            .in0(N__33821),
            .in1(N__56466),
            .in2(N__45358),
            .in3(N__44298),
            .lcout(acadc_skipCount_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54353),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i0_LC_12_18_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i0_LC_12_18_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i0_LC_12_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i0_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(N__37954),
            .in2(N__38451),
            .in3(_gnd_net_),
            .lcout(acadc_skipcnt_0),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(n19610),
            .clk(INVacadc_skipcnt_i0_i0C_net),
            .ce(N__32656),
            .sr(N__32346));
    defparam add_73_2_THRU_CRY_0_LC_12_18_1.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_0_LC_12_18_1.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_0_LC_12_18_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_0_LC_12_18_1 (
            .in0(_gnd_net_),
            .in1(N__58608),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19610),
            .carryout(n19610_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_1_LC_12_18_2.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_1_LC_12_18_2.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_1_LC_12_18_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_1_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__58621),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19610_THRU_CRY_0_THRU_CO),
            .carryout(n19610_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_2_LC_12_18_3.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_2_LC_12_18_3.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_2_LC_12_18_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_2_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(N__58612),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19610_THRU_CRY_1_THRU_CO),
            .carryout(n19610_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_3_LC_12_18_4.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_3_LC_12_18_4.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_3_LC_12_18_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_3_LC_12_18_4 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__58622),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19610_THRU_CRY_2_THRU_CO),
            .carryout(n19610_THRU_CRY_3_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_4_LC_12_18_5.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_4_LC_12_18_5.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_4_LC_12_18_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_4_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(N__58616),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19610_THRU_CRY_3_THRU_CO),
            .carryout(n19610_THRU_CRY_4_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_5_LC_12_18_6.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_5_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_5_LC_12_18_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_5_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__58623),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19610_THRU_CRY_4_THRU_CO),
            .carryout(n19610_THRU_CRY_5_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_6_LC_12_18_7.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_6_LC_12_18_7.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_6_LC_12_18_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_6_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(N__58620),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19610_THRU_CRY_5_THRU_CO),
            .carryout(n19610_THRU_CRY_6_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i1_LC_12_19_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i1_LC_12_19_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i1_LC_12_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i1_LC_12_19_0 (
            .in0(_gnd_net_),
            .in1(N__32418),
            .in2(_gnd_net_),
            .in3(N__32406),
            .lcout(acadc_skipcnt_1),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(n19611),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i2_LC_12_19_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i2_LC_12_19_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i2_LC_12_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i2_LC_12_19_1 (
            .in0(_gnd_net_),
            .in1(N__41579),
            .in2(_gnd_net_),
            .in3(N__32403),
            .lcout(acadc_skipcnt_2),
            .ltout(),
            .carryin(n19611),
            .carryout(n19612),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i3_LC_12_19_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i3_LC_12_19_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i3_LC_12_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i3_LC_12_19_2 (
            .in0(_gnd_net_),
            .in1(N__32399),
            .in2(_gnd_net_),
            .in3(N__32385),
            .lcout(acadc_skipcnt_3),
            .ltout(),
            .carryin(n19612),
            .carryout(n19613),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i4_LC_12_19_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i4_LC_12_19_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i4_LC_12_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i4_LC_12_19_3 (
            .in0(_gnd_net_),
            .in1(N__32555),
            .in2(_gnd_net_),
            .in3(N__32541),
            .lcout(acadc_skipcnt_4),
            .ltout(),
            .carryin(n19613),
            .carryout(n19614),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i5_LC_12_19_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i5_LC_12_19_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i5_LC_12_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i5_LC_12_19_4 (
            .in0(_gnd_net_),
            .in1(N__32537),
            .in2(_gnd_net_),
            .in3(N__32523),
            .lcout(acadc_skipcnt_5),
            .ltout(),
            .carryin(n19614),
            .carryout(n19615),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i6_LC_12_19_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i6_LC_12_19_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i6_LC_12_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i6_LC_12_19_5 (
            .in0(_gnd_net_),
            .in1(N__38426),
            .in2(_gnd_net_),
            .in3(N__32520),
            .lcout(acadc_skipcnt_6),
            .ltout(),
            .carryin(n19615),
            .carryout(n19616),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i7_LC_12_19_6.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i7_LC_12_19_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i7_LC_12_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i7_LC_12_19_6 (
            .in0(_gnd_net_),
            .in1(N__41597),
            .in2(_gnd_net_),
            .in3(N__32517),
            .lcout(acadc_skipcnt_7),
            .ltout(),
            .carryin(n19616),
            .carryout(n19617),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i8_LC_12_19_7.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i8_LC_12_19_7.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i8_LC_12_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i8_LC_12_19_7 (
            .in0(_gnd_net_),
            .in1(N__32513),
            .in2(_gnd_net_),
            .in3(N__32499),
            .lcout(acadc_skipcnt_8),
            .ltout(),
            .carryin(n19617),
            .carryout(n19618),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32658),
            .sr(N__32622));
    defparam acadc_skipcnt_i0_i9_LC_12_20_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i9_LC_12_20_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i9_LC_12_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i9_LC_12_20_0 (
            .in0(_gnd_net_),
            .in1(N__32495),
            .in2(_gnd_net_),
            .in3(N__32481),
            .lcout(acadc_skipcnt_9),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(n19619),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32657),
            .sr(N__32618));
    defparam acadc_skipcnt_i0_i10_LC_12_20_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i10_LC_12_20_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i10_LC_12_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i10_LC_12_20_1 (
            .in0(_gnd_net_),
            .in1(N__32474),
            .in2(_gnd_net_),
            .in3(N__32460),
            .lcout(acadc_skipcnt_10),
            .ltout(),
            .carryin(n19619),
            .carryout(n19620),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32657),
            .sr(N__32618));
    defparam acadc_skipcnt_i0_i11_LC_12_20_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i11_LC_12_20_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i11_LC_12_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i11_LC_12_20_2 (
            .in0(_gnd_net_),
            .in1(N__32456),
            .in2(_gnd_net_),
            .in3(N__32442),
            .lcout(acadc_skipcnt_11),
            .ltout(),
            .carryin(n19620),
            .carryout(n19621),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32657),
            .sr(N__32618));
    defparam acadc_skipcnt_i0_i12_LC_12_20_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i12_LC_12_20_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i12_LC_12_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i12_LC_12_20_3 (
            .in0(_gnd_net_),
            .in1(N__32435),
            .in2(_gnd_net_),
            .in3(N__32421),
            .lcout(acadc_skipcnt_12),
            .ltout(),
            .carryin(n19621),
            .carryout(n19622),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32657),
            .sr(N__32618));
    defparam acadc_skipcnt_i0_i13_LC_12_20_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i13_LC_12_20_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i13_LC_12_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i13_LC_12_20_4 (
            .in0(_gnd_net_),
            .in1(N__32711),
            .in2(_gnd_net_),
            .in3(N__32697),
            .lcout(acadc_skipcnt_13),
            .ltout(),
            .carryin(n19622),
            .carryout(n19623),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32657),
            .sr(N__32618));
    defparam acadc_skipcnt_i0_i14_LC_12_20_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i14_LC_12_20_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i14_LC_12_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i14_LC_12_20_5 (
            .in0(_gnd_net_),
            .in1(N__32693),
            .in2(_gnd_net_),
            .in3(N__32679),
            .lcout(acadc_skipcnt_14),
            .ltout(),
            .carryin(n19623),
            .carryout(n19624),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32657),
            .sr(N__32618));
    defparam acadc_skipcnt_i0_i15_LC_12_20_6.C_ON=1'b0;
    defparam acadc_skipcnt_i0_i15_LC_12_20_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i15_LC_12_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i15_LC_12_20_6 (
            .in0(_gnd_net_),
            .in1(N__32672),
            .in2(_gnd_net_),
            .in3(N__32676),
            .lcout(acadc_skipcnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32657),
            .sr(N__32618));
    defparam \ADC_VDC.i19363_4_lut_LC_13_3_0 .C_ON=1'b0;
    defparam \ADC_VDC.i19363_4_lut_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19363_4_lut_LC_13_3_0 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \ADC_VDC.i19363_4_lut_LC_13_3_0  (
            .in0(N__48481),
            .in1(N__32567),
            .in2(N__48835),
            .in3(N__34338),
            .lcout(\ADC_VDC.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i2_LC_13_3_2 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i2_LC_13_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i2_LC_13_3_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ADC_VDC.adc_state_i2_LC_13_3_2  (
            .in0(N__48758),
            .in1(N__48277),
            .in2(_gnd_net_),
            .in3(N__47359),
            .lcout(adc_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53261),
            .ce(N__32598),
            .sr(N__32589));
    defparam \ADC_VDC.i19412_4_lut_LC_13_3_3 .C_ON=1'b0;
    defparam \ADC_VDC.i19412_4_lut_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19412_4_lut_LC_13_3_3 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \ADC_VDC.i19412_4_lut_LC_13_3_3  (
            .in0(N__48480),
            .in1(N__32577),
            .in2(N__48773),
            .in3(N__47480),
            .lcout(\ADC_VDC.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i2_2_lut_LC_13_3_4 .C_ON=1'b0;
    defparam \ADC_VDC.i2_2_lut_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i2_2_lut_LC_13_3_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i2_2_lut_LC_13_3_4  (
            .in0(_gnd_net_),
            .in1(N__48275),
            .in2(_gnd_net_),
            .in3(N__47358),
            .lcout(\ADC_VDC.n7_adj_1398 ),
            .ltout(\ADC_VDC.n7_adj_1398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_11_LC_13_3_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_11_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_11_LC_13_3_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_11_LC_13_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32571),
            .in3(N__47481),
            .lcout(\ADC_VDC.n77 ),
            .ltout(\ADC_VDC.n77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_16_LC_13_3_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_16_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_16_LC_13_3_6 .LUT_INIT=16'b1011111110101110;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_16_LC_13_3_6  (
            .in0(N__48754),
            .in1(N__48479),
            .in2(N__32787),
            .in3(N__32784),
            .lcout(),
            .ltout(\ADC_VDC.n72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_17_LC_13_3_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_17_LC_13_3_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_17_LC_13_3_7 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_17_LC_13_3_7  (
            .in0(N__48276),
            .in1(N__32778),
            .in2(N__32772),
            .in3(N__34806),
            .lcout(\ADC_VDC.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i37_4_lut_LC_13_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.i37_4_lut_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i37_4_lut_LC_13_4_0 .LUT_INIT=16'b1101101001010010;
    LogicCell40 \ADC_VDC.i37_4_lut_LC_13_4_0  (
            .in0(N__47334),
            .in1(N__48288),
            .in2(N__47491),
            .in3(N__32904),
            .lcout(),
            .ltout(\ADC_VDC.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_13_LC_13_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_13_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_13_LC_13_4_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_13_LC_13_4_1  (
            .in0(N__48455),
            .in1(N__48774),
            .in2(N__32769),
            .in3(N__34323),
            .lcout(\ADC_VDC.n20811 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_13_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_13_4_2 .LUT_INIT=16'b0010110001101100;
    LogicCell40 \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_13_4_2  (
            .in0(N__47333),
            .in1(N__48287),
            .in2(N__48844),
            .in3(N__32726),
            .lcout(),
            .ltout(\ADC_VDC.n22195_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.n22195_bdd_4_lut_4_lut_LC_13_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.n22195_bdd_4_lut_4_lut_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.n22195_bdd_4_lut_4_lut_LC_13_4_3 .LUT_INIT=16'b1010010011110100;
    LogicCell40 \ADC_VDC.n22195_bdd_4_lut_4_lut_LC_13_4_3  (
            .in0(N__48709),
            .in1(N__34329),
            .in2(N__32766),
            .in3(N__47335),
            .lcout(),
            .ltout(\ADC_VDC.n22198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i1_LC_13_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i1_LC_13_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i1_LC_13_4_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.adc_state_i1_LC_13_4_4  (
            .in0(N__48778),
            .in1(N__48456),
            .in2(N__32763),
            .in3(N__32760),
            .lcout(\ADC_VDC.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53265),
            .ce(N__32745),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_14_LC_13_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_14_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_14_LC_13_4_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_14_LC_13_4_5  (
            .in0(_gnd_net_),
            .in1(N__36708),
            .in2(_gnd_net_),
            .in3(N__34845),
            .lcout(),
            .ltout(\ADC_VDC.n6_adj_1399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_adj_15_LC_13_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_adj_15_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_adj_15_LC_13_4_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \ADC_VDC.i4_4_lut_adj_15_LC_13_4_6  (
            .in0(N__36920),
            .in1(N__36611),
            .in2(N__32736),
            .in3(N__36645),
            .lcout(\ADC_VDC.n10536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18983_4_lut_LC_13_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i18983_4_lut_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18983_4_lut_LC_13_4_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ADC_VDC.i18983_4_lut_LC_13_4_7  (
            .in0(N__36612),
            .in1(N__36921),
            .in2(N__48529),
            .in3(N__34311),
            .lcout(\ADC_VDC.n21229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i0_LC_13_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i0_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i0_LC_13_5_4 .LUT_INIT=16'b0000000001110110;
    LogicCell40 \ADC_VDC.adc_state_i0_LC_13_5_4  (
            .in0(N__48784),
            .in1(N__48530),
            .in2(N__47489),
            .in3(N__47357),
            .lcout(\ADC_VDC.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53207),
            .ce(N__32898),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i7_12189_12190_reset_LC_13_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12189_12190_reset_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i7_12189_12190_reset_LC_13_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_12189_12190_reset_LC_13_6_0  (
            .in0(N__37344),
            .in1(N__44445),
            .in2(_gnd_net_),
            .in3(N__42387),
            .lcout(\comm_spi.n14608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52546),
            .ce(),
            .sr(N__35108));
    defparam comm_buf_2__i1_LC_13_7_0.C_ON=1'b0;
    defparam comm_buf_2__i1_LC_13_7_0.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i1_LC_13_7_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i1_LC_13_7_0 (
            .in0(N__45725),
            .in1(N__32802),
            .in2(_gnd_net_),
            .in3(N__51800),
            .lcout(comm_buf_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54274),
            .ce(N__33093),
            .sr(N__33071));
    defparam mux_130_Mux_1_i19_3_lut_LC_13_7_1.C_ON=1'b0;
    defparam mux_130_Mux_1_i19_3_lut_LC_13_7_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i19_3_lut_LC_13_7_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_130_Mux_1_i19_3_lut_LC_13_7_1 (
            .in0(N__57757),
            .in1(_gnd_net_),
            .in2(N__32871),
            .in3(N__33713),
            .lcout(),
            .ltout(n19_adj_1491_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i22_3_lut_LC_13_7_2.C_ON=1'b0;
    defparam mux_130_Mux_1_i22_3_lut_LC_13_7_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i22_3_lut_LC_13_7_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_1_i22_3_lut_LC_13_7_2 (
            .in0(_gnd_net_),
            .in1(N__32846),
            .in2(N__32823),
            .in3(N__53720),
            .lcout(),
            .ltout(n22_adj_1488_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i30_3_lut_LC_13_7_3.C_ON=1'b0;
    defparam mux_130_Mux_1_i30_3_lut_LC_13_7_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i30_3_lut_LC_13_7_3.LUT_INIT=16'b1101100011011000;
    LogicCell40 mux_130_Mux_1_i30_3_lut_LC_13_7_3 (
            .in0(N__54707),
            .in1(N__32820),
            .in2(N__32805),
            .in3(_gnd_net_),
            .lcout(n30_adj_1506),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19734_LC_13_7_4.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19734_LC_13_7_4.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19734_LC_13_7_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_0__bdd_4_lut_19734_LC_13_7_4 (
            .in0(N__32796),
            .in1(N__50658),
            .in2(N__45684),
            .in3(N__52331),
            .lcout(),
            .ltout(n22249_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22249_bdd_4_lut_LC_13_7_5.C_ON=1'b0;
    defparam n22249_bdd_4_lut_LC_13_7_5.SEQ_MODE=4'b0000;
    defparam n22249_bdd_4_lut_LC_13_7_5.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22249_bdd_4_lut_LC_13_7_5 (
            .in0(N__52332),
            .in1(N__40145),
            .in2(N__32790),
            .in3(N__37447),
            .lcout(n22252),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19739_LC_13_7_6.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19739_LC_13_7_6.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19739_LC_13_7_6.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_0__bdd_4_lut_19739_LC_13_7_6 (
            .in0(N__32967),
            .in1(N__50657),
            .in2(N__45504),
            .in3(N__52330),
            .lcout(n22381),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i0_LC_13_8_0.C_ON=1'b0;
    defparam comm_buf_2__i0_LC_13_8_0.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i0_LC_13_8_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_2__i0_LC_13_8_0 (
            .in0(N__32994),
            .in1(N__51868),
            .in2(_gnd_net_),
            .in3(N__53038),
            .lcout(comm_buf_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__33092),
            .sr(N__33072));
    defparam comm_buf_2__i7_LC_13_8_1.C_ON=1'b0;
    defparam comm_buf_2__i7_LC_13_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i7_LC_13_8_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i7_LC_13_8_1 (
            .in0(N__51867),
            .in1(N__50349),
            .in2(_gnd_net_),
            .in3(N__32982),
            .lcout(comm_buf_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__33092),
            .sr(N__33072));
    defparam comm_buf_2__i6_LC_13_8_2.C_ON=1'b0;
    defparam comm_buf_2__i6_LC_13_8_2.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i6_LC_13_8_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i6_LC_13_8_2 (
            .in0(N__46405),
            .in1(N__32961),
            .in2(_gnd_net_),
            .in3(N__51871),
            .lcout(comm_buf_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__33092),
            .sr(N__33072));
    defparam comm_buf_2__i5_LC_13_8_3.C_ON=1'b0;
    defparam comm_buf_2__i5_LC_13_8_3.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i5_LC_13_8_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i5_LC_13_8_3 (
            .in0(N__51866),
            .in1(N__52059),
            .in2(_gnd_net_),
            .in3(N__32946),
            .lcout(comm_buf_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__33092),
            .sr(N__33072));
    defparam comm_buf_2__i4_LC_13_8_4.C_ON=1'b0;
    defparam comm_buf_2__i4_LC_13_8_4.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i4_LC_13_8_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i4_LC_13_8_4 (
            .in0(N__46730),
            .in1(N__32934),
            .in2(_gnd_net_),
            .in3(N__51870),
            .lcout(comm_buf_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__33092),
            .sr(N__33072));
    defparam comm_buf_2__i3_LC_13_8_5.C_ON=1'b0;
    defparam comm_buf_2__i3_LC_13_8_5.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i3_LC_13_8_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i3_LC_13_8_5 (
            .in0(N__51865),
            .in1(N__51055),
            .in2(_gnd_net_),
            .in3(N__32925),
            .lcout(comm_buf_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__33092),
            .sr(N__33072));
    defparam comm_buf_2__i2_LC_13_8_6.C_ON=1'b0;
    defparam comm_buf_2__i2_LC_13_8_6.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i2_LC_13_8_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_2__i2_LC_13_8_6 (
            .in0(N__32916),
            .in1(N__47175),
            .in2(_gnd_net_),
            .in3(N__51869),
            .lcout(comm_buf_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54278),
            .ce(N__33092),
            .sr(N__33072));
    defparam mux_137_Mux_3_i4_3_lut_LC_13_9_0.C_ON=1'b0;
    defparam mux_137_Mux_3_i4_3_lut_LC_13_9_0.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_3_i4_3_lut_LC_13_9_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_137_Mux_3_i4_3_lut_LC_13_9_0 (
            .in0(N__39861),
            .in1(N__50669),
            .in2(_gnd_net_),
            .in3(N__42576),
            .lcout(),
            .ltout(n4_adj_1594_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18583_4_lut_LC_13_9_1.C_ON=1'b0;
    defparam i18583_4_lut_LC_13_9_1.SEQ_MODE=4'b0000;
    defparam i18583_4_lut_LC_13_9_1.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18583_4_lut_LC_13_9_1 (
            .in0(N__52344),
            .in1(N__33780),
            .in2(N__32907),
            .in3(N__50688),
            .lcout(n21193),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19744_LC_13_9_2.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19744_LC_13_9_2.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19744_LC_13_9_2.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_0__bdd_4_lut_19744_LC_13_9_2 (
            .in0(N__33024),
            .in1(N__50668),
            .in2(N__45435),
            .in3(N__52345),
            .lcout(),
            .ltout(n22387_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22387_bdd_4_lut_LC_13_9_3.C_ON=1'b0;
    defparam n22387_bdd_4_lut_LC_13_9_3.SEQ_MODE=4'b0000;
    defparam n22387_bdd_4_lut_LC_13_9_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22387_bdd_4_lut_LC_13_9_3 (
            .in0(N__52346),
            .in1(N__44222),
            .in2(N__33018),
            .in3(N__51012),
            .lcout(),
            .ltout(n22390_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i3_LC_13_9_4.C_ON=1'b0;
    defparam comm_tx_buf_i3_LC_13_9_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i3_LC_13_9_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_tx_buf_i3_LC_13_9_4 (
            .in0(_gnd_net_),
            .in1(N__33015),
            .in2(N__33009),
            .in3(N__50538),
            .lcout(comm_tx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__45234),
            .sr(N__45172));
    defparam mux_137_Mux_7_i4_3_lut_LC_13_9_5.C_ON=1'b0;
    defparam mux_137_Mux_7_i4_3_lut_LC_13_9_5.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_7_i4_3_lut_LC_13_9_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_137_Mux_7_i4_3_lut_LC_13_9_5 (
            .in0(N__50670),
            .in1(N__39942),
            .in2(_gnd_net_),
            .in3(N__42675),
            .lcout(),
            .ltout(n4_adj_1587_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18565_4_lut_LC_13_9_6.C_ON=1'b0;
    defparam i18565_4_lut_LC_13_9_6.SEQ_MODE=4'b0000;
    defparam i18565_4_lut_LC_13_9_6.LUT_INIT=16'b0010001011110000;
    LogicCell40 i18565_4_lut_LC_13_9_6 (
            .in0(N__33047),
            .in1(N__50671),
            .in2(N__33006),
            .in3(N__52347),
            .lcout(),
            .ltout(n21175_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i7_LC_13_9_7.C_ON=1'b0;
    defparam comm_tx_buf_i7_LC_13_9_7.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i7_LC_13_9_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_tx_buf_i7_LC_13_9_7 (
            .in0(N__50539),
            .in1(_gnd_net_),
            .in2(N__33003),
            .in3(N__34221),
            .lcout(comm_tx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54281),
            .ce(N__45234),
            .sr(N__45172));
    defparam i458_2_lut_LC_13_10_0.C_ON=1'b0;
    defparam i458_2_lut_LC_13_10_0.SEQ_MODE=4'b0000;
    defparam i458_2_lut_LC_13_10_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 i458_2_lut_LC_13_10_0 (
            .in0(N__50038),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49846),
            .lcout(n2358),
            .ltout(n2358_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_255_LC_13_10_1.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_255_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_255_LC_13_10_1.LUT_INIT=16'b0000000001000000;
    LogicCell40 i1_2_lut_4_lut_adj_255_LC_13_10_1 (
            .in0(N__50753),
            .in1(N__52370),
            .in2(N__33000),
            .in3(N__52266),
            .lcout(n20850),
            .ltout(n20850_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i36_4_lut_LC_13_10_2.C_ON=1'b0;
    defparam i36_4_lut_LC_13_10_2.SEQ_MODE=4'b0000;
    defparam i36_4_lut_LC_13_10_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 i36_4_lut_LC_13_10_2 (
            .in0(N__51799),
            .in1(N__45636),
            .in2(N__32997),
            .in3(N__33894),
            .lcout(),
            .ltout(n31_adj_1613_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_270_LC_13_10_3.C_ON=1'b0;
    defparam i1_3_lut_adj_270_LC_13_10_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_270_LC_13_10_3.LUT_INIT=16'b1100110011000000;
    LogicCell40 i1_3_lut_adj_270_LC_13_10_3 (
            .in0(_gnd_net_),
            .in1(N__45927),
            .in2(N__33096),
            .in3(N__45881),
            .lcout(n12085),
            .ltout(n12085_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12351_2_lut_LC_13_10_4.C_ON=1'b0;
    defparam i12351_2_lut_LC_13_10_4.SEQ_MODE=4'b0000;
    defparam i12351_2_lut_LC_13_10_4.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12351_2_lut_LC_13_10_4 (
            .in0(N__56863),
            .in1(_gnd_net_),
            .in2(N__33075),
            .in3(_gnd_net_),
            .lcout(n14764),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_214_LC_13_10_5.C_ON=1'b0;
    defparam i1_3_lut_adj_214_LC_13_10_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_214_LC_13_10_5.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_3_lut_adj_214_LC_13_10_5 (
            .in0(N__49586),
            .in1(N__33030),
            .in2(_gnd_net_),
            .in3(N__56864),
            .lcout(n12228),
            .ltout(n12228_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i7_LC_13_10_6.C_ON=1'b0;
    defparam comm_buf_6__i7_LC_13_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i7_LC_13_10_6.LUT_INIT=16'b0100111101000000;
    LogicCell40 comm_buf_6__i7_LC_13_10_6 (
            .in0(N__56865),
            .in1(N__50380),
            .in2(N__33051),
            .in3(N__33048),
            .lcout(comm_buf_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i6_LC_13_10_7.C_ON=1'b0;
    defparam comm_buf_6__i6_LC_13_10_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i6_LC_13_10_7.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i6_LC_13_10_7 (
            .in0(N__45593),
            .in1(N__56866),
            .in2(N__46448),
            .in3(N__34993),
            .lcout(comm_buf_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54289),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_213_LC_13_11_0.C_ON=1'b0;
    defparam i3_4_lut_adj_213_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_213_LC_13_11_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i3_4_lut_adj_213_LC_13_11_0 (
            .in0(N__51792),
            .in1(N__33036),
            .in2(N__37671),
            .in3(N__55518),
            .lcout(n20852),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i4_LC_13_11_1.C_ON=1'b0;
    defparam comm_cmd_i4_LC_13_11_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i4_LC_13_11_1.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i4_LC_13_11_1 (
            .in0(N__46000),
            .in1(N__46071),
            .in2(N__46755),
            .in3(N__49776),
            .lcout(comm_cmd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54294),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i0_LC_13_11_2.C_ON=1'b0;
    defparam comm_cmd_i0_LC_13_11_2.SEQ_MODE=4'b1000;
    defparam comm_cmd_i0_LC_13_11_2.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i0_LC_13_11_2 (
            .in0(N__57388),
            .in1(N__53040),
            .in2(N__46082),
            .in3(N__45999),
            .lcout(comm_cmd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54294),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_13_11_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_13_11_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_104_2_lut_LC_13_11_3  (
            .in0(N__55865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34897),
            .lcout(\comm_spi.data_tx_7__N_786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i5_LC_13_11_4.C_ON=1'b0;
    defparam comm_buf_6__i5_LC_13_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i5_LC_13_11_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_buf_6__i5_LC_13_11_4 (
            .in0(N__34996),
            .in1(N__52092),
            .in2(N__57088),
            .in3(N__42446),
            .lcout(comm_buf_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54294),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i0_LC_13_11_5.C_ON=1'b0;
    defparam comm_buf_6__i0_LC_13_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i0_LC_13_11_5.LUT_INIT=16'b0010001011110000;
    LogicCell40 comm_buf_6__i0_LC_13_11_5 (
            .in0(N__53039),
            .in1(N__56992),
            .in2(N__42317),
            .in3(N__34994),
            .lcout(comm_buf_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54294),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i3_LC_13_11_6.C_ON=1'b0;
    defparam comm_buf_6__i3_LC_13_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i3_LC_13_11_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_buf_6__i3_LC_13_11_6 (
            .in0(N__34995),
            .in1(N__51071),
            .in2(N__57087),
            .in3(N__33776),
            .lcout(comm_buf_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54294),
            .ce(),
            .sr(_gnd_net_));
    defparam i38_3_lut_LC_13_11_7.C_ON=1'b0;
    defparam i38_3_lut_LC_13_11_7.SEQ_MODE=4'b0000;
    defparam i38_3_lut_LC_13_11_7.LUT_INIT=16'b0101010110001000;
    LogicCell40 i38_3_lut_LC_13_11_7 (
            .in0(N__54868),
            .in1(N__57387),
            .in2(_gnd_net_),
            .in3(N__53489),
            .lcout(n22_adj_1615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i1_LC_13_12_0.C_ON=1'b0;
    defparam buf_dds1_i1_LC_13_12_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i1_LC_13_12_0.LUT_INIT=16'b1101000010000000;
    LogicCell40 buf_dds1_i1_LC_13_12_0 (
            .in0(N__44934),
            .in1(N__37440),
            .in2(N__40656),
            .in3(N__33758),
            .lcout(buf_dds1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54306),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i1_LC_13_12_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i1_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i1_LC_13_12_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i1_LC_13_12_1  (
            .in0(N__33458),
            .in1(N__33678),
            .in2(N__33709),
            .in3(N__33738),
            .lcout(buf_adcdata_vac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54306),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i10_LC_13_12_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i10_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i10_LC_13_12_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i10_LC_13_12_2  (
            .in0(N__33677),
            .in1(N__33459),
            .in2(N__35954),
            .in3(N__33128),
            .lcout(buf_adcdata_vac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54306),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i1_LC_13_12_3.C_ON=1'b0;
    defparam comm_cmd_i1_LC_13_12_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i1_LC_13_12_3.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i1_LC_13_12_3 (
            .in0(N__46001),
            .in1(N__46070),
            .in2(N__45794),
            .in3(N__54837),
            .lcout(comm_cmd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54306),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_13_12_4.C_ON=1'b0;
    defparam comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_13_12_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_13_12_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_13_12_4 (
            .in0(N__54836),
            .in1(N__57262),
            .in2(_gnd_net_),
            .in3(N__53458),
            .lcout(n9_adj_1416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i0_LC_13_12_5.C_ON=1'b0;
    defparam buf_dds1_i0_LC_13_12_5.SEQ_MODE=4'b1000;
    defparam buf_dds1_i0_LC_13_12_5.LUT_INIT=16'b1100000010001000;
    LogicCell40 buf_dds1_i0_LC_13_12_5 (
            .in0(N__33923),
            .in1(N__40631),
            .in2(N__43299),
            .in3(N__44935),
            .lcout(buf_dds1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54306),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_13_12_6.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_13_12_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_13_12_6.LUT_INIT=16'b1101110111111111;
    LogicCell40 i2_2_lut_3_lut_LC_13_12_6 (
            .in0(N__54835),
            .in1(N__57261),
            .in2(_gnd_net_),
            .in3(N__53457),
            .lcout(n10717),
            .ltout(n10717_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19112_4_lut_LC_13_12_7.C_ON=1'b0;
    defparam i19112_4_lut_LC_13_12_7.SEQ_MODE=4'b0000;
    defparam i19112_4_lut_LC_13_12_7.LUT_INIT=16'b0000101010001000;
    LogicCell40 i19112_4_lut_LC_13_12_7 (
            .in0(N__49271),
            .in1(N__33903),
            .in2(N__33897),
            .in3(N__54569),
            .lcout(n21344),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i5_LC_13_13_0.C_ON=1'b0;
    defparam buf_dds1_i5_LC_13_13_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i5_LC_13_13_0.LUT_INIT=16'b1110010011101110;
    LogicCell40 buf_dds1_i5_LC_13_13_0 (
            .in0(N__44931),
            .in1(N__33883),
            .in2(N__37496),
            .in3(N__57049),
            .lcout(buf_dds1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i3_LC_13_13_1.C_ON=1'b0;
    defparam comm_cmd_i3_LC_13_13_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i3_LC_13_13_1.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i3_LC_13_13_1 (
            .in0(N__46012),
            .in1(N__46079),
            .in2(N__51106),
            .in3(N__54601),
            .lcout(comm_cmd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i7_LC_13_13_2.C_ON=1'b0;
    defparam buf_dds1_i7_LC_13_13_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i7_LC_13_13_2.LUT_INIT=16'b1110010000000000;
    LogicCell40 buf_dds1_i7_LC_13_13_2 (
            .in0(N__44932),
            .in1(N__33847),
            .in2(N__50321),
            .in3(N__40637),
            .lcout(buf_dds1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_6_i23_3_lut_LC_13_13_3.C_ON=1'b0;
    defparam mux_128_Mux_6_i23_3_lut_LC_13_13_3.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_6_i23_3_lut_LC_13_13_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_128_Mux_6_i23_3_lut_LC_13_13_3 (
            .in0(N__57589),
            .in1(N__38674),
            .in2(_gnd_net_),
            .in3(N__33828),
            .lcout(n23_adj_1538),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i16_3_lut_LC_13_13_4.C_ON=1'b0;
    defparam mux_129_Mux_4_i16_3_lut_LC_13_13_4.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i16_3_lut_LC_13_13_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_4_i16_3_lut_LC_13_13_4 (
            .in0(N__33988),
            .in1(N__33807),
            .in2(_gnd_net_),
            .in3(N__57588),
            .lcout(n16_adj_1510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i8_LC_13_13_5.C_ON=1'b0;
    defparam req_data_cnt_i8_LC_13_13_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i8_LC_13_13_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i8_LC_13_13_5 (
            .in0(N__41741),
            .in1(N__37851),
            .in2(_gnd_net_),
            .in3(N__43876),
            .lcout(req_data_cnt_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i6_LC_13_13_6.C_ON=1'b0;
    defparam req_data_cnt_i6_LC_13_13_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i6_LC_13_13_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i6_LC_13_13_6 (
            .in0(N__47832),
            .in1(N__41740),
            .in2(_gnd_net_),
            .in3(N__40781),
            .lcout(req_data_cnt_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i4_LC_13_13_7.C_ON=1'b0;
    defparam buf_dds1_i4_LC_13_13_7.SEQ_MODE=4'b1000;
    defparam buf_dds1_i4_LC_13_13_7.LUT_INIT=16'b1100000010001000;
    LogicCell40 buf_dds1_i4_LC_13_13_7 (
            .in0(N__33992),
            .in1(N__40635),
            .in2(N__47784),
            .in3(N__44933),
            .lcout(buf_dds1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54319),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_284_LC_13_14_0.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_284_LC_13_14_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_284_LC_13_14_0.LUT_INIT=16'b0000000000000010;
    LogicCell40 i1_2_lut_4_lut_adj_284_LC_13_14_0 (
            .in0(N__49786),
            .in1(N__49732),
            .in2(N__49496),
            .in3(N__49696),
            .lcout(n20804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i6_LC_13_14_1.C_ON=1'b0;
    defparam comm_cmd_i6_LC_13_14_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i6_LC_13_14_1.LUT_INIT=16'b1110001000100010;
    LogicCell40 comm_cmd_i6_LC_13_14_1 (
            .in0(N__49733),
            .in1(N__46013),
            .in2(N__46464),
            .in3(N__46080),
            .lcout(comm_cmd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54332),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i3_LC_13_14_2.C_ON=1'b0;
    defparam acadc_skipCount_i3_LC_13_14_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i3_LC_13_14_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i3_LC_13_14_2 (
            .in0(N__56474),
            .in1(N__44325),
            .in2(N__51020),
            .in3(N__50080),
            .lcout(acadc_skipCount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54332),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i0_LC_13_14_3.C_ON=1'b0;
    defparam buf_dds0_i0_LC_13_14_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i0_LC_13_14_3.LUT_INIT=16'b0010001011110000;
    LogicCell40 buf_dds0_i0_LC_13_14_3 (
            .in0(N__43290),
            .in1(N__56475),
            .in2(N__33972),
            .in3(N__48012),
            .lcout(buf_dds0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54332),
            .ce(),
            .sr(_gnd_net_));
    defparam i15337_2_lut_3_lut_LC_13_14_6.C_ON=1'b0;
    defparam i15337_2_lut_3_lut_LC_13_14_6.SEQ_MODE=4'b0000;
    defparam i15337_2_lut_3_lut_LC_13_14_6.LUT_INIT=16'b0000000001010000;
    LogicCell40 i15337_2_lut_3_lut_LC_13_14_6 (
            .in0(N__55548),
            .in1(_gnd_net_),
            .in2(N__41491),
            .in3(N__51880),
            .lcout(n14_adj_1577),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_184_LC_13_14_7.C_ON=1'b0;
    defparam i3_4_lut_adj_184_LC_13_14_7.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_184_LC_13_14_7.LUT_INIT=16'b0111110110111110;
    LogicCell40 i3_4_lut_adj_184_LC_13_14_7 (
            .in0(N__38127),
            .in1(N__41049),
            .in2(N__43877),
            .in3(N__33940),
            .lcout(n19_adj_1607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i2_LC_13_15_0.C_ON=1'b0;
    defparam req_data_cnt_i2_LC_13_15_0.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i2_LC_13_15_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i2_LC_13_15_0 (
            .in0(N__37547),
            .in1(N__41729),
            .in2(_gnd_net_),
            .in3(N__46607),
            .lcout(req_data_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54346),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_312_LC_13_15_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_312_LC_13_15_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_312_LC_13_15_1.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_312_LC_13_15_1 (
            .in0(N__49695),
            .in1(N__49777),
            .in2(_gnd_net_),
            .in3(N__49731),
            .lcout(n20893),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i9_LC_13_15_2.C_ON=1'b0;
    defparam req_data_cnt_i9_LC_13_15_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i9_LC_13_15_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i9_LC_13_15_2 (
            .in0(N__37827),
            .in1(N__41730),
            .in2(_gnd_net_),
            .in3(N__34265),
            .lcout(req_data_cnt_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54346),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_264_LC_13_15_3.C_ON=1'b0;
    defparam i1_2_lut_adj_264_LC_13_15_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_264_LC_13_15_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_264_LC_13_15_3 (
            .in0(_gnd_net_),
            .in1(N__34112),
            .in2(_gnd_net_),
            .in3(N__41764),
            .lcout(n10697),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_13_15_4.C_ON=1'b0;
    defparam i13_4_lut_LC_13_15_4.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_13_15_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_LC_13_15_4 (
            .in0(N__34053),
            .in1(N__36066),
            .in2(N__36009),
            .in3(N__34122),
            .lcout(),
            .ltout(n29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_198_LC_13_15_5.C_ON=1'b0;
    defparam i1_3_lut_adj_198_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_198_LC_13_15_5.LUT_INIT=16'b1100110011001111;
    LogicCell40 i1_3_lut_adj_198_LC_13_15_5 (
            .in0(_gnd_net_),
            .in1(N__34284),
            .in2(N__34044),
            .in3(N__34005),
            .lcout(n16_adj_1603),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_stop_328_LC_13_15_6.C_ON=1'b0;
    defparam eis_stop_328_LC_13_15_6.SEQ_MODE=4'b1000;
    defparam eis_stop_328_LC_13_15_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 eis_stop_328_LC_13_15_6 (
            .in0(N__34285),
            .in1(N__40135),
            .in2(_gnd_net_),
            .in3(N__36247),
            .lcout(eis_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54346),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_173_LC_13_16_2.C_ON=1'b0;
    defparam i8_4_lut_adj_173_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_173_LC_13_16_2.LUT_INIT=16'b0111101111011110;
    LogicCell40 i8_4_lut_adj_173_LC_13_16_2 (
            .in0(N__38088),
            .in1(N__41175),
            .in2(N__36230),
            .in3(N__34261),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_178_LC_13_16_3.C_ON=1'b0;
    defparam i5_4_lut_adj_178_LC_13_16_3.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_178_LC_13_16_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_adj_178_LC_13_16_3 (
            .in0(N__38148),
            .in1(N__41229),
            .in2(N__40820),
            .in3(N__34087),
            .lcout(),
            .ltout(n21_adj_1492_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_187_LC_13_16_4.C_ON=1'b0;
    defparam i14_4_lut_adj_187_LC_13_16_4.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_187_LC_13_16_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_187_LC_13_16_4 (
            .in0(N__36039),
            .in1(N__34014),
            .in2(N__34008),
            .in3(N__36072),
            .lcout(n30_adj_1618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19084_2_lut_LC_13_16_5.C_ON=1'b0;
    defparam i19084_2_lut_LC_13_16_5.SEQ_MODE=4'b0000;
    defparam i19084_2_lut_LC_13_16_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19084_2_lut_LC_13_16_5 (
            .in0(_gnd_net_),
            .in1(N__57554),
            .in2(_gnd_net_),
            .in3(N__34088),
            .lcout(n21309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_306_LC_13_16_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_306_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_306_LC_13_16_6.LUT_INIT=16'b1111110111111101;
    LogicCell40 i1_2_lut_3_lut_adj_306_LC_13_16_6 (
            .in0(N__54602),
            .in1(N__37644),
            .in2(N__49495),
            .in3(_gnd_net_),
            .lcout(n20907),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_179_LC_13_16_7.C_ON=1'b0;
    defparam i4_4_lut_adj_179_LC_13_16_7.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_179_LC_13_16_7.LUT_INIT=16'b0111101111011110;
    LogicCell40 i4_4_lut_adj_179_LC_13_16_7 (
            .in0(N__50862),
            .in1(N__51155),
            .in2(N__50113),
            .in3(N__52840),
            .lcout(n20_adj_1617),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_13_17_0.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_13_17_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_13_17_0.LUT_INIT=16'b1111111111111011;
    LogicCell40 i2_3_lut_4_lut_LC_13_17_0 (
            .in0(N__41762),
            .in1(N__55542),
            .in2(N__51958),
            .in3(N__34111),
            .lcout(n10598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i12_LC_13_17_1.C_ON=1'b0;
    defparam req_data_cnt_i12_LC_13_17_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i12_LC_13_17_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i12_LC_13_17_1 (
            .in0(N__41699),
            .in1(N__37769),
            .in2(_gnd_net_),
            .in3(N__34089),
            .lcout(req_data_cnt_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54372),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i1_LC_13_17_2.C_ON=1'b0;
    defparam req_data_cnt_i1_LC_13_17_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i1_LC_13_17_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i1_LC_13_17_2 (
            .in0(N__37589),
            .in1(N__41700),
            .in2(_gnd_net_),
            .in3(N__37085),
            .lcout(req_data_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54372),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i3_LC_13_17_3.C_ON=1'b0;
    defparam req_data_cnt_i3_LC_13_17_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i3_LC_13_17_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 req_data_cnt_i3_LC_13_17_3 (
            .in0(N__41701),
            .in1(_gnd_net_),
            .in2(N__50117),
            .in3(N__47096),
            .lcout(req_data_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54372),
            .ce(),
            .sr(_gnd_net_));
    defparam n22375_bdd_4_lut_LC_13_17_4.C_ON=1'b0;
    defparam n22375_bdd_4_lut_LC_13_17_4.SEQ_MODE=4'b0000;
    defparam n22375_bdd_4_lut_LC_13_17_4.LUT_INIT=16'b1011101010011000;
    LogicCell40 n22375_bdd_4_lut_LC_13_17_4 (
            .in0(N__34245),
            .in1(N__55022),
            .in2(N__36366),
            .in3(N__34072),
            .lcout(n22378),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_263_LC_13_17_5.C_ON=1'b0;
    defparam i1_4_lut_adj_263_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_263_LC_13_17_5.LUT_INIT=16'b1000100010001100;
    LogicCell40 i1_4_lut_adj_263_LC_13_17_5 (
            .in0(N__56400),
            .in1(N__57126),
            .in2(N__44409),
            .in3(N__41763),
            .lcout(n12399),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15347_2_lut_3_lut_LC_13_17_6.C_ON=1'b0;
    defparam i15347_2_lut_3_lut_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam i15347_2_lut_3_lut_LC_13_17_6.LUT_INIT=16'b0001000100000000;
    LogicCell40 i15347_2_lut_3_lut_LC_13_17_6 (
            .in0(N__51876),
            .in1(N__55543),
            .in2(_gnd_net_),
            .in3(N__43815),
            .lcout(n14_adj_1550),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15339_2_lut_3_lut_LC_13_17_7.C_ON=1'b0;
    defparam i15339_2_lut_3_lut_LC_13_17_7.SEQ_MODE=4'b0000;
    defparam i15339_2_lut_3_lut_LC_13_17_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15339_2_lut_3_lut_LC_13_17_7 (
            .in0(N__55544),
            .in1(N__44749),
            .in2(_gnd_net_),
            .in3(N__51877),
            .lcout(n14_adj_1579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6449_3_lut_LC_13_18_1.C_ON=1'b0;
    defparam i6449_3_lut_LC_13_18_1.SEQ_MODE=4'b0000;
    defparam i6449_3_lut_LC_13_18_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6449_3_lut_LC_13_18_1 (
            .in0(N__37424),
            .in1(N__36288),
            .in2(_gnd_net_),
            .in3(N__47683),
            .lcout(n8_adj_1573),
            .ltout(n8_adj_1573_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i1_LC_13_18_2.C_ON=1'b0;
    defparam data_index_i1_LC_13_18_2.SEQ_MODE=4'b1000;
    defparam data_index_i1_LC_13_18_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 data_index_i1_LC_13_18_2 (
            .in0(N__57133),
            .in1(N__56512),
            .in2(N__34299),
            .in3(N__36477),
            .lcout(data_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54386),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19754_LC_13_18_3.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19754_LC_13_18_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19754_LC_13_18_3.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19754_LC_13_18_3 (
            .in0(N__57553),
            .in1(N__34295),
            .in2(N__55146),
            .in3(N__34266),
            .lcout(n22375),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22381_bdd_4_lut_LC_13_18_6.C_ON=1'b0;
    defparam n22381_bdd_4_lut_LC_13_18_6.SEQ_MODE=4'b0000;
    defparam n22381_bdd_4_lut_LC_13_18_6.LUT_INIT=16'b1110001111100000;
    LogicCell40 n22381_bdd_4_lut_LC_13_18_6 (
            .in0(N__50318),
            .in1(N__52413),
            .in2(N__34239),
            .in3(N__42802),
            .lcout(n22384),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds0_304_LC_13_18_7.C_ON=1'b0;
    defparam trig_dds0_304_LC_13_18_7.SEQ_MODE=4'b1000;
    defparam trig_dds0_304_LC_13_18_7.LUT_INIT=16'b0010111000100010;
    LogicCell40 trig_dds0_304_LC_13_18_7 (
            .in0(N__42124),
            .in1(N__34206),
            .in2(N__56556),
            .in3(N__57134),
            .lcout(trig_dds0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54386),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.SCLK_27_LC_13_19_2 .C_ON=1'b0;
    defparam \SIG_DDS.SCLK_27_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.SCLK_27_LC_13_19_2 .LUT_INIT=16'b0100000011101101;
    LogicCell40 \SIG_DDS.SCLK_27_LC_13_19_2  (
            .in0(N__42958),
            .in1(N__34178),
            .in2(N__41336),
            .in3(N__42189),
            .lcout(DDS_SCK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54399),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i23_4_lut_LC_13_19_3 .C_ON=1'b0;
    defparam \SIG_DDS.i23_4_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i23_4_lut_LC_13_19_3 .LUT_INIT=16'b1010101110011001;
    LogicCell40 \SIG_DDS.i23_4_lut_LC_13_19_3  (
            .in0(N__42188),
            .in1(N__42956),
            .in2(N__42120),
            .in3(N__41327),
            .lcout(\SIG_DDS.n9_adj_1393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i2_LC_13_19_4 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i2_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i2_LC_13_19_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \SIG_DDS.dds_state_i2_LC_13_19_4  (
            .in0(N__42957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42190),
            .lcout(dds_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54399),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i1_LC_13_20_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i1_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i1_LC_13_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \SIG_DDS.dds_state_i1_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__41337),
            .in2(_gnd_net_),
            .in3(N__42197),
            .lcout(dds_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54413),
            .ce(N__36096),
            .sr(N__43060));
    defparam \comm_spi.i12188_3_lut_LC_14_3_0 .C_ON=1'b0;
    defparam \comm_spi.i12188_3_lut_LC_14_3_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12188_3_lut_LC_14_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i12188_3_lut_LC_14_3_0  (
            .in0(N__34167),
            .in1(N__34155),
            .in2(_gnd_net_),
            .in3(N__35165),
            .lcout(ICE_SPI_MISO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_14_3_4 .C_ON=1'b0;
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_14_3_4 .LUT_INIT=16'b1100101101000011;
    LogicCell40 \ADC_VDC.i40_3_lut_4_lut_LC_14_3_4  (
            .in0(N__48298),
            .in1(N__47377),
            .in2(N__47492),
            .in3(N__34826),
            .lcout(\ADC_VDC.n19_adj_1401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19327_4_lut_LC_14_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.i19327_4_lut_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19327_4_lut_LC_14_4_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \ADC_VDC.i19327_4_lut_LC_14_4_1  (
            .in0(N__36639),
            .in1(N__36604),
            .in2(N__36707),
            .in3(N__36668),
            .lcout(),
            .ltout(\ADC_VDC.n21323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19100_4_lut_LC_14_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.i19100_4_lut_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19100_4_lut_LC_14_4_2 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \ADC_VDC.i19100_4_lut_LC_14_4_2  (
            .in0(N__36912),
            .in1(N__34305),
            .in2(N__34332),
            .in3(N__47332),
            .lcout(\ADC_VDC.n21320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18357_2_lut_LC_14_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i18357_2_lut_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18357_2_lut_LC_14_4_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ADC_VDC.i18357_2_lut_LC_14_4_3  (
            .in0(N__47482),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48300),
            .lcout(\ADC_VDC.n20965 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_2_lut_LC_14_4_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_2_lut_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_2_lut_LC_14_4_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_2_lut_LC_14_4_4  (
            .in0(N__42495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55810),
            .lcout(\comm_spi.data_tx_7__N_795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_adj_12_LC_14_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_adj_12_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_adj_12_LC_14_4_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ADC_VDC.i4_4_lut_adj_12_LC_14_4_5  (
            .in0(N__36638),
            .in1(N__36879),
            .in2(N__36706),
            .in3(N__36667),
            .lcout(),
            .ltout(\ADC_VDC.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i5_3_lut_LC_14_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.i5_3_lut_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i5_3_lut_LC_14_4_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \ADC_VDC.i5_3_lut_LC_14_4_6  (
            .in0(_gnd_net_),
            .in1(N__36826),
            .in2(N__34314),
            .in3(N__36853),
            .lcout(\ADC_VDC.n20812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i2_3_lut_LC_14_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i2_3_lut_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i2_3_lut_LC_14_4_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ADC_VDC.i2_3_lut_LC_14_4_7  (
            .in0(N__36854),
            .in1(N__36880),
            .in2(_gnd_net_),
            .in3(N__36827),
            .lcout(\ADC_VDC.n20784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_LC_14_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_LC_14_5_0 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \ADC_VDC.i1_4_lut_LC_14_5_0  (
            .in0(N__47348),
            .in1(N__48536),
            .in2(N__34854),
            .in3(N__48219),
            .lcout(\ADC_VDC.n18550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_9_LC_14_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_9_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_9_LC_14_5_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_9_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__36603),
            .in2(_gnd_net_),
            .in3(N__36640),
            .lcout(\ADC_VDC.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i15111_2_lut_LC_14_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.i15111_2_lut_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i15111_2_lut_LC_14_5_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i15111_2_lut_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__48792),
            .in2(_gnd_net_),
            .in3(N__48297),
            .lcout(\ADC_VDC.n17509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_4_lut_LC_14_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_4_lut_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_4_lut_LC_14_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i1_2_lut_4_lut_LC_14_5_3  (
            .in0(N__36825),
            .in1(N__36852),
            .in2(N__36882),
            .in3(N__36666),
            .lcout(\ADC_VDC.n11265 ),
            .ltout(\ADC_VDC.n11265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_LC_14_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_LC_14_5_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \ADC_VDC.i4_4_lut_LC_14_5_4  (
            .in0(N__36919),
            .in1(N__34839),
            .in2(N__34833),
            .in3(N__36704),
            .lcout(\ADC_VDC.n15 ),
            .ltout(\ADC_VDC.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18386_2_lut_LC_14_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i18386_2_lut_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18386_2_lut_LC_14_5_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ADC_VDC.i18386_2_lut_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34809),
            .in3(N__47347),
            .lcout(\ADC_VDC.n20996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i19328_4_lut_LC_14_5_7 .C_ON=1'b0;
    defparam \CLK_DDS.i19328_4_lut_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19328_4_lut_LC_14_5_7 .LUT_INIT=16'b1000100111001100;
    LogicCell40 \CLK_DDS.i19328_4_lut_LC_14_5_7  (
            .in0(N__34771),
            .in1(N__34620),
            .in2(N__44059),
            .in3(N__34464),
            .lcout(\CLK_DDS.n12784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i7_12189_12190_set_LC_14_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12189_12190_set_LC_14_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i7_12189_12190_set_LC_14_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_12189_12190_set_LC_14_6_0  (
            .in0(N__37343),
            .in1(N__44441),
            .in2(_gnd_net_),
            .in3(N__42386),
            .lcout(\comm_spi.n14607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52547),
            .ce(),
            .sr(N__35044));
    defparam comm_clear_301_LC_14_7_0.C_ON=1'b0;
    defparam comm_clear_301_LC_14_7_0.SEQ_MODE=4'b1000;
    defparam comm_clear_301_LC_14_7_0.LUT_INIT=16'b0111011100110011;
    LogicCell40 comm_clear_301_LC_14_7_0 (
            .in0(N__56958),
            .in1(N__51761),
            .in2(_gnd_net_),
            .in3(N__49489),
            .lcout(comm_clear),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54279),
            .ce(N__34866),
            .sr(_gnd_net_));
    defparam comm_index_i1_LC_14_8_0.C_ON=1'b0;
    defparam comm_index_i1_LC_14_8_0.SEQ_MODE=4'b1000;
    defparam comm_index_i1_LC_14_8_0.LUT_INIT=16'b1101111100100000;
    LogicCell40 comm_index_i1_LC_14_8_0 (
            .in0(N__49876),
            .in1(N__49965),
            .in2(N__50780),
            .in3(N__52355),
            .lcout(comm_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54282),
            .ce(N__36030),
            .sr(N__39429));
    defparam comm_index_i0_LC_14_8_1.C_ON=1'b0;
    defparam comm_index_i0_LC_14_8_1.SEQ_MODE=4'b1000;
    defparam comm_index_i0_LC_14_8_1.LUT_INIT=16'b1001100111001100;
    LogicCell40 comm_index_i0_LC_14_8_1 (
            .in0(N__49964),
            .in1(N__50733),
            .in2(_gnd_net_),
            .in3(N__49875),
            .lcout(comm_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54282),
            .ce(N__36030),
            .sr(N__39429));
    defparam comm_index_i2_LC_14_8_2.C_ON=1'b0;
    defparam comm_index_i2_LC_14_8_2.SEQ_MODE=4'b1000;
    defparam comm_index_i2_LC_14_8_2.LUT_INIT=16'b0110101010101010;
    LogicCell40 comm_index_i2_LC_14_8_2 (
            .in0(N__50578),
            .in1(N__52354),
            .in2(N__50781),
            .in3(N__49087),
            .lcout(comm_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54282),
            .ce(N__36030),
            .sr(N__39429));
    defparam i18512_4_lut_LC_14_9_0.C_ON=1'b0;
    defparam i18512_4_lut_LC_14_9_0.SEQ_MODE=4'b0000;
    defparam i18512_4_lut_LC_14_9_0.LUT_INIT=16'b1110111011110000;
    LogicCell40 i18512_4_lut_LC_14_9_0 (
            .in0(N__49171),
            .in1(N__52212),
            .in2(N__34875),
            .in3(N__55407),
            .lcout(),
            .ltout(n21122_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i0_LC_14_9_1.C_ON=1'b0;
    defparam comm_state_i0_LC_14_9_1.SEQ_MODE=4'b1000;
    defparam comm_state_i0_LC_14_9_1.LUT_INIT=16'b0101000011111010;
    LogicCell40 comm_state_i0_LC_14_9_1 (
            .in0(N__56826),
            .in1(_gnd_net_),
            .in2(N__34878),
            .in3(N__56544),
            .lcout(comm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54290),
            .ce(N__36981),
            .sr(_gnd_net_));
    defparam i18510_3_lut_LC_14_9_2.C_ON=1'b0;
    defparam i18510_3_lut_LC_14_9_2.SEQ_MODE=4'b0000;
    defparam i18510_3_lut_LC_14_9_2.LUT_INIT=16'b1110111001010101;
    LogicCell40 i18510_3_lut_LC_14_9_2 (
            .in0(N__49407),
            .in1(N__50008),
            .in2(_gnd_net_),
            .in3(N__51644),
            .lcout(n21120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_313_LC_14_9_3.C_ON=1'b0;
    defparam i2_2_lut_adj_313_LC_14_9_3.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_313_LC_14_9_3.LUT_INIT=16'b1010101011111111;
    LogicCell40 i2_2_lut_adj_313_LC_14_9_3 (
            .in0(N__50012),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49404),
            .lcout(n14529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_adj_271_LC_14_9_4.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_271_LC_14_9_4.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_271_LC_14_9_4.LUT_INIT=16'b1110111011111111;
    LogicCell40 i2_2_lut_3_lut_adj_271_LC_14_9_4 (
            .in0(N__49406),
            .in1(N__51643),
            .in2(_gnd_net_),
            .in3(N__56825),
            .lcout(n11361),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i22_4_lut_4_lut_LC_14_9_5.C_ON=1'b0;
    defparam i22_4_lut_4_lut_LC_14_9_5.SEQ_MODE=4'b0000;
    defparam i22_4_lut_4_lut_LC_14_9_5.LUT_INIT=16'b0101010100001000;
    LogicCell40 i22_4_lut_4_lut_LC_14_9_5 (
            .in0(N__51642),
            .in1(N__49849),
            .in2(N__50037),
            .in3(N__49405),
            .lcout(),
            .ltout(n7_adj_1616_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_219_LC_14_9_6.C_ON=1'b0;
    defparam i1_4_lut_adj_219_LC_14_9_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_219_LC_14_9_6.LUT_INIT=16'b1010101000100000;
    LogicCell40 i1_4_lut_adj_219_LC_14_9_6 (
            .in0(N__49562),
            .in1(N__55406),
            .in2(N__34857),
            .in3(N__56824),
            .lcout(n11896),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_valid_85_LC_14_10_0 .C_ON=1'b0;
    defparam \comm_spi.data_valid_85_LC_14_10_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_valid_85_LC_14_10_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.data_valid_85_LC_14_10_0  (
            .in0(N__35898),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35853),
            .lcout(comm_data_vld),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.data_valid_85C_net ),
            .ce(),
            .sr(N__55820));
    defparam \ADC_IAC.ADC_DATA_i13_LC_14_11_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i13_LC_14_11_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i13_LC_14_11_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i13_LC_14_11_0  (
            .in0(N__35807),
            .in1(N__35637),
            .in2(N__35250),
            .in3(N__53813),
            .lcout(buf_adcdata_iac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54307),
            .ce(),
            .sr(_gnd_net_));
    defparam i18514_4_lut_LC_14_11_1.C_ON=1'b0;
    defparam i18514_4_lut_LC_14_11_1.SEQ_MODE=4'b0000;
    defparam i18514_4_lut_LC_14_11_1.LUT_INIT=16'b0100010010100000;
    LogicCell40 i18514_4_lut_LC_14_11_1 (
            .in0(N__57385),
            .in1(N__35214),
            .in2(N__37698),
            .in3(N__54884),
            .lcout(n21124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19425_4_lut_3_lut_LC_14_11_2 .C_ON=1'b0;
    defparam \comm_spi.i19425_4_lut_3_lut_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19425_4_lut_3_lut_LC_14_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19425_4_lut_3_lut_LC_14_11_2  (
            .in0(N__35146),
            .in1(N__35065),
            .in2(_gnd_net_),
            .in3(N__55817),
            .lcout(\comm_spi.n14603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_11_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_11_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.RESET_I_0_100_2_lut_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__55816),
            .in2(_gnd_net_),
            .in3(N__35067),
            .lcout(\comm_spi.data_tx_7__N_774 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_14_11_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_14_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_92_2_lut_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__35066),
            .in2(_gnd_net_),
            .in3(N__55818),
            .lcout(\comm_spi.data_tx_7__N_766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i1_LC_14_11_5.C_ON=1'b0;
    defparam comm_buf_6__i1_LC_14_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i1_LC_14_11_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i1_LC_14_11_5 (
            .in0(N__39638),
            .in1(N__56831),
            .in2(N__45791),
            .in3(N__34997),
            .lcout(comm_buf_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54307),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i19_3_lut_LC_14_11_6.C_ON=1'b0;
    defparam mux_129_Mux_1_i19_3_lut_LC_14_11_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i19_3_lut_LC_14_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_1_i19_3_lut_LC_14_11_6 (
            .in0(N__34968),
            .in1(N__34937),
            .in2(_gnd_net_),
            .in3(N__57386),
            .lcout(n19_adj_1522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19445_4_lut_3_lut_LC_14_11_7 .C_ON=1'b0;
    defparam \comm_spi.i19445_4_lut_3_lut_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19445_4_lut_3_lut_LC_14_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.i19445_4_lut_3_lut_LC_14_11_7  (
            .in0(N__55819),
            .in1(N__39118),
            .in2(_gnd_net_),
            .in3(N__34901),
            .lcout(\comm_spi.n22875 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i2_LC_14_12_2.C_ON=1'b0;
    defparam buf_dds1_i2_LC_14_12_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i2_LC_14_12_2.LUT_INIT=16'b1101100000000000;
    LogicCell40 buf_dds1_i2_LC_14_12_2 (
            .in0(N__44908),
            .in1(N__48084),
            .in2(N__46891),
            .in3(N__40636),
            .lcout(buf_dds1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54320),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_51_LC_14_12_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_51_LC_14_12_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_51_LC_14_12_3.LUT_INIT=16'b0001000011111111;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_51_LC_14_12_3 (
            .in0(N__55522),
            .in1(N__51858),
            .in2(N__57109),
            .in3(N__44907),
            .lcout(n16891),
            .ltout(n16891_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i9_LC_14_12_4.C_ON=1'b0;
    defparam buf_dds1_i9_LC_14_12_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i9_LC_14_12_4.LUT_INIT=16'b1101000010000000;
    LogicCell40 buf_dds1_i9_LC_14_12_4 (
            .in0(N__44909),
            .in1(N__40119),
            .in2(N__36000),
            .in3(N__40237),
            .lcout(buf_dds1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54320),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19009_2_lut_LC_14_12_5 .C_ON=1'b0;
    defparam \SIG_DDS.i19009_2_lut_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19009_2_lut_LC_14_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \SIG_DDS.i19009_2_lut_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__43188),
            .in2(_gnd_net_),
            .in3(N__42286),
            .lcout(\SIG_DDS.n21571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i19_3_lut_LC_14_12_6.C_ON=1'b0;
    defparam mux_129_Mux_2_i19_3_lut_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i19_3_lut_LC_14_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_2_i19_3_lut_LC_14_12_6 (
            .in0(N__35982),
            .in1(N__35947),
            .in2(_gnd_net_),
            .in3(N__57499),
            .lcout(n19_adj_1518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i2_LC_14_12_7.C_ON=1'b0;
    defparam comm_cmd_i2_LC_14_12_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i2_LC_14_12_7.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i2_LC_14_12_7 (
            .in0(N__46078),
            .in1(N__45998),
            .in2(N__47224),
            .in3(N__53670),
            .lcout(comm_cmd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54320),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_response_302_LC_14_13_0.C_ON=1'b0;
    defparam comm_response_302_LC_14_13_0.SEQ_MODE=4'b1000;
    defparam comm_response_302_LC_14_13_0.LUT_INIT=16'b0000010100110000;
    LogicCell40 comm_response_302_LC_14_13_0 (
            .in0(N__49485),
            .in1(N__55525),
            .in2(N__57028),
            .in3(N__51826),
            .lcout(ICE_GPMI_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54333),
            .ce(N__35907),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_292_LC_14_13_1.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_292_LC_14_13_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_292_LC_14_13_1.LUT_INIT=16'b1101110111010000;
    LogicCell40 i1_3_lut_4_lut_adj_292_LC_14_13_1 (
            .in0(N__55524),
            .in1(N__56901),
            .in2(N__49591),
            .in3(N__49484),
            .lcout(n11385),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i17_3_lut_3_lut_LC_14_13_2.C_ON=1'b0;
    defparam i17_3_lut_3_lut_LC_14_13_2.SEQ_MODE=4'b0000;
    defparam i17_3_lut_3_lut_LC_14_13_2.LUT_INIT=16'b0100010000100010;
    LogicCell40 i17_3_lut_3_lut_LC_14_13_2 (
            .in0(N__49483),
            .in1(N__55523),
            .in2(_gnd_net_),
            .in3(N__51825),
            .lcout(),
            .ltout(n10_adj_1554_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_261_LC_14_13_3.C_ON=1'b0;
    defparam i1_3_lut_adj_261_LC_14_13_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_261_LC_14_13_3.LUT_INIT=16'b1010101010100000;
    LogicCell40 i1_3_lut_adj_261_LC_14_13_3 (
            .in0(N__49575),
            .in1(_gnd_net_),
            .in2(N__36033),
            .in3(N__56900),
            .lcout(n11850),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_241_LC_14_13_4.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_241_LC_14_13_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_241_LC_14_13_4.LUT_INIT=16'b1111111111111011;
    LogicCell40 i1_2_lut_4_lut_adj_241_LC_14_13_4 (
            .in0(N__54913),
            .in1(N__57498),
            .in2(N__41532),
            .in3(N__53548),
            .lcout(n20914),
            .ltout(n20914_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_226_LC_14_13_5.C_ON=1'b0;
    defparam i1_4_lut_adj_226_LC_14_13_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_226_LC_14_13_5.LUT_INIT=16'b1010111100100011;
    LogicCell40 i1_4_lut_adj_226_LC_14_13_5 (
            .in0(N__49574),
            .in1(N__36015),
            .in2(N__36018),
            .in3(N__56899),
            .lcout(n11819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18404_2_lut_3_lut_LC_14_13_7.C_ON=1'b0;
    defparam i18404_2_lut_3_lut_LC_14_13_7.SEQ_MODE=4'b0000;
    defparam i18404_2_lut_3_lut_LC_14_13_7.LUT_INIT=16'b1111111111101110;
    LogicCell40 i18404_2_lut_3_lut_LC_14_13_7 (
            .in0(N__51824),
            .in1(N__55500),
            .in2(_gnd_net_),
            .in3(N__49482),
            .lcout(n21014),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i0_LC_14_14_0.C_ON=1'b0;
    defparam req_data_cnt_i0_LC_14_14_0.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i0_LC_14_14_0.LUT_INIT=16'b1101100011011000;
    LogicCell40 req_data_cnt_i0_LC_14_14_0 (
            .in0(N__41723),
            .in1(N__37614),
            .in2(N__43334),
            .in3(_gnd_net_),
            .lcout(req_data_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54347),
            .ce(),
            .sr(_gnd_net_));
    defparam i15327_2_lut_3_lut_LC_14_14_1.C_ON=1'b0;
    defparam i15327_2_lut_3_lut_LC_14_14_1.SEQ_MODE=4'b0000;
    defparam i15327_2_lut_3_lut_LC_14_14_1.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15327_2_lut_3_lut_LC_14_14_1 (
            .in0(N__55550),
            .in1(N__51428),
            .in2(_gnd_net_),
            .in3(N__51862),
            .lcout(n14_adj_1584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_186_LC_14_14_2.C_ON=1'b0;
    defparam i1_4_lut_adj_186_LC_14_14_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_186_LC_14_14_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_186_LC_14_14_2 (
            .in0(N__46511),
            .in1(N__43391),
            .in2(N__43333),
            .in3(N__40777),
            .lcout(n17_adj_1489),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15344_2_lut_3_lut_LC_14_14_3.C_ON=1'b0;
    defparam i15344_2_lut_3_lut_LC_14_14_3.SEQ_MODE=4'b0000;
    defparam i15344_2_lut_3_lut_LC_14_14_3.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15344_2_lut_3_lut_LC_14_14_3 (
            .in0(N__55551),
            .in1(N__48068),
            .in2(_gnd_net_),
            .in3(N__51863),
            .lcout(n14_adj_1555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_251_LC_14_14_4.C_ON=1'b0;
    defparam i1_3_lut_adj_251_LC_14_14_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_251_LC_14_14_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_3_lut_adj_251_LC_14_14_4 (
            .in0(N__54554),
            .in1(N__49481),
            .in2(_gnd_net_),
            .in3(N__37645),
            .lcout(n20912),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15346_2_lut_3_lut_LC_14_14_5.C_ON=1'b0;
    defparam i15346_2_lut_3_lut_LC_14_14_5.SEQ_MODE=4'b0000;
    defparam i15346_2_lut_3_lut_LC_14_14_5.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15346_2_lut_3_lut_LC_14_14_5 (
            .in0(N__55549),
            .in1(N__42770),
            .in2(_gnd_net_),
            .in3(N__51861),
            .lcout(n14_adj_1549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i5_LC_14_14_6.C_ON=1'b0;
    defparam comm_cmd_i5_LC_14_14_6.SEQ_MODE=4'b1000;
    defparam comm_cmd_i5_LC_14_14_6.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i5_LC_14_14_6 (
            .in0(N__46081),
            .in1(N__46008),
            .in2(N__52125),
            .in3(N__49700),
            .lcout(comm_cmd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54347),
            .ce(),
            .sr(_gnd_net_));
    defparam i15385_2_lut_3_lut_LC_14_14_7.C_ON=1'b0;
    defparam i15385_2_lut_3_lut_LC_14_14_7.SEQ_MODE=4'b0000;
    defparam i15385_2_lut_3_lut_LC_14_14_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15385_2_lut_3_lut_LC_14_14_7 (
            .in0(N__55552),
            .in1(N__43292),
            .in2(_gnd_net_),
            .in3(N__51864),
            .lcout(n14_adj_1533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i12_LC_14_15_0.C_ON=1'b0;
    defparam buf_dds1_i12_LC_14_15_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i12_LC_14_15_0.LUT_INIT=16'b1100000010001000;
    LogicCell40 buf_dds1_i12_LC_14_15_0 (
            .in0(N__40309),
            .in1(N__40655),
            .in2(N__41492),
            .in3(N__44947),
            .lcout(buf_dds1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54360),
            .ce(),
            .sr(_gnd_net_));
    defparam i19064_2_lut_LC_14_15_1.C_ON=1'b0;
    defparam i19064_2_lut_LC_14_15_1.SEQ_MODE=4'b0000;
    defparam i19064_2_lut_LC_14_15_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19064_2_lut_LC_14_15_1 (
            .in0(_gnd_net_),
            .in1(N__57661),
            .in2(_gnd_net_),
            .in3(N__36055),
            .lcout(n21286),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i14_LC_14_15_2.C_ON=1'b0;
    defparam req_data_cnt_i14_LC_14_15_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i14_LC_14_15_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i14_LC_14_15_2 (
            .in0(N__36056),
            .in1(N__38070),
            .in2(_gnd_net_),
            .in3(N__41725),
            .lcout(req_data_cnt_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54360),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19372_4_lut_LC_14_15_4 .C_ON=1'b0;
    defparam \SIG_DDS.i19372_4_lut_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19372_4_lut_LC_14_15_4 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \SIG_DDS.i19372_4_lut_LC_14_15_4  (
            .in0(N__42131),
            .in1(N__41311),
            .in2(N__43059),
            .in3(N__42266),
            .lcout(\SIG_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i7_LC_14_15_5.C_ON=1'b0;
    defparam req_data_cnt_i7_LC_14_15_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i7_LC_14_15_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 req_data_cnt_i7_LC_14_15_5 (
            .in0(_gnd_net_),
            .in1(N__46993),
            .in2(N__41739),
            .in3(N__37878),
            .lcout(req_data_cnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54360),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_174_LC_14_15_6.C_ON=1'b0;
    defparam i6_4_lut_adj_174_LC_14_15_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_174_LC_14_15_6.LUT_INIT=16'b0111110110111110;
    LogicCell40 i6_4_lut_adj_174_LC_14_15_6 (
            .in0(N__47122),
            .in1(N__50452),
            .in2(N__46997),
            .in3(N__46603),
            .lcout(n22_adj_1499),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_182_LC_14_16_0.C_ON=1'b0;
    defparam i2_4_lut_adj_182_LC_14_16_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_182_LC_14_16_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_182_LC_14_16_0 (
            .in0(N__37918),
            .in1(N__46192),
            .in2(N__46817),
            .in3(N__37081),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_177_LC_14_16_1.C_ON=1'b0;
    defparam i7_4_lut_adj_177_LC_14_16_1.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_177_LC_14_16_1.LUT_INIT=16'b0111101111011110;
    LogicCell40 i7_4_lut_adj_177_LC_14_16_1 (
            .in0(N__38105),
            .in1(N__40936),
            .in2(N__36060),
            .in3(N__41020),
            .lcout(n23_adj_1614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i10_LC_14_16_2.C_ON=1'b0;
    defparam req_data_cnt_i10_LC_14_16_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i10_LC_14_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i10_LC_14_16_2 (
            .in0(N__37790),
            .in1(N__41702),
            .in2(_gnd_net_),
            .in3(N__40813),
            .lcout(req_data_cnt_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54373),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i11_LC_14_16_3.C_ON=1'b0;
    defparam req_data_cnt_i11_LC_14_16_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i11_LC_14_16_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i11_LC_14_16_3 (
            .in0(N__41703),
            .in1(N__44427),
            .in2(_gnd_net_),
            .in3(N__41021),
            .lcout(req_data_cnt_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54373),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_130_LC_14_16_4.C_ON=1'b0;
    defparam i2_4_lut_adj_130_LC_14_16_4.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_130_LC_14_16_4.LUT_INIT=16'b0000000000010000;
    LogicCell40 i2_4_lut_adj_130_LC_14_16_4 (
            .in0(N__49426),
            .in1(N__47058),
            .in2(N__57108),
            .in3(N__36333),
            .lcout(n10520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i4_LC_14_16_5.C_ON=1'b0;
    defparam req_data_cnt_i4_LC_14_16_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i4_LC_14_16_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 req_data_cnt_i4_LC_14_16_5 (
            .in0(_gnd_net_),
            .in1(N__37526),
            .in2(N__41724),
            .in3(N__46813),
            .lcout(req_data_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54373),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i15_LC_14_16_6.C_ON=1'b0;
    defparam req_data_cnt_i15_LC_14_16_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i15_LC_14_16_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i15_LC_14_16_6 (
            .in0(N__38028),
            .in1(N__41704),
            .in2(_gnd_net_),
            .in3(N__36223),
            .lcout(req_data_cnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54373),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_267_LC_14_17_0.C_ON=1'b0;
    defparam i15_4_lut_adj_267_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_267_LC_14_17_0.LUT_INIT=16'b1100111101000111;
    LogicCell40 i15_4_lut_adj_267_LC_14_17_0 (
            .in0(N__47690),
            .in1(N__57014),
            .in2(N__36558),
            .in3(N__56228),
            .lcout(n12280),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4408_3_lut_LC_14_17_1.C_ON=1'b0;
    defparam i4408_3_lut_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam i4408_3_lut_LC_14_17_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i4408_3_lut_LC_14_17_1 (
            .in0(N__43283),
            .in1(N__36321),
            .in2(_gnd_net_),
            .in3(N__47689),
            .lcout(n8_adj_1532),
            .ltout(n8_adj_1532_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_14_17_2.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_14_17_2.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_14_17_2 (
            .in0(N__36302),
            .in1(N__56227),
            .in2(N__36204),
            .in3(N__57013),
            .lcout(data_index_9_N_216_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i0_LC_14_17_3.C_ON=1'b0;
    defparam data_index_i0_LC_14_17_3.SEQ_MODE=4'b1000;
    defparam data_index_i0_LC_14_17_3.LUT_INIT=16'b0100111001000100;
    LogicCell40 data_index_i0_LC_14_17_3 (
            .in0(N__57015),
            .in1(N__36303),
            .in2(N__56344),
            .in3(N__36102),
            .lcout(data_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54387),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_310_LC_14_17_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_310_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_310_LC_14_17_4.LUT_INIT=16'b1111111101110111;
    LogicCell40 i1_2_lut_3_lut_adj_310_LC_14_17_4 (
            .in0(N__57654),
            .in1(N__54747),
            .in2(_gnd_net_),
            .in3(N__37652),
            .lcout(n11338),
            .ltout(n11338_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_14_17_5.C_ON=1'b0;
    defparam i3_4_lut_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_14_17_5.LUT_INIT=16'b1111111011111111;
    LogicCell40 i3_4_lut_LC_14_17_5 (
            .in0(N__49425),
            .in1(N__55056),
            .in2(N__36327),
            .in3(N__53679),
            .lcout(n8813),
            .ltout(n8813_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6429_3_lut_LC_14_17_6.C_ON=1'b0;
    defparam i6429_3_lut_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam i6429_3_lut_LC_14_17_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 i6429_3_lut_LC_14_17_6 (
            .in0(_gnd_net_),
            .in1(N__51019),
            .in2(N__36324),
            .in3(N__41099),
            .lcout(n8_adj_1569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i5_LC_14_17_7.C_ON=1'b0;
    defparam req_data_cnt_i5_LC_14_17_7.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i5_LC_14_17_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i5_LC_14_17_7 (
            .in0(N__37497),
            .in1(N__41698),
            .in2(_gnd_net_),
            .in3(N__52844),
            .lcout(req_data_cnt_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54387),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_2_lut_LC_14_18_0.C_ON=1'b1;
    defparam add_125_2_lut_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam add_125_2_lut_LC_14_18_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_2_lut_LC_14_18_0 (
            .in0(N__36320),
            .in1(N__36319),
            .in2(N__36536),
            .in3(N__36291),
            .lcout(n7),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(n19625),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_3_lut_LC_14_18_1.C_ON=1'b1;
    defparam add_125_3_lut_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam add_125_3_lut_LC_14_18_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_3_lut_LC_14_18_1 (
            .in0(N__36287),
            .in1(N__36286),
            .in2(N__36559),
            .in3(N__36270),
            .lcout(n7_adj_1572),
            .ltout(),
            .carryin(n19625),
            .carryout(n19626),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_4_lut_LC_14_18_2.C_ON=1'b1;
    defparam add_125_4_lut_LC_14_18_2.SEQ_MODE=4'b0000;
    defparam add_125_4_lut_LC_14_18_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_4_lut_LC_14_18_2 (
            .in0(N__41004),
            .in1(N__41003),
            .in2(N__36537),
            .in3(N__36267),
            .lcout(n7_adj_1570),
            .ltout(),
            .carryin(n19626),
            .carryout(n19627),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_5_lut_LC_14_18_3.C_ON=1'b1;
    defparam add_125_5_lut_LC_14_18_3.SEQ_MODE=4'b0000;
    defparam add_125_5_lut_LC_14_18_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_5_lut_LC_14_18_3 (
            .in0(N__41100),
            .in1(N__41098),
            .in2(N__36560),
            .in3(N__36264),
            .lcout(n7_adj_1568),
            .ltout(),
            .carryin(n19627),
            .carryout(n19628),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_6_lut_LC_14_18_4.C_ON=1'b1;
    defparam add_125_6_lut_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam add_125_6_lut_LC_14_18_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_6_lut_LC_14_18_4 (
            .in0(N__47723),
            .in1(N__47722),
            .in2(N__36538),
            .in3(N__36261),
            .lcout(n7_adj_1566),
            .ltout(),
            .carryin(n19628),
            .carryout(n19629),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_7_lut_LC_14_18_5.C_ON=1'b1;
    defparam add_125_7_lut_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam add_125_7_lut_LC_14_18_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_7_lut_LC_14_18_5 (
            .in0(N__40569),
            .in1(N__40567),
            .in2(N__36561),
            .in3(N__36579),
            .lcout(n17487),
            .ltout(),
            .carryin(n19629),
            .carryout(n19630),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_8_lut_LC_14_18_6.C_ON=1'b1;
    defparam add_125_8_lut_LC_14_18_6.SEQ_MODE=4'b0000;
    defparam add_125_8_lut_LC_14_18_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_8_lut_LC_14_18_6 (
            .in0(N__38393),
            .in1(N__38392),
            .in2(N__36539),
            .in3(N__36576),
            .lcout(n7_adj_1564),
            .ltout(),
            .carryin(n19630),
            .carryout(n19631),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_9_lut_LC_14_18_7.C_ON=1'b1;
    defparam add_125_9_lut_LC_14_18_7.SEQ_MODE=4'b0000;
    defparam add_125_9_lut_LC_14_18_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_9_lut_LC_14_18_7 (
            .in0(N__41991),
            .in1(N__41990),
            .in2(N__36562),
            .in3(N__36573),
            .lcout(n7_adj_1562),
            .ltout(),
            .carryin(n19631),
            .carryout(n19632),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_10_lut_LC_14_19_0.C_ON=1'b1;
    defparam add_125_10_lut_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam add_125_10_lut_LC_14_19_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_10_lut_LC_14_19_0 (
            .in0(N__42062),
            .in1(N__42058),
            .in2(N__36567),
            .in3(N__36570),
            .lcout(n7_adj_1560),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(n19633),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_11_lut_LC_14_19_1.C_ON=1'b0;
    defparam add_125_11_lut_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam add_125_11_lut_LC_14_19_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_11_lut_LC_14_19_1 (
            .in0(N__39076),
            .in1(N__39077),
            .in2(N__36566),
            .in3(N__36480),
            .lcout(n7_adj_1558),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i8_LC_14_19_2.C_ON=1'b0;
    defparam data_index_i8_LC_14_19_2.SEQ_MODE=4'b1000;
    defparam data_index_i8_LC_14_19_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i8_LC_14_19_2 (
            .in0(N__57059),
            .in1(N__42042),
            .in2(N__56473),
            .in3(N__38952),
            .lcout(data_index_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54414),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i3_LC_14_19_3.C_ON=1'b0;
    defparam buf_control_i3_LC_14_19_3.SEQ_MODE=4'b1000;
    defparam buf_control_i3_LC_14_19_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i3_LC_14_19_3 (
            .in0(N__56357),
            .in1(N__41887),
            .in2(N__44228),
            .in3(N__41953),
            .lcout(SELIRNG1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54414),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4.LUT_INIT=16'b0010111000100010;
    LogicCell40 comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4 (
            .in0(N__36476),
            .in1(N__57090),
            .in2(N__56472),
            .in3(N__36465),
            .lcout(data_index_9_N_216_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i1_LC_14_19_5.C_ON=1'b0;
    defparam buf_control_i1_LC_14_19_5.SEQ_MODE=4'b1000;
    defparam buf_control_i1_LC_14_19_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i1_LC_14_19_5 (
            .in0(N__56356),
            .in1(N__41886),
            .in2(N__40155),
            .in3(N__36352),
            .lcout(DDS_RNG_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54414),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.MOSI_31_LC_14_19_6 .C_ON=1'b0;
    defparam \SIG_DDS.MOSI_31_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.MOSI_31_LC_14_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \SIG_DDS.MOSI_31_LC_14_19_6  (
            .in0(N__36780),
            .in1(N__36752),
            .in2(_gnd_net_),
            .in3(N__42976),
            .lcout(DDS_MOSI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54414),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i9_LC_14_19_7.C_ON=1'b0;
    defparam data_index_i9_LC_14_19_7.SEQ_MODE=4'b1000;
    defparam data_index_i9_LC_14_19_7.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i9_LC_14_19_7 (
            .in0(N__39060),
            .in1(N__57060),
            .in2(N__56476),
            .in3(N__39054),
            .lcout(data_index_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54414),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.CS_28_LC_14_20_1 .C_ON=1'b0;
    defparam \SIG_DDS.CS_28_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.CS_28_LC_14_20_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \SIG_DDS.CS_28_LC_14_20_1  (
            .in0(N__42196),
            .in1(N__42983),
            .in2(_gnd_net_),
            .in3(N__41335),
            .lcout(DDS_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54421),
            .ce(N__36720),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i2_12204_12205_reset_LC_15_2_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12204_12205_reset_LC_15_2_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i2_12204_12205_reset_LC_15_2_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12204_12205_reset_LC_15_2_0  (
            .in0(N__39344),
            .in1(N__38573),
            .in2(_gnd_net_),
            .in3(N__38618),
            .lcout(\comm_spi.n14623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52641),
            .ce(),
            .sr(N__39321));
    defparam \comm_spi.data_tx_i0_12174_12175_reset_LC_15_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12174_12175_reset_LC_15_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i0_12174_12175_reset_LC_15_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_12174_12175_reset_LC_15_3_0  (
            .in0(N__58335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52639),
            .ce(),
            .sr(N__36714));
    defparam \ADC_VDC.bit_cnt_3769__i0_LC_15_4_0 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i0_LC_15_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i0_LC_15_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i0_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__36705),
            .in2(_gnd_net_),
            .in3(N__36672),
            .lcout(\ADC_VDC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\ADC_VDC.n19772 ),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam \ADC_VDC.bit_cnt_3769__i1_LC_15_4_1 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i1_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i1_LC_15_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i1_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__36669),
            .in2(_gnd_net_),
            .in3(N__36648),
            .lcout(\ADC_VDC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19772 ),
            .carryout(\ADC_VDC.n19773 ),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam \ADC_VDC.bit_cnt_3769__i2_LC_15_4_2 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i2_LC_15_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i2_LC_15_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i2_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__36644),
            .in2(_gnd_net_),
            .in3(N__36615),
            .lcout(\ADC_VDC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19773 ),
            .carryout(\ADC_VDC.n19774 ),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam \ADC_VDC.bit_cnt_3769__i3_LC_15_4_3 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i3_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i3_LC_15_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i3_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__36610),
            .in2(_gnd_net_),
            .in3(N__36582),
            .lcout(\ADC_VDC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19774 ),
            .carryout(\ADC_VDC.n19775 ),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam \ADC_VDC.bit_cnt_3769__i4_LC_15_4_4 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i4_LC_15_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i4_LC_15_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i4_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(N__36913),
            .in2(_gnd_net_),
            .in3(N__36885),
            .lcout(\ADC_VDC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19775 ),
            .carryout(\ADC_VDC.n19776 ),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam \ADC_VDC.bit_cnt_3769__i5_LC_15_4_5 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i5_LC_15_4_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i5_LC_15_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i5_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__36881),
            .in2(_gnd_net_),
            .in3(N__36858),
            .lcout(\ADC_VDC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19776 ),
            .carryout(\ADC_VDC.n19777 ),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam \ADC_VDC.bit_cnt_3769__i6_LC_15_4_6 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i6_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i6_LC_15_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i6_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__36855),
            .in2(_gnd_net_),
            .in3(N__36834),
            .lcout(\ADC_VDC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19777 ),
            .carryout(\ADC_VDC.n19778 ),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam \ADC_VDC.bit_cnt_3769__i7_LC_15_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.bit_cnt_3769__i7_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i7_LC_15_4_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i7_LC_15_4_7  (
            .in0(_gnd_net_),
            .in1(N__36828),
            .in2(_gnd_net_),
            .in3(N__36831),
            .lcout(\ADC_VDC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53194),
            .ce(N__47508),
            .sr(N__36804));
    defparam wdtick_flag_289_LC_15_5_0.C_ON=1'b0;
    defparam wdtick_flag_289_LC_15_5_0.SEQ_MODE=4'b1010;
    defparam wdtick_flag_289_LC_15_5_0.LUT_INIT=16'b1111111100010000;
    LogicCell40 wdtick_flag_289_LC_15_5_0 (
            .in0(N__39245),
            .in1(N__39225),
            .in2(N__39264),
            .in3(N__44633),
            .lcout(wdtick_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39205),
            .ce(),
            .sr(N__39417));
    defparam \comm_spi.data_tx_i4_12212_12213_reset_LC_15_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12212_12213_reset_LC_15_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i4_12212_12213_reset_LC_15_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_12212_12213_reset_LC_15_6_0  (
            .in0(N__39131),
            .in1(N__39095),
            .in2(_gnd_net_),
            .in3(N__39146),
            .lcout(\comm_spi.n14631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52548),
            .ce(),
            .sr(N__39492));
    defparam \comm_spi.data_tx_i3_12208_12209_reset_LC_15_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12208_12209_reset_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i3_12208_12209_reset_LC_15_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_12208_12209_reset_LC_15_7_0  (
            .in0(N__39287),
            .in1(N__37359),
            .in2(_gnd_net_),
            .in3(N__37385),
            .lcout(\comm_spi.n14627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(),
            .sr(N__36795));
    defparam i2_3_lut_LC_15_8_0.C_ON=1'b0;
    defparam i2_3_lut_LC_15_8_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_15_8_0.LUT_INIT=16'b1110111011111111;
    LogicCell40 i2_3_lut_LC_15_8_0 (
            .in0(N__45861),
            .in1(N__36968),
            .in2(_gnd_net_),
            .in3(N__49086),
            .lcout(n19902),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_258_LC_15_8_1.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_258_LC_15_8_1.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_258_LC_15_8_1.LUT_INIT=16'b1111111011111111;
    LogicCell40 i2_3_lut_4_lut_adj_258_LC_15_8_1 (
            .in0(N__51645),
            .in1(N__49167),
            .in2(N__45878),
            .in3(N__49874),
            .lcout(),
            .ltout(n20944_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_15_8_2.C_ON=1'b0;
    defparam i2_4_lut_LC_15_8_2.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_15_8_2.LUT_INIT=16'b1110000000000000;
    LogicCell40 i2_4_lut_LC_15_8_2 (
            .in0(N__49654),
            .in1(N__36975),
            .in2(N__36984),
            .in3(N__36954),
            .lcout(n20964),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_4_lut_LC_15_8_3.C_ON=1'b0;
    defparam i3_4_lut_4_lut_LC_15_8_3.SEQ_MODE=4'b0000;
    defparam i3_4_lut_4_lut_LC_15_8_3.LUT_INIT=16'b0111011111110011;
    LogicCell40 i3_4_lut_4_lut_LC_15_8_3 (
            .in0(N__49409),
            .in1(N__51636),
            .in2(N__50031),
            .in3(N__49873),
            .lcout(n20962),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_317_LC_15_8_4.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_317_LC_15_8_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_317_LC_15_8_4.LUT_INIT=16'b0111111100101111;
    LogicCell40 i1_4_lut_4_lut_adj_317_LC_15_8_4 (
            .in0(N__49872),
            .in1(N__49408),
            .in2(N__51759),
            .in3(N__49994),
            .lcout(n4_adj_1586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_298_LC_15_8_5.C_ON=1'b0;
    defparam i2_4_lut_adj_298_LC_15_8_5.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_298_LC_15_8_5.LUT_INIT=16'b1110111100000000;
    LogicCell40 i2_4_lut_adj_298_LC_15_8_5 (
            .in0(N__36969),
            .in1(N__49653),
            .in2(N__50030),
            .in3(N__37035),
            .lcout(n20801),
            .ltout(n20801_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_15_8_6.C_ON=1'b0;
    defparam i1_4_lut_LC_15_8_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_15_8_6.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_LC_15_8_6 (
            .in0(N__49655),
            .in1(N__36948),
            .in2(N__36942),
            .in3(N__36939),
            .lcout(n20829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19129_2_lut_3_lut_LC_15_8_7.C_ON=1'b0;
    defparam i19129_2_lut_3_lut_LC_15_8_7.SEQ_MODE=4'b0000;
    defparam i19129_2_lut_3_lut_LC_15_8_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i19129_2_lut_3_lut_LC_15_8_7 (
            .in0(N__49993),
            .in1(N__51632),
            .in2(_gnd_net_),
            .in3(N__49871),
            .lcout(n21369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_1__bdd_4_lut_LC_15_9_0.C_ON=1'b0;
    defparam comm_state_1__bdd_4_lut_LC_15_9_0.SEQ_MODE=4'b0000;
    defparam comm_state_1__bdd_4_lut_LC_15_9_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_state_1__bdd_4_lut_LC_15_9_0 (
            .in0(N__37626),
            .in1(N__51637),
            .in2(N__49172),
            .in3(N__55404),
            .lcout(n22423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_15_9_1.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_15_9_1.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_15_9_1.LUT_INIT=16'b0011000010111000;
    LogicCell40 comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_15_9_1 (
            .in0(N__51641),
            .in1(N__49412),
            .in2(N__50047),
            .in3(N__37028),
            .lcout(),
            .ltout(n2_adj_1581_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22423_bdd_4_lut_LC_15_9_2.C_ON=1'b0;
    defparam n22423_bdd_4_lut_LC_15_9_2.SEQ_MODE=4'b0000;
    defparam n22423_bdd_4_lut_LC_15_9_2.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22423_bdd_4_lut_LC_15_9_2 (
            .in0(N__49413),
            .in1(N__36933),
            .in2(N__36924),
            .in3(N__55405),
            .lcout(n22426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19296_4_lut_LC_15_9_3.C_ON=1'b0;
    defparam i19296_4_lut_LC_15_9_3.SEQ_MODE=4'b0000;
    defparam i19296_4_lut_LC_15_9_3.LUT_INIT=16'b0000111000000010;
    LogicCell40 i19296_4_lut_LC_15_9_3 (
            .in0(N__50035),
            .in1(N__55451),
            .in2(N__51760),
            .in3(N__49088),
            .lcout(),
            .ltout(n21370_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19388_4_lut_LC_15_9_4.C_ON=1'b0;
    defparam i19388_4_lut_LC_15_9_4.SEQ_MODE=4'b0000;
    defparam i19388_4_lut_LC_15_9_4.LUT_INIT=16'b1100111011011111;
    LogicCell40 i19388_4_lut_LC_15_9_4 (
            .in0(N__49411),
            .in1(N__56822),
            .in2(N__37065),
            .in3(N__37062),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i1_LC_15_9_5.C_ON=1'b0;
    defparam comm_state_i1_LC_15_9_5.SEQ_MODE=4'b1000;
    defparam comm_state_i1_LC_15_9_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_i1_LC_15_9_5 (
            .in0(N__56823),
            .in1(N__37017),
            .in2(N__56567),
            .in3(N__37056),
            .lcout(comm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54296),
            .ce(N__37050),
            .sr(_gnd_net_));
    defparam i227_2_lut_LC_15_9_6.C_ON=1'b0;
    defparam i227_2_lut_LC_15_9_6.SEQ_MODE=4'b0000;
    defparam i227_2_lut_LC_15_9_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 i227_2_lut_LC_15_9_6 (
            .in0(_gnd_net_),
            .in1(N__50036),
            .in2(_gnd_net_),
            .in3(N__49848),
            .lcout(n1264),
            .ltout(n1264_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_296_LC_15_9_7.C_ON=1'b0;
    defparam i1_4_lut_adj_296_LC_15_9_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_296_LC_15_9_7.LUT_INIT=16'b1111101100000000;
    LogicCell40 i1_4_lut_adj_296_LC_15_9_7 (
            .in0(N__49566),
            .in1(N__49410),
            .in2(N__37038),
            .in3(N__37215),
            .lcout(n4_adj_1643),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_15_10_0.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_15_10_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_15_10_0.LUT_INIT=16'b0000001110001011;
    LogicCell40 comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_15_10_0 (
            .in0(N__51574),
            .in1(N__49402),
            .in2(N__37011),
            .in3(N__37029),
            .lcout(n8_adj_1582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_84_LC_15_10_1.C_ON=1'b0;
    defparam i1_4_lut_adj_84_LC_15_10_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_84_LC_15_10_1.LUT_INIT=16'b1100000011000100;
    LogicCell40 i1_4_lut_adj_84_LC_15_10_1 (
            .in0(N__55136),
            .in1(N__45666),
            .in2(N__40038),
            .in3(N__53671),
            .lcout(comm_state_3_N_420_3),
            .ltout(comm_state_3_N_420_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19114_2_lut_LC_15_10_2.C_ON=1'b0;
    defparam i19114_2_lut_LC_15_10_2.SEQ_MODE=4'b0000;
    defparam i19114_2_lut_LC_15_10_2.LUT_INIT=16'b0000000011110000;
    LogicCell40 i19114_2_lut_LC_15_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37002),
            .in3(N__49403),
            .lcout(),
            .ltout(n21435_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i3_LC_15_10_3.C_ON=1'b0;
    defparam comm_state_i3_LC_15_10_3.SEQ_MODE=4'b1000;
    defparam comm_state_i3_LC_15_10_3.LUT_INIT=16'b0010000001110101;
    LogicCell40 comm_state_i3_LC_15_10_3 (
            .in0(N__56830),
            .in1(N__56452),
            .in2(N__36999),
            .in3(N__49143),
            .lcout(comm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54308),
            .ce(N__36996),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_275_LC_15_10_4.C_ON=1'b0;
    defparam i1_2_lut_adj_275_LC_15_10_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_275_LC_15_10_4.LUT_INIT=16'b1111111101010101;
    LogicCell40 i1_2_lut_adj_275_LC_15_10_4 (
            .in0(N__51573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49401),
            .lcout(),
            .ltout(n20937_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_268_LC_15_10_5.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_268_LC_15_10_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_268_LC_15_10_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i2_3_lut_4_lut_adj_268_LC_15_10_5 (
            .in0(N__50045),
            .in1(N__49847),
            .in2(N__37218),
            .in3(N__45846),
            .lcout(n20939),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_101_LC_15_10_6.C_ON=1'b0;
    defparam i1_2_lut_adj_101_LC_15_10_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_101_LC_15_10_6.LUT_INIT=16'b1010101011111111;
    LogicCell40 i1_2_lut_adj_101_LC_15_10_6 (
            .in0(N__56693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55430),
            .lcout(n20917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_311_LC_15_10_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_311_LC_15_10_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_311_LC_15_10_7.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_311_LC_15_10_7 (
            .in0(N__55429),
            .in1(N__56692),
            .in2(_gnd_net_),
            .in3(N__51572),
            .lcout(n12226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19644_LC_15_11_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19644_LC_15_11_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19644_LC_15_11_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19644_LC_15_11_0 (
            .in0(N__37209),
            .in1(N__55140),
            .in2(N__37203),
            .in3(N__53552),
            .lcout(),
            .ltout(n22261_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22261_bdd_4_lut_LC_15_11_1.C_ON=1'b0;
    defparam n22261_bdd_4_lut_LC_15_11_1.SEQ_MODE=4'b0000;
    defparam n22261_bdd_4_lut_LC_15_11_1.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22261_bdd_4_lut_LC_15_11_1 (
            .in0(N__53553),
            .in1(N__37172),
            .in2(N__37140),
            .in3(N__37137),
            .lcout(n22264),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i26_3_lut_LC_15_11_2.C_ON=1'b0;
    defparam mux_129_Mux_1_i26_3_lut_LC_15_11_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i26_3_lut_LC_15_11_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_129_Mux_1_i26_3_lut_LC_15_11_2 (
            .in0(N__57477),
            .in1(_gnd_net_),
            .in2(N__37575),
            .in3(N__37923),
            .lcout(),
            .ltout(n26_adj_1523_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19773_LC_15_11_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19773_LC_15_11_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19773_LC_15_11_3.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19773_LC_15_11_3 (
            .in0(N__53554),
            .in1(N__55059),
            .in2(N__37125),
            .in3(N__57156),
            .lcout(),
            .ltout(n22411_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22411_bdd_4_lut_LC_15_11_4.C_ON=1'b0;
    defparam n22411_bdd_4_lut_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam n22411_bdd_4_lut_LC_15_11_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22411_bdd_4_lut_LC_15_11_4 (
            .in0(N__53555),
            .in1(N__37122),
            .in2(N__37095),
            .in3(N__37092),
            .lcout(),
            .ltout(n22414_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1553761_i1_3_lut_LC_15_11_5.C_ON=1'b0;
    defparam i1553761_i1_3_lut_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam i1553761_i1_3_lut_LC_15_11_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1553761_i1_3_lut_LC_15_11_5 (
            .in0(_gnd_net_),
            .in1(N__37467),
            .in2(N__37461),
            .in3(N__54745),
            .lcout(),
            .ltout(n30_adj_1524_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i1_LC_15_11_6.C_ON=1'b0;
    defparam comm_buf_1__i1_LC_15_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i1_LC_15_11_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i1_LC_15_11_6 (
            .in0(_gnd_net_),
            .in1(N__45768),
            .in2(N__37458),
            .in3(N__51758),
            .lcout(comm_buf_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54321),
            .ce(N__51383),
            .sr(N__51302));
    defparam \comm_spi.data_tx_i3_12208_12209_set_LC_15_12_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12208_12209_set_LC_15_12_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i3_12208_12209_set_LC_15_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_12208_12209_set_LC_15_12_0  (
            .in0(N__39291),
            .in1(N__37355),
            .in2(_gnd_net_),
            .in3(N__37389),
            .lcout(\comm_spi.n14626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52638),
            .ce(),
            .sr(N__37371));
    defparam i19037_2_lut_LC_15_12_2.C_ON=1'b0;
    defparam i19037_2_lut_LC_15_12_2.SEQ_MODE=4'b0000;
    defparam i19037_2_lut_LC_15_12_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 i19037_2_lut_LC_15_12_2 (
            .in0(N__57701),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38048),
            .lcout(n21272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19106_2_lut_LC_15_12_5.C_ON=1'b0;
    defparam i19106_2_lut_LC_15_12_5.SEQ_MODE=4'b0000;
    defparam i19106_2_lut_LC_15_12_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i19106_2_lut_LC_15_12_5 (
            .in0(_gnd_net_),
            .in1(N__37748),
            .in2(_gnd_net_),
            .in3(N__57700),
            .lcout(n21568),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i2_12204_12205_set_LC_15_13_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12204_12205_set_LC_15_13_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i2_12204_12205_set_LC_15_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_tx_i2_12204_12205_set_LC_15_13_0  (
            .in0(N__38580),
            .in1(N__39351),
            .in2(_gnd_net_),
            .in3(N__38628),
            .lcout(\comm_spi.n14622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52609),
            .ce(),
            .sr(N__39309));
    defparam \comm_spi.i19450_4_lut_3_lut_LC_15_13_1 .C_ON=1'b0;
    defparam \comm_spi.i19450_4_lut_3_lut_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19450_4_lut_3_lut_LC_15_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.i19450_4_lut_3_lut_LC_15_13_1  (
            .in0(N__55874),
            .in1(N__44546),
            .in2(_gnd_net_),
            .in3(N__39483),
            .lcout(\comm_spi.n22872 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19460_4_lut_3_lut_LC_15_13_3 .C_ON=1'b0;
    defparam \comm_spi.i19460_4_lut_3_lut_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19460_4_lut_3_lut_LC_15_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.i19460_4_lut_3_lut_LC_15_13_3  (
            .in0(N__37328),
            .in1(N__55875),
            .in2(_gnd_net_),
            .in3(N__45270),
            .lcout(\comm_spi.n22857 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12225_2_lut_LC_15_13_4.C_ON=1'b0;
    defparam i12225_2_lut_LC_15_13_4.SEQ_MODE=4'b0000;
    defparam i12225_2_lut_LC_15_13_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 i12225_2_lut_LC_15_13_4 (
            .in0(_gnd_net_),
            .in1(N__37316),
            .in2(_gnd_net_),
            .in3(N__38556),
            .lcout(n14647),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i17178_2_lut_LC_15_13_5.C_ON=1'b0;
    defparam i17178_2_lut_LC_15_13_5.SEQ_MODE=4'b0000;
    defparam i17178_2_lut_LC_15_13_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i17178_2_lut_LC_15_13_5 (
            .in0(_gnd_net_),
            .in1(N__50579),
            .in2(_gnd_net_),
            .in3(N__49497),
            .lcout(n19783),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_211_LC_15_13_6.C_ON=1'b0;
    defparam i1_2_lut_adj_211_LC_15_13_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_211_LC_15_13_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 i1_2_lut_adj_211_LC_15_13_6 (
            .in0(N__49498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50580),
            .lcout(n26_adj_1644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19281_2_lut_LC_15_13_7.C_ON=1'b0;
    defparam i19281_2_lut_LC_15_13_7.SEQ_MODE=4'b0000;
    defparam i19281_2_lut_LC_15_13_7.LUT_INIT=16'b1111111111001100;
    LogicCell40 i19281_2_lut_LC_15_13_7 (
            .in0(_gnd_net_),
            .in1(N__49499),
            .in2(_gnd_net_),
            .in3(N__37656),
            .lcout(n21521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_idxvec_i0_LC_15_14_0.C_ON=1'b1;
    defparam data_idxvec_i0_LC_15_14_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i0_LC_15_14_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i0_LC_15_14_0 (
            .in0(N__37613),
            .in1(N__56929),
            .in2(N__43412),
            .in3(N__37602),
            .lcout(data_idxvec_0),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(n19634),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i1_LC_15_14_1.C_ON=1'b1;
    defparam data_idxvec_i1_LC_15_14_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i1_LC_15_14_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i1_LC_15_14_1 (
            .in0(N__37599),
            .in1(N__56933),
            .in2(N__37574),
            .in3(N__37554),
            .lcout(data_idxvec_1),
            .ltout(),
            .carryin(n19634),
            .carryout(n19635),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i2_LC_15_14_2.C_ON=1'b1;
    defparam data_idxvec_i2_LC_15_14_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i2_LC_15_14_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i2_LC_15_14_2 (
            .in0(N__37551),
            .in1(N__56930),
            .in2(N__47147),
            .in3(N__37533),
            .lcout(data_idxvec_2),
            .ltout(),
            .carryin(n19635),
            .carryout(n19636),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i3_LC_15_14_3.C_ON=1'b1;
    defparam data_idxvec_i3_LC_15_14_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i3_LC_15_14_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i3_LC_15_14_3 (
            .in0(N__47097),
            .in1(N__56934),
            .in2(N__50882),
            .in3(N__37530),
            .lcout(data_idxvec_3),
            .ltout(),
            .carryin(n19636),
            .carryout(n19637),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i4_LC_15_14_4.C_ON=1'b1;
    defparam data_idxvec_i4_LC_15_14_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i4_LC_15_14_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i4_LC_15_14_4 (
            .in0(N__37527),
            .in1(N__56931),
            .in2(N__46217),
            .in3(N__37500),
            .lcout(data_idxvec_4),
            .ltout(),
            .carryin(n19637),
            .carryout(n19638),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i5_LC_15_14_5.C_ON=1'b1;
    defparam data_idxvec_i5_LC_15_14_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i5_LC_15_14_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i5_LC_15_14_5 (
            .in0(N__37486),
            .in1(N__56935),
            .in2(N__51176),
            .in3(N__37470),
            .lcout(data_idxvec_5),
            .ltout(),
            .carryin(n19638),
            .carryout(n19639),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i6_LC_15_14_6.C_ON=1'b1;
    defparam data_idxvec_i6_LC_15_14_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i6_LC_15_14_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i6_LC_15_14_6 (
            .in0(N__47828),
            .in1(N__56932),
            .in2(N__46535),
            .in3(N__37881),
            .lcout(data_idxvec_6),
            .ltout(),
            .carryin(n19639),
            .carryout(n19640),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i7_LC_15_14_7.C_ON=1'b1;
    defparam data_idxvec_i7_LC_15_14_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i7_LC_15_14_7.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i7_LC_15_14_7 (
            .in0(N__37877),
            .in1(N__56936),
            .in2(N__50477),
            .in3(N__37854),
            .lcout(data_idxvec_7),
            .ltout(),
            .carryin(n19640),
            .carryout(n19641),
            .clk(N__54361),
            .ce(N__37986),
            .sr(_gnd_net_));
    defparam data_idxvec_i8_LC_15_15_0.C_ON=1'b1;
    defparam data_idxvec_i8_LC_15_15_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i8_LC_15_15_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i8_LC_15_15_0 (
            .in0(N__37847),
            .in1(N__57021),
            .in2(N__41069),
            .in3(N__37830),
            .lcout(data_idxvec_8),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(n19642),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_idxvec_i9_LC_15_15_1.C_ON=1'b1;
    defparam data_idxvec_i9_LC_15_15_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i9_LC_15_15_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i9_LC_15_15_1 (
            .in0(N__37823),
            .in1(N__56945),
            .in2(N__41195),
            .in3(N__37797),
            .lcout(data_idxvec_9),
            .ltout(),
            .carryin(n19642),
            .carryout(n19643),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_idxvec_i10_LC_15_15_2.C_ON=1'b1;
    defparam data_idxvec_i10_LC_15_15_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i10_LC_15_15_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i10_LC_15_15_2 (
            .in0(N__37794),
            .in1(N__57022),
            .in2(N__41244),
            .in3(N__37776),
            .lcout(data_idxvec_10),
            .ltout(),
            .carryin(n19643),
            .carryout(n19644),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_idxvec_i11_LC_15_15_3.C_ON=1'b1;
    defparam data_idxvec_i11_LC_15_15_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i11_LC_15_15_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i11_LC_15_15_3 (
            .in0(N__44426),
            .in1(N__56946),
            .in2(N__40953),
            .in3(N__37773),
            .lcout(data_idxvec_11),
            .ltout(),
            .carryin(n19644),
            .carryout(n19645),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_idxvec_i12_LC_15_15_4.C_ON=1'b1;
    defparam data_idxvec_i12_LC_15_15_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i12_LC_15_15_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i12_LC_15_15_4 (
            .in0(N__37770),
            .in1(N__57023),
            .in2(N__37749),
            .in3(N__37731),
            .lcout(data_idxvec_12),
            .ltout(),
            .carryin(n19645),
            .carryout(n19646),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_idxvec_i13_LC_15_15_5.C_ON=1'b1;
    defparam data_idxvec_i13_LC_15_15_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i13_LC_15_15_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i13_LC_15_15_5 (
            .in0(N__37727),
            .in1(N__56947),
            .in2(N__37694),
            .in3(N__37674),
            .lcout(data_idxvec_13),
            .ltout(),
            .carryin(n19646),
            .carryout(n19647),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_idxvec_i14_LC_15_15_6.C_ON=1'b1;
    defparam data_idxvec_i14_LC_15_15_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i14_LC_15_15_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i14_LC_15_15_6 (
            .in0(N__38069),
            .in1(N__57024),
            .in2(N__38049),
            .in3(N__38031),
            .lcout(data_idxvec_14),
            .ltout(),
            .carryin(n19647),
            .carryout(n19648),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_idxvec_i15_LC_15_15_7.C_ON=1'b0;
    defparam data_idxvec_i15_LC_15_15_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i15_LC_15_15_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i15_LC_15_15_7 (
            .in0(N__38018),
            .in1(N__38000),
            .in2(N__57095),
            .in3(N__38007),
            .lcout(data_idxvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54374),
            .ce(N__37982),
            .sr(_gnd_net_));
    defparam data_cntvec_i0_i0_LC_15_16_0.C_ON=1'b1;
    defparam data_cntvec_i0_i0_LC_15_16_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i0_LC_15_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i0_LC_15_16_0 (
            .in0(_gnd_net_),
            .in1(N__43387),
            .in2(N__37962),
            .in3(_gnd_net_),
            .lcout(data_cntvec_0),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(n19595),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i1_LC_15_16_1.C_ON=1'b1;
    defparam data_cntvec_i0_i1_LC_15_16_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i1_LC_15_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i1_LC_15_16_1 (
            .in0(_gnd_net_),
            .in1(N__37919),
            .in2(_gnd_net_),
            .in3(N__37899),
            .lcout(data_cntvec_1),
            .ltout(),
            .carryin(n19595),
            .carryout(n19596),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i2_LC_15_16_2.C_ON=1'b1;
    defparam data_cntvec_i0_i2_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i2_LC_15_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i2_LC_15_16_2 (
            .in0(_gnd_net_),
            .in1(N__47123),
            .in2(_gnd_net_),
            .in3(N__37896),
            .lcout(data_cntvec_2),
            .ltout(),
            .carryin(n19596),
            .carryout(n19597),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i3_LC_15_16_3.C_ON=1'b1;
    defparam data_cntvec_i0_i3_LC_15_16_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i3_LC_15_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i3_LC_15_16_3 (
            .in0(_gnd_net_),
            .in1(N__50854),
            .in2(_gnd_net_),
            .in3(N__37893),
            .lcout(data_cntvec_3),
            .ltout(),
            .carryin(n19597),
            .carryout(n19598),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i4_LC_15_16_4.C_ON=1'b1;
    defparam data_cntvec_i0_i4_LC_15_16_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i4_LC_15_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i4_LC_15_16_4 (
            .in0(_gnd_net_),
            .in1(N__46193),
            .in2(_gnd_net_),
            .in3(N__37890),
            .lcout(data_cntvec_4),
            .ltout(),
            .carryin(n19598),
            .carryout(n19599),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i5_LC_15_16_5.C_ON=1'b1;
    defparam data_cntvec_i0_i5_LC_15_16_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i5_LC_15_16_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i5_LC_15_16_5 (
            .in0(_gnd_net_),
            .in1(N__51151),
            .in2(_gnd_net_),
            .in3(N__37887),
            .lcout(data_cntvec_5),
            .ltout(),
            .carryin(n19599),
            .carryout(n19600),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i6_LC_15_16_6.C_ON=1'b1;
    defparam data_cntvec_i0_i6_LC_15_16_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i6_LC_15_16_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i6_LC_15_16_6 (
            .in0(_gnd_net_),
            .in1(N__46507),
            .in2(_gnd_net_),
            .in3(N__37884),
            .lcout(data_cntvec_6),
            .ltout(),
            .carryin(n19600),
            .carryout(n19601),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i7_LC_15_16_7.C_ON=1'b1;
    defparam data_cntvec_i0_i7_LC_15_16_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i7_LC_15_16_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i7_LC_15_16_7 (
            .in0(_gnd_net_),
            .in1(N__50453),
            .in2(_gnd_net_),
            .in3(N__38163),
            .lcout(data_cntvec_7),
            .ltout(),
            .carryin(n19601),
            .carryout(n19602),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38559),
            .sr(N__38481));
    defparam data_cntvec_i0_i8_LC_15_17_0.C_ON=1'b1;
    defparam data_cntvec_i0_i8_LC_15_17_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i8_LC_15_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i8_LC_15_17_0 (
            .in0(_gnd_net_),
            .in1(N__41045),
            .in2(_gnd_net_),
            .in3(N__38160),
            .lcout(data_cntvec_8),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(n19603),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam data_cntvec_i0_i9_LC_15_17_1.C_ON=1'b1;
    defparam data_cntvec_i0_i9_LC_15_17_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i9_LC_15_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i9_LC_15_17_1 (
            .in0(_gnd_net_),
            .in1(N__41171),
            .in2(_gnd_net_),
            .in3(N__38157),
            .lcout(data_cntvec_9),
            .ltout(),
            .carryin(n19603),
            .carryout(n19604),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam data_cntvec_i0_i10_LC_15_17_2.C_ON=1'b1;
    defparam data_cntvec_i0_i10_LC_15_17_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i10_LC_15_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i10_LC_15_17_2 (
            .in0(_gnd_net_),
            .in1(N__41225),
            .in2(_gnd_net_),
            .in3(N__38154),
            .lcout(data_cntvec_10),
            .ltout(),
            .carryin(n19604),
            .carryout(n19605),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam data_cntvec_i0_i11_LC_15_17_3.C_ON=1'b1;
    defparam data_cntvec_i0_i11_LC_15_17_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i11_LC_15_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i11_LC_15_17_3 (
            .in0(_gnd_net_),
            .in1(N__40937),
            .in2(_gnd_net_),
            .in3(N__38151),
            .lcout(data_cntvec_11),
            .ltout(),
            .carryin(n19605),
            .carryout(n19606),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam data_cntvec_i0_i12_LC_15_17_4.C_ON=1'b1;
    defparam data_cntvec_i0_i12_LC_15_17_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i12_LC_15_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i12_LC_15_17_4 (
            .in0(_gnd_net_),
            .in1(N__38144),
            .in2(_gnd_net_),
            .in3(N__38130),
            .lcout(data_cntvec_12),
            .ltout(),
            .carryin(n19606),
            .carryout(n19607),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam data_cntvec_i0_i13_LC_15_17_5.C_ON=1'b1;
    defparam data_cntvec_i0_i13_LC_15_17_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i13_LC_15_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i13_LC_15_17_5 (
            .in0(_gnd_net_),
            .in1(N__38123),
            .in2(_gnd_net_),
            .in3(N__38109),
            .lcout(data_cntvec_13),
            .ltout(),
            .carryin(n19607),
            .carryout(n19608),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam data_cntvec_i0_i14_LC_15_17_6.C_ON=1'b1;
    defparam data_cntvec_i0_i14_LC_15_17_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i14_LC_15_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i14_LC_15_17_6 (
            .in0(_gnd_net_),
            .in1(N__38106),
            .in2(_gnd_net_),
            .in3(N__38094),
            .lcout(data_cntvec_14),
            .ltout(),
            .carryin(n19608),
            .carryout(n19609),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam data_cntvec_i0_i15_LC_15_17_7.C_ON=1'b0;
    defparam data_cntvec_i0_i15_LC_15_17_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i15_LC_15_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i15_LC_15_17_7 (
            .in0(_gnd_net_),
            .in1(N__38084),
            .in2(_gnd_net_),
            .in3(N__38091),
            .lcout(data_cntvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38557),
            .sr(N__38489));
    defparam i6389_3_lut_LC_15_18_0.C_ON=1'b0;
    defparam i6389_3_lut_LC_15_18_0.SEQ_MODE=4'b0000;
    defparam i6389_3_lut_LC_15_18_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i6389_3_lut_LC_15_18_0 (
            .in0(N__41978),
            .in1(N__50302),
            .in2(_gnd_net_),
            .in3(N__47681),
            .lcout(n8_adj_1563),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_171_LC_15_18_1.C_ON=1'b0;
    defparam i1_4_lut_adj_171_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_171_LC_15_18_1.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_171_LC_15_18_1 (
            .in0(N__38450),
            .in1(N__41350),
            .in2(N__38433),
            .in3(N__43357),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6399_3_lut_LC_15_18_2.C_ON=1'b0;
    defparam i6399_3_lut_LC_15_18_2.SEQ_MODE=4'b0000;
    defparam i6399_3_lut_LC_15_18_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6399_3_lut_LC_15_18_2 (
            .in0(N__47895),
            .in1(N__38394),
            .in2(_gnd_net_),
            .in3(N__47682),
            .lcout(n8_adj_1565),
            .ltout(n8_adj_1565_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i6_LC_15_18_3.C_ON=1'b0;
    defparam data_index_i6_LC_15_18_3.SEQ_MODE=4'b1000;
    defparam data_index_i6_LC_15_18_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 data_index_i6_LC_15_18_3 (
            .in0(N__56169),
            .in1(N__56924),
            .in2(N__38397),
            .in3(N__38268),
            .lcout(data_index_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54415),
            .ce(),
            .sr(_gnd_net_));
    defparam i15090_3_lut_LC_15_18_4.C_ON=1'b0;
    defparam i15090_3_lut_LC_15_18_4.SEQ_MODE=4'b0000;
    defparam i15090_3_lut_LC_15_18_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i15090_3_lut_LC_15_18_4 (
            .in0(N__51435),
            .in1(N__40568),
            .in2(_gnd_net_),
            .in3(N__47680),
            .lcout(n17489),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_188_i9_2_lut_3_lut_LC_15_18_5.C_ON=1'b0;
    defparam equal_188_i9_2_lut_3_lut_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam equal_188_i9_2_lut_3_lut_LC_15_18_5.LUT_INIT=16'b1111111111011101;
    LogicCell40 equal_188_i9_2_lut_3_lut_LC_15_18_5 (
            .in0(N__55176),
            .in1(N__57781),
            .in2(_gnd_net_),
            .in3(N__53723),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_15_18_6.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_15_18_6.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_15_18_6.LUT_INIT=16'b0111001001010000;
    LogicCell40 comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_15_18_6 (
            .in0(N__56923),
            .in1(N__56168),
            .in2(N__41123),
            .in3(N__41135),
            .lcout(data_index_9_N_216_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_15_19_2.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_15_19_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_15_19_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_15_19_2 (
            .in0(N__56925),
            .in1(N__56420),
            .in2(N__38280),
            .in3(N__38267),
            .lcout(data_index_9_N_216_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6369_3_lut_LC_15_19_3.C_ON=1'b0;
    defparam i6369_3_lut_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam i6369_3_lut_LC_15_19_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i6369_3_lut_LC_15_19_3 (
            .in0(N__39078),
            .in1(N__40122),
            .in2(_gnd_net_),
            .in3(N__47703),
            .lcout(n8_adj_1559),
            .ltout(n8_adj_1559_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_4 (
            .in0(N__56419),
            .in1(N__39053),
            .in2(N__39042),
            .in3(N__56928),
            .lcout(data_index_9_N_216_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_15_19_5.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_15_19_5.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_15_19_5.LUT_INIT=16'b0100111001000100;
    LogicCell40 comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_15_19_5 (
            .in0(N__56927),
            .in1(N__38951),
            .in2(N__56517),
            .in3(N__42035),
            .lcout(data_index_9_N_216_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_15_19_7.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_15_19_7.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_15_19_7.LUT_INIT=16'b0011101100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_15_19_7 (
            .in0(N__42023),
            .in1(N__56926),
            .in2(N__56516),
            .in3(N__42002),
            .lcout(data_index_9_N_216_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_16MHz_I_0_3_lut_LC_15_20_1.C_ON=1'b0;
    defparam clk_16MHz_I_0_3_lut_LC_15_20_1.SEQ_MODE=4'b0000;
    defparam clk_16MHz_I_0_3_lut_LC_15_20_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 clk_16MHz_I_0_3_lut_LC_15_20_1 (
            .in0(N__38766),
            .in1(N__38703),
            .in2(_gnd_net_),
            .in3(N__38679),
            .lcout(DDS_MCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i1_12200_12201_reset_LC_16_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12200_12201_reset_LC_16_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i1_12200_12201_reset_LC_16_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12200_12201_reset_LC_16_3_0  (
            .in0(N__38607),
            .in1(N__41790),
            .in2(_gnd_net_),
            .in3(N__38591),
            .lcout(\comm_spi.n14619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52626),
            .ce(),
            .sr(N__39363));
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_16_4_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_16_4_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_16_4_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \comm_spi.RESET_I_0_98_2_lut_LC_16_4_0  (
            .in0(N__39605),
            .in1(_gnd_net_),
            .in2(N__55872),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19465_4_lut_3_lut_LC_16_4_1 .C_ON=1'b0;
    defparam \comm_spi.i19465_4_lut_3_lut_LC_16_4_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19465_4_lut_3_lut_LC_16_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19465_4_lut_3_lut_LC_16_4_1  (
            .in0(N__38606),
            .in1(N__42494),
            .in2(_gnd_net_),
            .in3(N__55858),
            .lcout(\comm_spi.n22884 ),
            .ltout(\comm_spi.n22884_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i1_12200_12201_set_LC_16_4_2 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12200_12201_set_LC_16_4_2 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i1_12200_12201_set_LC_16_4_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.data_tx_i1_12200_12201_set_LC_16_4_2  (
            .in0(N__41789),
            .in1(_gnd_net_),
            .in2(N__38595),
            .in3(N__38592),
            .lcout(\comm_spi.n14618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52640),
            .ce(),
            .sr(N__39375));
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_16_4_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_16_4_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_16_4_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_106_2_lut_LC_16_4_3  (
            .in0(_gnd_net_),
            .in1(N__39604),
            .in2(_gnd_net_),
            .in3(N__55849),
            .lcout(\comm_spi.data_tx_7__N_792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19430_4_lut_3_lut_LC_16_4_4 .C_ON=1'b0;
    defparam \comm_spi.i19430_4_lut_3_lut_LC_16_4_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19430_4_lut_3_lut_LC_16_4_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.i19430_4_lut_3_lut_LC_16_4_4  (
            .in0(N__39606),
            .in1(_gnd_net_),
            .in2(N__55873),
            .in3(N__39337),
            .lcout(\comm_spi.n22881 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_16_4_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_16_4_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_16_4_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_105_2_lut_LC_16_4_5  (
            .in0(N__39658),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55848),
            .lcout(\comm_spi.data_tx_7__N_789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_16_4_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_16_4_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_16_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_97_2_lut_LC_16_4_6  (
            .in0(N__55850),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39659),
            .lcout(\comm_spi.data_tx_7__N_771 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19440_4_lut_3_lut_LC_16_4_7 .C_ON=1'b0;
    defparam \comm_spi.i19440_4_lut_3_lut_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19440_4_lut_3_lut_LC_16_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19440_4_lut_3_lut_LC_16_4_7  (
            .in0(N__39660),
            .in1(N__39275),
            .in2(_gnd_net_),
            .in3(N__55857),
            .lcout(\comm_spi.n22878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam wdtick_cnt_3763_3764__i1_LC_16_5_0.C_ON=1'b0;
    defparam wdtick_cnt_3763_3764__i1_LC_16_5_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i1_LC_16_5_0.LUT_INIT=16'b0011001100010001;
    LogicCell40 wdtick_cnt_3763_3764__i1_LC_16_5_0 (
            .in0(N__39259),
            .in1(N__39241),
            .in2(_gnd_net_),
            .in3(N__39222),
            .lcout(wdtick_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39206),
            .ce(N__39447),
            .sr(N__39413));
    defparam wdtick_cnt_3763_3764__i3_LC_16_5_1.C_ON=1'b0;
    defparam wdtick_cnt_3763_3764__i3_LC_16_5_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i3_LC_16_5_1.LUT_INIT=16'b0101101010100000;
    LogicCell40 wdtick_cnt_3763_3764__i3_LC_16_5_1 (
            .in0(N__39224),
            .in1(_gnd_net_),
            .in2(N__39246),
            .in3(N__39260),
            .lcout(wdtick_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39206),
            .ce(N__39447),
            .sr(N__39413));
    defparam wdtick_cnt_3763_3764__i2_LC_16_5_2.C_ON=1'b0;
    defparam wdtick_cnt_3763_3764__i2_LC_16_5_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i2_LC_16_5_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 wdtick_cnt_3763_3764__i2_LC_16_5_2 (
            .in0(_gnd_net_),
            .in1(N__39240),
            .in2(_gnd_net_),
            .in3(N__39223),
            .lcout(wdtick_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39206),
            .ce(N__39447),
            .sr(N__39413));
    defparam \comm_spi.data_tx_i4_12212_12213_set_LC_16_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12212_12213_set_LC_16_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i4_12212_12213_set_LC_16_6_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.data_tx_i4_12212_12213_set_LC_16_6_0  (
            .in0(N__39147),
            .in1(N__39135),
            .in2(_gnd_net_),
            .in3(N__39102),
            .lcout(\comm_spi.n14630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52610),
            .ce(),
            .sr(N__39462));
    defparam i46_2_lut_LC_16_6_2.C_ON=1'b0;
    defparam i46_2_lut_LC_16_6_2.SEQ_MODE=4'b0000;
    defparam i46_2_lut_LC_16_6_2.LUT_INIT=16'b0101010110101010;
    LogicCell40 i46_2_lut_LC_16_6_2 (
            .in0(N__50013),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51720),
            .lcout(n23_adj_1620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9325_1_lut_LC_16_6_4.C_ON=1'b0;
    defparam i9325_1_lut_LC_16_6_4.SEQ_MODE=4'b0000;
    defparam i9325_1_lut_LC_16_6_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i9325_1_lut_LC_16_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44632),
            .lcout(n11741),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_244_LC_16_7_0.C_ON=1'b0;
    defparam i1_4_lut_adj_244_LC_16_7_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_244_LC_16_7_0.LUT_INIT=16'b1010101100000000;
    LogicCell40 i1_4_lut_adj_244_LC_16_7_0 (
            .in0(N__56956),
            .in1(N__39438),
            .in2(N__55512),
            .in3(N__49590),
            .lcout(n11390),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18382_2_lut_LC_16_7_1.C_ON=1'b0;
    defparam i18382_2_lut_LC_16_7_1.SEQ_MODE=4'b0000;
    defparam i18382_2_lut_LC_16_7_1.LUT_INIT=16'b1010000010100000;
    LogicCell40 i18382_2_lut_LC_16_7_1 (
            .in0(N__49487),
            .in1(_gnd_net_),
            .in2(N__51859),
            .in3(_gnd_net_),
            .lcout(n20992),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6834_2_lut_LC_16_7_2.C_ON=1'b0;
    defparam i6834_2_lut_LC_16_7_2.SEQ_MODE=4'b0000;
    defparam i6834_2_lut_LC_16_7_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i6834_2_lut_LC_16_7_2 (
            .in0(_gnd_net_),
            .in1(N__51714),
            .in2(_gnd_net_),
            .in3(N__49486),
            .lcout(n9255),
            .ltout(n9255_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_259_LC_16_7_3.C_ON=1'b0;
    defparam i1_4_lut_adj_259_LC_16_7_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_259_LC_16_7_3.LUT_INIT=16'b1010101000100000;
    LogicCell40 i1_4_lut_adj_259_LC_16_7_3 (
            .in0(N__49589),
            .in1(N__55447),
            .in2(N__39432),
            .in3(N__56957),
            .lcout(n14737),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam flagcntwd_303_LC_16_7_4.C_ON=1'b0;
    defparam flagcntwd_303_LC_16_7_4.SEQ_MODE=4'b1000;
    defparam flagcntwd_303_LC_16_7_4.LUT_INIT=16'b1100110011111111;
    LogicCell40 flagcntwd_303_LC_16_7_4 (
            .in0(_gnd_net_),
            .in1(N__51719),
            .in2(_gnd_net_),
            .in3(N__49488),
            .lcout(flagcntwd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54291),
            .ce(N__39390),
            .sr(N__39569));
    defparam i1_4_lut_adj_279_LC_16_7_5.C_ON=1'b0;
    defparam i1_4_lut_adj_279_LC_16_7_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_279_LC_16_7_5.LUT_INIT=16'b1010100010001000;
    LogicCell40 i1_4_lut_adj_279_LC_16_7_5 (
            .in0(N__49588),
            .in1(N__56953),
            .in2(N__55510),
            .in3(N__49619),
            .lcout(n12336),
            .ltout(n12336_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12386_3_lut_LC_16_7_6.C_ON=1'b0;
    defparam i12386_3_lut_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam i12386_3_lut_LC_16_7_6.LUT_INIT=16'b1010000011110000;
    LogicCell40 i12386_3_lut_LC_16_7_6 (
            .in0(N__56954),
            .in1(_gnd_net_),
            .in2(N__39378),
            .in3(N__52265),
            .lcout(n14799),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_63_LC_16_7_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_63_LC_16_7_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_63_LC_16_7_7.LUT_INIT=16'b1111101000000000;
    LogicCell40 i1_2_lut_3_lut_adj_63_LC_16_7_7 (
            .in0(N__51718),
            .in1(_gnd_net_),
            .in2(N__55511),
            .in3(N__56955),
            .lcout(n20378),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_4_i1_3_lut_LC_16_8_0.C_ON=1'b0;
    defparam mux_137_Mux_4_i1_3_lut_LC_16_8_0.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_4_i1_3_lut_LC_16_8_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_137_Mux_4_i1_3_lut_LC_16_8_0 (
            .in0(N__50732),
            .in1(N__41484),
            .in2(_gnd_net_),
            .in3(N__47783),
            .lcout(n1_adj_1591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_4_i2_3_lut_LC_16_8_1.C_ON=1'b0;
    defparam mux_137_Mux_4_i2_3_lut_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_4_i2_3_lut_LC_16_8_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_4_i2_3_lut_LC_16_8_1 (
            .in0(N__45531),
            .in1(N__39546),
            .in2(_gnd_net_),
            .in3(N__50731),
            .lcout(n2_adj_1592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19294_2_lut_LC_16_8_2.C_ON=1'b0;
    defparam i19294_2_lut_LC_16_8_2.SEQ_MODE=4'b0000;
    defparam i19294_2_lut_LC_16_8_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 i19294_2_lut_LC_16_8_2 (
            .in0(N__50730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39537),
            .lcout(),
            .ltout(n21538_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_LC_16_8_3.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_LC_16_8_3.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_LC_16_8_3.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_1__bdd_4_lut_LC_16_8_3 (
            .in0(N__39498),
            .in1(N__50571),
            .in2(N__39516),
            .in3(N__52386),
            .lcout(),
            .ltout(n22369_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i4_LC_16_8_4.C_ON=1'b0;
    defparam comm_tx_buf_i4_LC_16_8_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i4_LC_16_8_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 comm_tx_buf_i4_LC_16_8_4 (
            .in0(N__50572),
            .in1(N__39513),
            .in2(N__39507),
            .in3(N__39504),
            .lcout(comm_tx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54297),
            .ce(N__45243),
            .sr(N__45164));
    defparam mux_137_Mux_4_i4_3_lut_LC_16_8_5.C_ON=1'b0;
    defparam mux_137_Mux_4_i4_3_lut_LC_16_8_5.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_4_i4_3_lut_LC_16_8_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_4_i4_3_lut_LC_16_8_5 (
            .in0(N__39885),
            .in1(N__42603),
            .in2(_gnd_net_),
            .in3(N__50729),
            .lcout(n4_adj_1593),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_16_8_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_16_8_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.RESET_I_0_103_2_lut_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__55843),
            .in2(_gnd_net_),
            .in3(N__39475),
            .lcout(\comm_spi.data_tx_7__N_783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_16_8_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_16_8_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \comm_spi.RESET_I_0_95_2_lut_LC_16_8_7  (
            .in0(N__39476),
            .in1(_gnd_net_),
            .in2(N__55871),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_LC_16_9_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_LC_16_9_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_LC_16_9_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_0__bdd_4_lut_LC_16_9_0 (
            .in0(N__39708),
            .in1(N__50754),
            .in2(N__45408),
            .in3(N__52404),
            .lcout(),
            .ltout(n22393_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22393_bdd_4_lut_LC_16_9_1.C_ON=1'b0;
    defparam n22393_bdd_4_lut_LC_16_9_1.SEQ_MODE=4'b0000;
    defparam n22393_bdd_4_lut_LC_16_9_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22393_bdd_4_lut_LC_16_9_1 (
            .in0(N__52405),
            .in1(N__44759),
            .in2(N__39696),
            .in3(N__48080),
            .lcout(n22396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_2_i4_3_lut_LC_16_9_2.C_ON=1'b0;
    defparam mux_137_Mux_2_i4_3_lut_LC_16_9_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_2_i4_3_lut_LC_16_9_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_2_i4_3_lut_LC_16_9_2 (
            .in0(N__39834),
            .in1(N__42546),
            .in2(_gnd_net_),
            .in3(N__50756),
            .lcout(),
            .ltout(n4_adj_1595_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18586_4_lut_LC_16_9_3.C_ON=1'b0;
    defparam i18586_4_lut_LC_16_9_3.SEQ_MODE=4'b0000;
    defparam i18586_4_lut_LC_16_9_3.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18586_4_lut_LC_16_9_3 (
            .in0(N__52406),
            .in1(N__39693),
            .in2(N__39672),
            .in3(N__50779),
            .lcout(),
            .ltout(n21196_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i2_LC_16_9_4.C_ON=1'b0;
    defparam comm_tx_buf_i2_LC_16_9_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i2_LC_16_9_4.LUT_INIT=16'b1110010011100100;
    LogicCell40 comm_tx_buf_i2_LC_16_9_4 (
            .in0(N__50598),
            .in1(N__39669),
            .in2(N__39663),
            .in3(_gnd_net_),
            .lcout(comm_tx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54309),
            .ce(N__45226),
            .sr(N__45157));
    defparam mux_137_Mux_1_i4_3_lut_LC_16_9_5.C_ON=1'b0;
    defparam mux_137_Mux_1_i4_3_lut_LC_16_9_5.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_1_i4_3_lut_LC_16_9_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_137_Mux_1_i4_3_lut_LC_16_9_5 (
            .in0(N__50755),
            .in1(N__39813),
            .in2(_gnd_net_),
            .in3(N__43194),
            .lcout(),
            .ltout(n4_adj_1596_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18442_4_lut_LC_16_9_6.C_ON=1'b0;
    defparam i18442_4_lut_LC_16_9_6.SEQ_MODE=4'b0000;
    defparam i18442_4_lut_LC_16_9_6.LUT_INIT=16'b0010001011110000;
    LogicCell40 i18442_4_lut_LC_16_9_6 (
            .in0(N__39642),
            .in1(N__50757),
            .in2(N__39624),
            .in3(N__52407),
            .lcout(),
            .ltout(n21052_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i1_LC_16_9_7.C_ON=1'b0;
    defparam comm_tx_buf_i1_LC_16_9_7.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i1_LC_16_9_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 comm_tx_buf_i1_LC_16_9_7 (
            .in0(_gnd_net_),
            .in1(N__39621),
            .in2(N__39609),
            .in3(N__50597),
            .lcout(comm_tx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54309),
            .ce(N__45226),
            .sr(N__45157));
    defparam comm_buf_5__i0_LC_16_10_0.C_ON=1'b0;
    defparam comm_buf_5__i0_LC_16_10_0.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i0_LC_16_10_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_5__i0_LC_16_10_0 (
            .in0(N__39588),
            .in1(N__51653),
            .in2(_gnd_net_),
            .in3(N__53037),
            .lcout(comm_buf_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_buf_5__i7_LC_16_10_1.C_ON=1'b0;
    defparam comm_buf_5__i7_LC_16_10_1.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i7_LC_16_10_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_5__i7_LC_16_10_1 (
            .in0(N__51652),
            .in1(_gnd_net_),
            .in2(N__39960),
            .in3(N__50389),
            .lcout(comm_buf_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_buf_5__i6_LC_16_10_2.C_ON=1'b0;
    defparam comm_buf_5__i6_LC_16_10_2.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i6_LC_16_10_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i6_LC_16_10_2 (
            .in0(N__46446),
            .in1(N__39930),
            .in2(_gnd_net_),
            .in3(N__51656),
            .lcout(comm_buf_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_buf_5__i5_LC_16_10_3.C_ON=1'b0;
    defparam comm_buf_5__i5_LC_16_10_3.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i5_LC_16_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i5_LC_16_10_3 (
            .in0(N__51651),
            .in1(N__52111),
            .in2(_gnd_net_),
            .in3(N__39915),
            .lcout(comm_buf_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_buf_5__i4_LC_16_10_4.C_ON=1'b0;
    defparam comm_buf_5__i4_LC_16_10_4.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i4_LC_16_10_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i4_LC_16_10_4 (
            .in0(N__46776),
            .in1(N__39900),
            .in2(_gnd_net_),
            .in3(N__51655),
            .lcout(comm_buf_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_buf_5__i3_LC_16_10_5.C_ON=1'b0;
    defparam comm_buf_5__i3_LC_16_10_5.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i3_LC_16_10_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i3_LC_16_10_5 (
            .in0(N__51650),
            .in1(N__51107),
            .in2(_gnd_net_),
            .in3(N__39876),
            .lcout(comm_buf_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_buf_5__i2_LC_16_10_6.C_ON=1'b0;
    defparam comm_buf_5__i2_LC_16_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i2_LC_16_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i2_LC_16_10_6 (
            .in0(N__47231),
            .in1(N__39849),
            .in2(_gnd_net_),
            .in3(N__51654),
            .lcout(comm_buf_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_buf_5__i1_LC_16_10_7.C_ON=1'b0;
    defparam comm_buf_5__i1_LC_16_10_7.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i1_LC_16_10_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i1_LC_16_10_7 (
            .in0(N__51649),
            .in1(N__45792),
            .in2(_gnd_net_),
            .in3(N__39828),
            .lcout(comm_buf_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54322),
            .ce(N__42858),
            .sr(N__42849));
    defparam comm_cmd_0__bdd_4_lut_19664_LC_16_11_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19664_LC_16_11_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19664_LC_16_11_0.LUT_INIT=16'b1110110000101100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19664_LC_16_11_0 (
            .in0(N__39800),
            .in1(N__57475),
            .in2(N__55211),
            .in3(N__39761),
            .lcout(),
            .ltout(n22237_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22237_bdd_4_lut_LC_16_11_1.C_ON=1'b0;
    defparam n22237_bdd_4_lut_LC_16_11_1.SEQ_MODE=4'b0000;
    defparam n22237_bdd_4_lut_LC_16_11_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22237_bdd_4_lut_LC_16_11_1 (
            .in0(N__55132),
            .in1(N__39738),
            .in2(N__40245),
            .in3(N__40242),
            .lcout(n22240),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18452_4_lut_LC_16_11_3.C_ON=1'b0;
    defparam i18452_4_lut_LC_16_11_3.SEQ_MODE=4'b0000;
    defparam i18452_4_lut_LC_16_11_3.LUT_INIT=16'b1110111111100000;
    LogicCell40 i18452_4_lut_LC_16_11_3 (
            .in0(N__57476),
            .in1(N__40215),
            .in2(N__55210),
            .in3(N__41151),
            .lcout(),
            .ltout(n21062_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_LC_16_11_4.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_LC_16_11_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_LC_16_11_4.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_2__bdd_4_lut_LC_16_11_4 (
            .in0(N__53750),
            .in1(N__40206),
            .in2(N__40191),
            .in3(N__54694),
            .lcout(),
            .ltout(n22447_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22447_bdd_4_lut_LC_16_11_5.C_ON=1'b0;
    defparam n22447_bdd_4_lut_LC_16_11_5.SEQ_MODE=4'b0000;
    defparam n22447_bdd_4_lut_LC_16_11_5.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22447_bdd_4_lut_LC_16_11_5 (
            .in0(N__40188),
            .in1(N__40182),
            .in2(N__40167),
            .in3(N__54693),
            .lcout(),
            .ltout(n22450_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i1_LC_16_11_6.C_ON=1'b0;
    defparam comm_buf_0__i1_LC_16_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i1_LC_16_11_6.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_0__i1_LC_16_11_6 (
            .in0(N__52026),
            .in1(N__45793),
            .in2(N__40164),
            .in3(_gnd_net_),
            .lcout(comm_buf_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54334),
            .ce(N__46164),
            .sr(N__43698));
    defparam i36_4_lut_4_lut_LC_16_11_7.C_ON=1'b0;
    defparam i36_4_lut_4_lut_LC_16_11_7.SEQ_MODE=4'b0000;
    defparam i36_4_lut_4_lut_LC_16_11_7.LUT_INIT=16'b0001100011011100;
    LogicCell40 i36_4_lut_4_lut_LC_16_11_7 (
            .in0(N__57474),
            .in1(N__54692),
            .in2(N__55209),
            .in3(N__53749),
            .lcout(n30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19649_LC_16_12_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19649_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19649_LC_16_12_0.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19649_LC_16_12_0 (
            .in0(N__41829),
            .in1(N__54979),
            .in2(N__40029),
            .in3(N__53667),
            .lcout(),
            .ltout(n22273_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22273_bdd_4_lut_LC_16_12_1.C_ON=1'b0;
    defparam n22273_bdd_4_lut_LC_16_12_1.SEQ_MODE=4'b0000;
    defparam n22273_bdd_4_lut_LC_16_12_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22273_bdd_4_lut_LC_16_12_1 (
            .in0(N__53668),
            .in1(N__40020),
            .in2(N__40008),
            .in3(N__40005),
            .lcout(n22276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22285_bdd_4_lut_LC_16_12_2.C_ON=1'b0;
    defparam n22285_bdd_4_lut_LC_16_12_2.SEQ_MODE=4'b0000;
    defparam n22285_bdd_4_lut_LC_16_12_2.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22285_bdd_4_lut_LC_16_12_2 (
            .in0(N__39993),
            .in1(N__40392),
            .in2(N__39978),
            .in3(N__53669),
            .lcout(),
            .ltout(n22288_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1552555_i1_3_lut_LC_16_12_3.C_ON=1'b0;
    defparam i1552555_i1_3_lut_LC_16_12_3.SEQ_MODE=4'b0000;
    defparam i1552555_i1_3_lut_LC_16_12_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 i1552555_i1_3_lut_LC_16_12_3 (
            .in0(N__54695),
            .in1(_gnd_net_),
            .in2(N__40473),
            .in3(N__40470),
            .lcout(),
            .ltout(n30_adj_1539_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i6_LC_16_12_4.C_ON=1'b0;
    defparam comm_buf_0__i6_LC_16_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i6_LC_16_12_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_0__i6_LC_16_12_4 (
            .in0(_gnd_net_),
            .in1(N__46447),
            .in2(N__40464),
            .in3(N__51872),
            .lcout(comm_buf_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54348),
            .ce(N__46167),
            .sr(N__43700));
    defparam mux_128_Mux_6_i19_3_lut_LC_16_12_5.C_ON=1'b0;
    defparam mux_128_Mux_6_i19_3_lut_LC_16_12_5.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_6_i19_3_lut_LC_16_12_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_6_i19_3_lut_LC_16_12_5 (
            .in0(N__40461),
            .in1(N__40433),
            .in2(_gnd_net_),
            .in3(N__57736),
            .lcout(),
            .ltout(n19_adj_1536_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19659_LC_16_12_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19659_LC_16_12_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19659_LC_16_12_6.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19659_LC_16_12_6 (
            .in0(N__40404),
            .in1(N__54978),
            .in2(N__40395),
            .in3(N__53666),
            .lcout(n22285),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19679_LC_16_13_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19679_LC_16_13_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19679_LC_16_13_0.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19679_LC_16_13_0 (
            .in0(N__57624),
            .in1(N__41387),
            .in2(N__40385),
            .in3(N__55215),
            .lcout(),
            .ltout(n22303_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22303_bdd_4_lut_LC_16_13_1.C_ON=1'b0;
    defparam n22303_bdd_4_lut_LC_16_13_1.SEQ_MODE=4'b0000;
    defparam n22303_bdd_4_lut_LC_16_13_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22303_bdd_4_lut_LC_16_13_1 (
            .in0(N__55216),
            .in1(N__40347),
            .in2(N__40320),
            .in3(N__40316),
            .lcout(n22306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22243_bdd_4_lut_LC_16_13_2.C_ON=1'b0;
    defparam n22243_bdd_4_lut_LC_16_13_2.SEQ_MODE=4'b0000;
    defparam n22243_bdd_4_lut_LC_16_13_2.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22243_bdd_4_lut_LC_16_13_2 (
            .in0(N__40287),
            .in1(N__40251),
            .in2(N__40275),
            .in3(N__53728),
            .lcout(n22246),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19634_LC_16_13_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19634_LC_16_13_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19634_LC_16_13_4.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19634_LC_16_13_4 (
            .in0(N__41805),
            .in1(N__55214),
            .in2(N__40260),
            .in3(N__53727),
            .lcout(n22243),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18482_3_lut_LC_16_13_5.C_ON=1'b0;
    defparam i18482_3_lut_LC_16_13_5.SEQ_MODE=4'b0000;
    defparam i18482_3_lut_LC_16_13_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 i18482_3_lut_LC_16_13_5 (
            .in0(N__53729),
            .in1(N__40545),
            .in2(_gnd_net_),
            .in3(N__40539),
            .lcout(),
            .ltout(n21092_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1551349_i1_3_lut_LC_16_13_6.C_ON=1'b0;
    defparam i1551349_i1_3_lut_LC_16_13_6.SEQ_MODE=4'b0000;
    defparam i1551349_i1_3_lut_LC_16_13_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 i1551349_i1_3_lut_LC_16_13_6 (
            .in0(_gnd_net_),
            .in1(N__40530),
            .in2(N__40524),
            .in3(N__54631),
            .lcout(),
            .ltout(n30_adj_1542_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i4_LC_16_13_7.C_ON=1'b0;
    defparam comm_buf_0__i4_LC_16_13_7.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i4_LC_16_13_7.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_0__i4_LC_16_13_7 (
            .in0(N__51904),
            .in1(N__46787),
            .in2(N__40521),
            .in3(_gnd_net_),
            .lcout(comm_buf_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54362),
            .ce(N__46168),
            .sr(N__43723));
    defparam comm_cmd_1__bdd_4_lut_19719_LC_16_14_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19719_LC_16_14_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19719_LC_16_14_1.LUT_INIT=16'b1110011010100010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19719_LC_16_14_1 (
            .in0(N__55217),
            .in1(N__53763),
            .in2(N__53865),
            .in3(N__41205),
            .lcout(),
            .ltout(n22357_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22357_bdd_4_lut_LC_16_14_2.C_ON=1'b0;
    defparam n22357_bdd_4_lut_LC_16_14_2.SEQ_MODE=4'b0000;
    defparam n22357_bdd_4_lut_LC_16_14_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22357_bdd_4_lut_LC_16_14_2 (
            .in0(N__53764),
            .in1(N__40518),
            .in2(N__40509),
            .in3(N__40791),
            .lcout(),
            .ltout(n22360_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18527_3_lut_LC_16_14_3.C_ON=1'b0;
    defparam i18527_3_lut_LC_16_14_3.SEQ_MODE=4'b0000;
    defparam i18527_3_lut_LC_16_14_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 i18527_3_lut_LC_16_14_3 (
            .in0(N__54691),
            .in1(_gnd_net_),
            .in2(N__40506),
            .in3(N__40479),
            .lcout(),
            .ltout(n21137_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i2_LC_16_14_4.C_ON=1'b0;
    defparam comm_buf_0__i2_LC_16_14_4.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i2_LC_16_14_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_0__i2_LC_16_14_4 (
            .in0(_gnd_net_),
            .in1(N__52032),
            .in2(N__40503),
            .in3(N__47244),
            .lcout(comm_buf_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54375),
            .ce(N__46169),
            .sr(N__43724));
    defparam n22327_bdd_4_lut_LC_16_14_6.C_ON=1'b0;
    defparam n22327_bdd_4_lut_LC_16_14_6.SEQ_MODE=4'b0000;
    defparam n22327_bdd_4_lut_LC_16_14_6.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22327_bdd_4_lut_LC_16_14_6 (
            .in0(N__53762),
            .in1(N__40680),
            .in2(N__40500),
            .in3(N__40488),
            .lcout(n22330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_6_i16_3_lut_LC_16_15_0.C_ON=1'b0;
    defparam mux_129_Mux_6_i16_3_lut_LC_16_15_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i16_3_lut_LC_16_15_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_6_i16_3_lut_LC_16_15_0 (
            .in0(N__40750),
            .in1(N__40729),
            .in2(_gnd_net_),
            .in3(N__57614),
            .lcout(n16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_3_i26_3_lut_LC_16_15_1.C_ON=1'b0;
    defparam mux_128_Mux_3_i26_3_lut_LC_16_15_1.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_3_i26_3_lut_LC_16_15_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_3_i26_3_lut_LC_16_15_1 (
            .in0(N__57615),
            .in1(N__40949),
            .in2(_gnd_net_),
            .in3(N__40938),
            .lcout(),
            .ltout(n26_adj_1544_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18475_4_lut_LC_16_15_2.C_ON=1'b0;
    defparam i18475_4_lut_LC_16_15_2.SEQ_MODE=4'b0000;
    defparam i18475_4_lut_LC_16_15_2.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18475_4_lut_LC_16_15_2 (
            .in0(N__55036),
            .in1(N__40917),
            .in2(N__40902),
            .in3(N__57616),
            .lcout(n21085),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18478_3_lut_LC_16_15_3.C_ON=1'b0;
    defparam i18478_3_lut_LC_16_15_3.SEQ_MODE=4'b0000;
    defparam i18478_3_lut_LC_16_15_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18478_3_lut_LC_16_15_3 (
            .in0(N__57618),
            .in1(N__40899),
            .in2(_gnd_net_),
            .in3(N__40821),
            .lcout(n21088),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18567_3_lut_LC_16_15_4.C_ON=1'b0;
    defparam i18567_3_lut_LC_16_15_4.SEQ_MODE=4'b0000;
    defparam i18567_3_lut_LC_16_15_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 i18567_3_lut_LC_16_15_4 (
            .in0(N__55035),
            .in1(N__41357),
            .in2(_gnd_net_),
            .in3(N__40785),
            .lcout(n21177),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i6_LC_16_15_5.C_ON=1'b0;
    defparam buf_dds1_i6_LC_16_15_5.SEQ_MODE=4'b1000;
    defparam buf_dds1_i6_LC_16_15_5.LUT_INIT=16'b1100000010001000;
    LogicCell40 buf_dds1_i6_LC_16_15_5 (
            .in0(N__40754),
            .in1(N__40668),
            .in2(N__47897),
            .in3(N__44971),
            .lcout(buf_dds1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54389),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i6_LC_16_15_6.C_ON=1'b0;
    defparam buf_dds0_i6_LC_16_15_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i6_LC_16_15_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i6_LC_16_15_6 (
            .in0(N__56450),
            .in1(N__40730),
            .in2(N__47896),
            .in3(N__48027),
            .lcout(buf_dds0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54389),
            .ce(),
            .sr(_gnd_net_));
    defparam i18463_3_lut_LC_16_15_7.C_ON=1'b0;
    defparam i18463_3_lut_LC_16_15_7.SEQ_MODE=4'b0000;
    defparam i18463_3_lut_LC_16_15_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18463_3_lut_LC_16_15_7 (
            .in0(N__57617),
            .in1(N__40715),
            .in2(_gnd_net_),
            .in3(N__44678),
            .lcout(n21073),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i11_LC_16_16_0.C_ON=1'b0;
    defparam buf_dds1_i11_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i11_LC_16_16_0.LUT_INIT=16'b1100100000001000;
    LogicCell40 buf_dds1_i11_LC_16_16_0 (
            .in0(N__43966),
            .in1(N__40666),
            .in2(N__44979),
            .in3(N__44177),
            .lcout(buf_dds1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54401),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i5_LC_16_16_1.C_ON=1'b0;
    defparam data_index_i5_LC_16_16_1.SEQ_MODE=4'b1000;
    defparam data_index_i5_LC_16_16_1.LUT_INIT=16'b0111010100100000;
    LogicCell40 data_index_i5_LC_16_16_1 (
            .in0(N__57124),
            .in1(N__56223),
            .in2(N__56598),
            .in3(N__56030),
            .lcout(data_index_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54401),
            .ce(),
            .sr(_gnd_net_));
    defparam i18540_3_lut_LC_16_16_2.C_ON=1'b0;
    defparam i18540_3_lut_LC_16_16_2.SEQ_MODE=4'b0000;
    defparam i18540_3_lut_LC_16_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 i18540_3_lut_LC_16_16_2 (
            .in0(N__41240),
            .in1(N__57803),
            .in2(_gnd_net_),
            .in3(N__41221),
            .lcout(n21150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18450_3_lut_LC_16_16_3.C_ON=1'b0;
    defparam i18450_3_lut_LC_16_16_3.SEQ_MODE=4'b0000;
    defparam i18450_3_lut_LC_16_16_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 i18450_3_lut_LC_16_16_3 (
            .in0(N__57802),
            .in1(_gnd_net_),
            .in2(N__41196),
            .in3(N__41167),
            .lcout(n21060),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i3_LC_16_16_4.C_ON=1'b0;
    defparam data_index_i3_LC_16_16_4.SEQ_MODE=4'b1000;
    defparam data_index_i3_LC_16_16_4.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i3_LC_16_16_4 (
            .in0(N__41142),
            .in1(N__57125),
            .in2(N__56343),
            .in3(N__41124),
            .lcout(data_index_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54401),
            .ce(),
            .sr(_gnd_net_));
    defparam i18555_3_lut_LC_16_16_6.C_ON=1'b0;
    defparam i18555_3_lut_LC_16_16_6.SEQ_MODE=4'b0000;
    defparam i18555_3_lut_LC_16_16_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 i18555_3_lut_LC_16_16_6 (
            .in0(N__41070),
            .in1(N__57801),
            .in2(_gnd_net_),
            .in3(N__41041),
            .lcout(n21165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18474_4_lut_LC_16_16_7.C_ON=1'b0;
    defparam i18474_4_lut_LC_16_16_7.SEQ_MODE=4'b0000;
    defparam i18474_4_lut_LC_16_16_7.LUT_INIT=16'b0111010000110000;
    LogicCell40 i18474_4_lut_LC_16_16_7 (
            .in0(N__57800),
            .in1(N__55125),
            .in2(N__41904),
            .in3(N__41025),
            .lcout(n21084),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i2_LC_16_17_0.C_ON=1'b0;
    defparam acadc_skipCount_i2_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i2_LC_16_17_0.LUT_INIT=16'b0000110010101010;
    LogicCell40 acadc_skipCount_i2_LC_16_17_0 (
            .in0(N__46579),
            .in1(N__48066),
            .in2(N__56321),
            .in3(N__44316),
            .lcout(acadc_skipCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54416),
            .ce(),
            .sr(_gnd_net_));
    defparam i6439_3_lut_LC_16_17_1.C_ON=1'b0;
    defparam i6439_3_lut_LC_16_17_1.SEQ_MODE=4'b0000;
    defparam i6439_3_lut_LC_16_17_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 i6439_3_lut_LC_16_17_1 (
            .in0(N__47691),
            .in1(N__48059),
            .in2(_gnd_net_),
            .in3(N__40996),
            .lcout(n8_adj_1571),
            .ltout(n8_adj_1571_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i2_LC_16_17_2.C_ON=1'b0;
    defparam data_index_i2_LC_16_17_2.SEQ_MODE=4'b1000;
    defparam data_index_i2_LC_16_17_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 data_index_i2_LC_16_17_2 (
            .in0(N__56202),
            .in1(N__57094),
            .in2(N__41007),
            .in3(N__45093),
            .lcout(data_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54416),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i10_LC_16_17_3.C_ON=1'b0;
    defparam buf_dds0_i10_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i10_LC_16_17_3.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_dds0_i10_LC_16_17_3 (
            .in0(N__40969),
            .in1(N__56203),
            .in2(N__44769),
            .in3(N__48024),
            .lcout(buf_dds0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54416),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_304_LC_16_17_4.C_ON=1'b0;
    defparam i1_4_lut_adj_304_LC_16_17_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_304_LC_16_17_4.LUT_INIT=16'b1100000011000100;
    LogicCell40 i1_4_lut_adj_304_LC_16_17_4 (
            .in0(N__41552),
            .in1(N__57093),
            .in2(N__56320),
            .in3(N__41777),
            .lcout(n12429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6973_2_lut_LC_16_17_5.C_ON=1'b0;
    defparam i6973_2_lut_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam i6973_2_lut_LC_16_17_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i6973_2_lut_LC_16_17_5 (
            .in0(_gnd_net_),
            .in1(N__51959),
            .in2(_gnd_net_),
            .in3(N__55499),
            .lcout(n9306),
            .ltout(n9306_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i13_LC_16_17_6.C_ON=1'b0;
    defparam buf_dds0_i13_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i13_LC_16_17_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_dds0_i13_LC_16_17_6 (
            .in0(N__48025),
            .in1(N__43593),
            .in2(N__41634),
            .in3(N__41617),
            .lcout(buf_dds0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54416),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_165_LC_16_17_7.C_ON=1'b0;
    defparam i6_4_lut_adj_165_LC_16_17_7.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_165_LC_16_17_7.LUT_INIT=16'b0111110110111110;
    LogicCell40 i6_4_lut_adj_165_LC_16_17_7 (
            .in0(N__41601),
            .in1(N__41583),
            .in2(N__46580),
            .in3(N__46972),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_248_LC_16_18_0.C_ON=1'b0;
    defparam i1_4_lut_adj_248_LC_16_18_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_248_LC_16_18_0.LUT_INIT=16'b1100110000000100;
    LogicCell40 i1_4_lut_adj_248_LC_16_18_0 (
            .in0(N__41553),
            .in1(N__57122),
            .in2(N__41541),
            .in3(N__56170),
            .lcout(n12381),
            .ltout(n12381_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i5_LC_16_18_1.C_ON=1'b0;
    defparam buf_device_acadc_i5_LC_16_18_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i5_LC_16_18_1.LUT_INIT=16'b0100111101000000;
    LogicCell40 buf_device_acadc_i5_LC_16_18_1 (
            .in0(N__56175),
            .in1(N__41465),
            .in2(N__41403),
            .in3(N__41377),
            .lcout(VAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54422),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i0_LC_16_18_3.C_ON=1'b0;
    defparam acadc_skipCount_i0_LC_16_18_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i0_LC_16_18_3.LUT_INIT=16'b0011101100001000;
    LogicCell40 acadc_skipCount_i0_LC_16_18_3 (
            .in0(N__43282),
            .in1(N__44329),
            .in2(N__56291),
            .in3(N__43361),
            .lcout(acadc_skipCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54422),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i6_LC_16_18_5.C_ON=1'b0;
    defparam acadc_skipCount_i6_LC_16_18_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i6_LC_16_18_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i6_LC_16_18_5 (
            .in0(N__56174),
            .in1(N__44330),
            .in2(N__47901),
            .in3(N__41358),
            .lcout(acadc_skipCount_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54422),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19329_4_lut_LC_16_18_7 .C_ON=1'b0;
    defparam \SIG_DDS.i19329_4_lut_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19329_4_lut_LC_16_18_7 .LUT_INIT=16'b1100110001000110;
    LogicCell40 \SIG_DDS.i19329_4_lut_LC_16_18_7  (
            .in0(N__41323),
            .in1(N__42267),
            .in2(N__42132),
            .in3(N__43020),
            .lcout(\SIG_DDS.n12722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6379_3_lut_LC_16_19_0.C_ON=1'b0;
    defparam i6379_3_lut_LC_16_19_0.SEQ_MODE=4'b0000;
    defparam i6379_3_lut_LC_16_19_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6379_3_lut_LC_16_19_0 (
            .in0(N__43783),
            .in1(N__42063),
            .in2(_gnd_net_),
            .in3(N__47702),
            .lcout(n8_adj_1561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i7_LC_16_19_2.C_ON=1'b0;
    defparam data_index_i7_LC_16_19_2.SEQ_MODE=4'b1000;
    defparam data_index_i7_LC_16_19_2.LUT_INIT=16'b0101000011011000;
    LogicCell40 data_index_i7_LC_16_19_2 (
            .in0(N__57123),
            .in1(N__42024),
            .in2(N__42012),
            .in3(N__56316),
            .lcout(data_index_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54429),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_3_i23_3_lut_LC_16_19_4.C_ON=1'b0;
    defparam mux_128_Mux_3_i23_3_lut_LC_16_19_4.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_3_i23_3_lut_LC_16_19_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_3_i23_3_lut_LC_16_19_4 (
            .in0(N__41954),
            .in1(N__57758),
            .in2(_gnd_net_),
            .in3(N__41934),
            .lcout(n23_adj_1543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i0_LC_16_19_5.C_ON=1'b0;
    defparam buf_control_i0_LC_16_19_5.SEQ_MODE=4'b1000;
    defparam buf_control_i0_LC_16_19_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i0_LC_16_19_5 (
            .in0(N__56315),
            .in1(N__41892),
            .in2(N__43808),
            .in3(N__44611),
            .lcout(buf_control_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54429),
            .ce(),
            .sr(_gnd_net_));
    defparam i19085_2_lut_LC_17_2_2.C_ON=1'b0;
    defparam i19085_2_lut_LC_17_2_2.SEQ_MODE=4'b0000;
    defparam i19085_2_lut_LC_17_2_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19085_2_lut_LC_17_2_2 (
            .in0(_gnd_net_),
            .in1(N__41838),
            .in2(_gnd_net_),
            .in3(N__57822),
            .lcout(n21273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19092_2_lut_LC_17_3_0.C_ON=1'b0;
    defparam i19092_2_lut_LC_17_3_0.SEQ_MODE=4'b0000;
    defparam i19092_2_lut_LC_17_3_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 i19092_2_lut_LC_17_3_0 (
            .in0(_gnd_net_),
            .in1(N__41817),
            .in2(_gnd_net_),
            .in3(N__57821),
            .lcout(n21569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12174_12175_set_LC_17_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12174_12175_set_LC_17_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i0_12174_12175_set_LC_17_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_12174_12175_set_LC_17_4_0  (
            .in0(N__58293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52602),
            .ce(),
            .sr(N__42465));
    defparam \comm_spi.data_tx_i5_12216_12217_reset_LC_17_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12216_12217_reset_LC_17_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i5_12216_12217_reset_LC_17_5_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_tx_i5_12216_12217_reset_LC_17_5_0  (
            .in0(N__44528),
            .in1(N__44561),
            .in2(_gnd_net_),
            .in3(N__44516),
            .lcout(\comm_spi.n14635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52586),
            .ce(),
            .sr(N__42360));
    defparam \comm_spi.data_tx_i6_12220_12221_reset_LC_17_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12220_12221_reset_LC_17_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i6_12220_12221_reset_LC_17_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_tx_i6_12220_12221_reset_LC_17_6_0  (
            .in0(N__44469),
            .in1(N__44486),
            .in2(_gnd_net_),
            .in3(N__44456),
            .lcout(\comm_spi.n14639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52552),
            .ce(),
            .sr(N__42372));
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_17_7_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_17_7_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_101_2_lut_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__45260),
            .in2(_gnd_net_),
            .in3(N__55757),
            .lcout(\comm_spi.data_tx_7__N_777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_17_7_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_17_7_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_102_2_lut_LC_17_7_5  (
            .in0(_gnd_net_),
            .in1(N__42734),
            .in2(_gnd_net_),
            .in3(N__55758),
            .lcout(\comm_spi.data_tx_7__N_780 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_6_i4_3_lut_LC_17_7_6.C_ON=1'b0;
    defparam mux_137_Mux_6_i4_3_lut_LC_17_7_6.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_6_i4_3_lut_LC_17_7_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_6_i4_3_lut_LC_17_7_6 (
            .in0(N__42348),
            .in1(N__42645),
            .in2(_gnd_net_),
            .in3(N__50790),
            .lcout(n4_adj_1590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19455_4_lut_3_lut_LC_17_7_7 .C_ON=1'b0;
    defparam \comm_spi.i19455_4_lut_3_lut_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19455_4_lut_3_lut_LC_17_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19455_4_lut_3_lut_LC_17_7_7  (
            .in0(N__44485),
            .in1(N__42735),
            .in2(_gnd_net_),
            .in3(N__55759),
            .lcout(\comm_spi.n22869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19580_LC_17_8_0.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19580_LC_17_8_0.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19580_LC_17_8_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_1__bdd_4_lut_19580_LC_17_8_0 (
            .in0(N__42324),
            .in1(N__50599),
            .in2(N__42297),
            .in3(N__52387),
            .lcout(),
            .ltout(n22183_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i0_LC_17_8_1.C_ON=1'b0;
    defparam comm_tx_buf_i0_LC_17_8_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i0_LC_17_8_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 comm_tx_buf_i0_LC_17_8_1 (
            .in0(N__50600),
            .in1(N__42522),
            .in2(N__42339),
            .in3(N__42501),
            .lcout(comm_tx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54310),
            .ce(N__45236),
            .sr(N__45171));
    defparam mux_137_Mux_0_i4_3_lut_LC_17_8_2.C_ON=1'b0;
    defparam mux_137_Mux_0_i4_3_lut_LC_17_8_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_0_i4_3_lut_LC_17_8_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_0_i4_3_lut_LC_17_8_2 (
            .in0(N__42336),
            .in1(N__42699),
            .in2(_gnd_net_),
            .in3(N__50795),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18964_2_lut_LC_17_8_3.C_ON=1'b0;
    defparam i18964_2_lut_LC_17_8_3.SEQ_MODE=4'b0000;
    defparam i18964_2_lut_LC_17_8_3.LUT_INIT=16'b0101010100000000;
    LogicCell40 i18964_2_lut_LC_17_8_3 (
            .in0(N__50794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42318),
            .lcout(n21211),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_0_i1_3_lut_LC_17_8_4.C_ON=1'b0;
    defparam mux_137_Mux_0_i1_3_lut_LC_17_8_4.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_0_i1_3_lut_LC_17_8_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_0_i1_3_lut_LC_17_8_4 (
            .in0(N__43291),
            .in1(N__43825),
            .in2(_gnd_net_),
            .in3(N__50797),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_0_i2_3_lut_LC_17_8_5.C_ON=1'b0;
    defparam mux_137_Mux_0_i2_3_lut_LC_17_8_5.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_0_i2_3_lut_LC_17_8_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_137_Mux_0_i2_3_lut_LC_17_8_5 (
            .in0(N__50796),
            .in1(N__45552),
            .in2(_gnd_net_),
            .in3(N__42513),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_17_8_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_17_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_99_2_lut_LC_17_8_7  (
            .in0(N__42481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55847),
            .lcout(\comm_spi.data_tx_7__N_773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15080_3_lut_LC_17_9_0.C_ON=1'b0;
    defparam i15080_3_lut_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam i15080_3_lut_LC_17_9_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i15080_3_lut_LC_17_9_0 (
            .in0(N__42621),
            .in1(N__43567),
            .in2(_gnd_net_),
            .in3(N__50596),
            .lcout(),
            .ltout(n17479_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i5_LC_17_9_1.C_ON=1'b0;
    defparam comm_tx_buf_i5_LC_17_9_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i5_LC_17_9_1.LUT_INIT=16'b1010101011011000;
    LogicCell40 comm_tx_buf_i5_LC_17_9_1 (
            .in0(N__42393),
            .in1(N__42417),
            .in2(N__42450),
            .in3(N__50778),
            .lcout(comm_tx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54323),
            .ce(N__45235),
            .sr(N__45173));
    defparam i19282_2_lut_LC_17_9_2.C_ON=1'b0;
    defparam i19282_2_lut_LC_17_9_2.SEQ_MODE=4'b0000;
    defparam i19282_2_lut_LC_17_9_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19282_2_lut_LC_17_9_2 (
            .in0(_gnd_net_),
            .in1(N__45450),
            .in2(_gnd_net_),
            .in3(N__50593),
            .lcout(n21212),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15081_3_lut_LC_17_9_3.C_ON=1'b0;
    defparam i15081_3_lut_LC_17_9_3.SEQ_MODE=4'b0000;
    defparam i15081_3_lut_LC_17_9_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i15081_3_lut_LC_17_9_3 (
            .in0(N__50595),
            .in1(N__42447),
            .in2(_gnd_net_),
            .in3(N__42429),
            .lcout(n17480),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15083_3_lut_LC_17_9_4.C_ON=1'b0;
    defparam i15083_3_lut_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam i15083_3_lut_LC_17_9_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 i15083_3_lut_LC_17_9_4 (
            .in0(N__42408),
            .in1(N__51436),
            .in2(_gnd_net_),
            .in3(N__50594),
            .lcout(),
            .ltout(n17482_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19699_LC_17_9_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19699_LC_17_9_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19699_LC_17_9_5.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_index_1__bdd_4_lut_19699_LC_17_9_5 (
            .in0(N__42402),
            .in1(N__50777),
            .in2(N__42396),
            .in3(N__52408),
            .lcout(n22189),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_17_9_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_17_9_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \comm_spi.RESET_I_0_94_2_lut_LC_17_9_7  (
            .in0(N__42728),
            .in1(N__55827),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i0_LC_17_10_0.C_ON=1'b0;
    defparam comm_buf_4__i0_LC_17_10_0.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i0_LC_17_10_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_4__i0_LC_17_10_0 (
            .in0(N__42717),
            .in1(N__52016),
            .in2(_gnd_net_),
            .in3(N__53036),
            .lcout(comm_buf_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam comm_buf_4__i7_LC_17_10_1.C_ON=1'b0;
    defparam comm_buf_4__i7_LC_17_10_1.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i7_LC_17_10_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i7_LC_17_10_1 (
            .in0(N__52015),
            .in1(N__50410),
            .in2(_gnd_net_),
            .in3(N__42690),
            .lcout(comm_buf_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam comm_buf_4__i6_LC_17_10_2.C_ON=1'b0;
    defparam comm_buf_4__i6_LC_17_10_2.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i6_LC_17_10_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_4__i6_LC_17_10_2 (
            .in0(N__42660),
            .in1(N__52017),
            .in2(_gnd_net_),
            .in3(N__46462),
            .lcout(comm_buf_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam comm_buf_4__i5_LC_17_10_3.C_ON=1'b0;
    defparam comm_buf_4__i5_LC_17_10_3.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i5_LC_17_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i5_LC_17_10_3 (
            .in0(N__52014),
            .in1(N__52113),
            .in2(_gnd_net_),
            .in3(N__42636),
            .lcout(comm_buf_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam comm_buf_4__i4_LC_17_10_4.C_ON=1'b0;
    defparam comm_buf_4__i4_LC_17_10_4.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i4_LC_17_10_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i4_LC_17_10_4 (
            .in0(N__46786),
            .in1(N__42615),
            .in2(_gnd_net_),
            .in3(N__52019),
            .lcout(comm_buf_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam comm_buf_4__i3_LC_17_10_5.C_ON=1'b0;
    defparam comm_buf_4__i3_LC_17_10_5.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i3_LC_17_10_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i3_LC_17_10_5 (
            .in0(N__52013),
            .in1(N__51110),
            .in2(_gnd_net_),
            .in3(N__42591),
            .lcout(comm_buf_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam comm_buf_4__i2_LC_17_10_6.C_ON=1'b0;
    defparam comm_buf_4__i2_LC_17_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i2_LC_17_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i2_LC_17_10_6 (
            .in0(N__47232),
            .in1(N__42564),
            .in2(_gnd_net_),
            .in3(N__52018),
            .lcout(comm_buf_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam comm_buf_4__i1_LC_17_10_7.C_ON=1'b0;
    defparam comm_buf_4__i1_LC_17_10_7.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i1_LC_17_10_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i1_LC_17_10_7 (
            .in0(N__52012),
            .in1(N__45787),
            .in2(_gnd_net_),
            .in3(N__42540),
            .lcout(comm_buf_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54335),
            .ce(N__45810),
            .sr(N__42843));
    defparam \SIG_DDS.bit_cnt_i3_LC_17_11_0 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i3_LC_17_11_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i3_LC_17_11_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \SIG_DDS.bit_cnt_i3_LC_17_11_0  (
            .in0(N__43170),
            .in1(N__43091),
            .in2(N__43127),
            .in3(N__43184),
            .lcout(\SIG_DDS.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54349),
            .ce(N__43074),
            .sr(N__42885));
    defparam \SIG_DDS.bit_cnt_i1_LC_17_11_1 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i1_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i1_LC_17_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \SIG_DDS.bit_cnt_i1_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__43116),
            .in2(_gnd_net_),
            .in3(N__43168),
            .lcout(\SIG_DDS.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54349),
            .ce(N__43074),
            .sr(N__42885));
    defparam \SIG_DDS.bit_cnt_i2_LC_17_11_2 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i2_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i2_LC_17_11_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \SIG_DDS.bit_cnt_i2_LC_17_11_2  (
            .in0(N__43169),
            .in1(_gnd_net_),
            .in2(N__43126),
            .in3(N__43090),
            .lcout(\SIG_DDS.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54349),
            .ce(N__43074),
            .sr(N__42885));
    defparam i1_3_lut_adj_277_LC_17_11_3.C_ON=1'b0;
    defparam i1_3_lut_adj_277_LC_17_11_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_277_LC_17_11_3.LUT_INIT=16'b1100110010001000;
    LogicCell40 i1_3_lut_adj_277_LC_17_11_3 (
            .in0(N__45882),
            .in1(N__45916),
            .in2(_gnd_net_),
            .in3(N__46092),
            .lcout(n12220),
            .ltout(n12220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12372_2_lut_LC_17_11_4.C_ON=1'b0;
    defparam i12372_2_lut_LC_17_11_4.SEQ_MODE=4'b0000;
    defparam i12372_2_lut_LC_17_11_4.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12372_2_lut_LC_17_11_4 (
            .in0(N__57069),
            .in1(_gnd_net_),
            .in2(N__42852),
            .in3(_gnd_net_),
            .lcout(n14785),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12337_2_lut_LC_17_11_5.C_ON=1'b0;
    defparam i12337_2_lut_LC_17_11_5.SEQ_MODE=4'b0000;
    defparam i12337_2_lut_LC_17_11_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12337_2_lut_LC_17_11_5 (
            .in0(_gnd_net_),
            .in1(N__57067),
            .in2(_gnd_net_),
            .in3(N__46123),
            .lcout(n14750),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12365_2_lut_LC_17_11_6.C_ON=1'b0;
    defparam i12365_2_lut_LC_17_11_6.SEQ_MODE=4'b0000;
    defparam i12365_2_lut_LC_17_11_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12365_2_lut_LC_17_11_6 (
            .in0(N__57068),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45806),
            .lcout(n14778),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i7_LC_17_12_0.C_ON=1'b0;
    defparam comm_buf_0__i7_LC_17_12_0.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i7_LC_17_12_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_0__i7_LC_17_12_0 (
            .in0(N__52020),
            .in1(N__50411),
            .in2(_gnd_net_),
            .in3(N__42831),
            .lcout(comm_buf_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54363),
            .ce(N__46165),
            .sr(N__43699));
    defparam comm_buf_0__i5_LC_17_12_1.C_ON=1'b0;
    defparam comm_buf_0__i5_LC_17_12_1.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i5_LC_17_12_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_0__i5_LC_17_12_1 (
            .in0(N__52117),
            .in1(N__43623),
            .in2(_gnd_net_),
            .in3(N__52021),
            .lcout(comm_buf_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54363),
            .ce(N__46165),
            .sr(N__43699));
    defparam n22213_bdd_4_lut_LC_17_13_0.C_ON=1'b0;
    defparam n22213_bdd_4_lut_LC_17_13_0.SEQ_MODE=4'b0000;
    defparam n22213_bdd_4_lut_LC_17_13_0.LUT_INIT=16'b1101100111001000;
    LogicCell40 n22213_bdd_4_lut_LC_17_13_0 (
            .in0(N__53755),
            .in1(N__43422),
            .in2(N__43521),
            .in3(N__43482),
            .lcout(n22216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19611_LC_17_13_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19611_LC_17_13_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19611_LC_17_13_1.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19611_LC_17_13_1 (
            .in0(N__43467),
            .in1(N__55151),
            .in2(N__43449),
            .in3(N__53754),
            .lcout(n22213),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_0_i26_3_lut_LC_17_13_2.C_ON=1'b0;
    defparam mux_129_Mux_0_i26_3_lut_LC_17_13_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i26_3_lut_LC_17_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_0_i26_3_lut_LC_17_13_2 (
            .in0(N__43416),
            .in1(N__57626),
            .in2(_gnd_net_),
            .in3(N__43392),
            .lcout(),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19593_LC_17_13_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19593_LC_17_13_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19593_LC_17_13_3.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19593_LC_17_13_3 (
            .in0(N__52695),
            .in1(N__55152),
            .in2(N__43368),
            .in3(N__53756),
            .lcout(),
            .ltout(n22201_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22201_bdd_4_lut_LC_17_13_4.C_ON=1'b0;
    defparam n22201_bdd_4_lut_LC_17_13_4.SEQ_MODE=4'b0000;
    defparam n22201_bdd_4_lut_LC_17_13_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22201_bdd_4_lut_LC_17_13_4 (
            .in0(N__53757),
            .in1(N__43365),
            .in2(N__43341),
            .in3(N__43338),
            .lcout(),
            .ltout(n22204_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1556173_i1_3_lut_LC_17_13_5.C_ON=1'b0;
    defparam i1556173_i1_3_lut_LC_17_13_5.SEQ_MODE=4'b0000;
    defparam i1556173_i1_3_lut_LC_17_13_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1556173_i1_3_lut_LC_17_13_5 (
            .in0(_gnd_net_),
            .in1(N__43311),
            .in2(N__43305),
            .in3(N__54746),
            .lcout(),
            .ltout(n30_adj_1485_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i0_LC_17_13_6.C_ON=1'b0;
    defparam comm_buf_1__i0_LC_17_13_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i0_LC_17_13_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_1__i0_LC_17_13_6 (
            .in0(N__52022),
            .in1(_gnd_net_),
            .in2(N__43302),
            .in3(N__53051),
            .lcout(comm_buf_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54376),
            .ce(N__51381),
            .sr(N__51277));
    defparam comm_cmd_0__bdd_4_lut_19669_LC_17_14_1.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19669_LC_17_14_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19669_LC_17_14_1.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19669_LC_17_14_1 (
            .in0(N__44108),
            .in1(N__55160),
            .in2(N__43229),
            .in3(N__57625),
            .lcout(),
            .ltout(n22297_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22297_bdd_4_lut_LC_17_14_2.C_ON=1'b0;
    defparam n22297_bdd_4_lut_LC_17_14_2.SEQ_MODE=4'b0000;
    defparam n22297_bdd_4_lut_LC_17_14_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22297_bdd_4_lut_LC_17_14_2 (
            .in0(N__55161),
            .in1(N__44001),
            .in2(N__43974),
            .in3(N__43970),
            .lcout(n22300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22309_bdd_4_lut_LC_17_14_5.C_ON=1'b0;
    defparam n22309_bdd_4_lut_LC_17_14_5.SEQ_MODE=4'b0000;
    defparam n22309_bdd_4_lut_LC_17_14_5.LUT_INIT=16'b1110111000110000;
    LogicCell40 n22309_bdd_4_lut_LC_17_14_5 (
            .in0(N__43941),
            .in1(N__54697),
            .in2(N__43932),
            .in3(N__44340),
            .lcout(),
            .ltout(n22312_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i3_LC_17_14_6.C_ON=1'b0;
    defparam comm_buf_0__i3_LC_17_14_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i3_LC_17_14_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_0__i3_LC_17_14_6 (
            .in0(N__51114),
            .in1(_gnd_net_),
            .in2(N__43923),
            .in3(N__51993),
            .lcout(comm_buf_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54390),
            .ce(N__46166),
            .sr(N__43710));
    defparam comm_cmd_0__bdd_4_lut_19616_LC_17_15_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19616_LC_17_15_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19616_LC_17_15_0.LUT_INIT=16'b1110011011000100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19616_LC_17_15_0 (
            .in0(N__55034),
            .in1(N__57604),
            .in2(N__43920),
            .in3(N__43881),
            .lcout(n22219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18461_3_lut_LC_17_15_5.C_ON=1'b0;
    defparam i18461_3_lut_LC_17_15_5.SEQ_MODE=4'b0000;
    defparam i18461_3_lut_LC_17_15_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 i18461_3_lut_LC_17_15_5 (
            .in0(N__43854),
            .in1(_gnd_net_),
            .in2(N__44361),
            .in3(N__54687),
            .lcout(),
            .ltout(n21071_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i0_LC_17_15_6.C_ON=1'b0;
    defparam comm_buf_0__i0_LC_17_15_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i0_LC_17_15_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_0__i0_LC_17_15_6 (
            .in0(_gnd_net_),
            .in1(N__51992),
            .in2(N__43839),
            .in3(N__53055),
            .lcout(comm_buf_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54402),
            .ce(N__46173),
            .sr(N__43725));
    defparam i19115_4_lut_4_lut_LC_17_15_7.C_ON=1'b0;
    defparam i19115_4_lut_4_lut_LC_17_15_7.SEQ_MODE=4'b0000;
    defparam i19115_4_lut_4_lut_LC_17_15_7.LUT_INIT=16'b1110111101101011;
    LogicCell40 i19115_4_lut_4_lut_LC_17_15_7 (
            .in0(N__57603),
            .in1(N__54686),
            .in2(N__55147),
            .in3(N__53672),
            .lcout(n21341),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22219_bdd_4_lut_LC_17_16_0.C_ON=1'b0;
    defparam n22219_bdd_4_lut_LC_17_16_0.SEQ_MODE=4'b0000;
    defparam n22219_bdd_4_lut_LC_17_16_0.LUT_INIT=16'b1011101010011000;
    LogicCell40 n22219_bdd_4_lut_LC_17_16_0 (
            .in0(N__43656),
            .in1(N__55188),
            .in2(N__44616),
            .in3(N__43650),
            .lcout(n22222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15338_2_lut_3_lut_LC_17_16_1.C_ON=1'b0;
    defparam i15338_2_lut_3_lut_LC_17_16_1.SEQ_MODE=4'b0000;
    defparam i15338_2_lut_3_lut_LC_17_16_1.LUT_INIT=16'b0000000000001010;
    LogicCell40 i15338_2_lut_3_lut_LC_17_16_1 (
            .in0(N__44187),
            .in1(_gnd_net_),
            .in2(N__55556),
            .in3(N__51960),
            .lcout(n14_adj_1578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_187_i9_2_lut_3_lut_LC_17_16_2.C_ON=1'b0;
    defparam equal_187_i9_2_lut_3_lut_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam equal_187_i9_2_lut_3_lut_LC_17_16_2.LUT_INIT=16'b1111111110111011;
    LogicCell40 equal_187_i9_2_lut_3_lut_LC_17_16_2 (
            .in0(N__53765),
            .in1(N__57759),
            .in2(_gnd_net_),
            .in3(N__55187),
            .lcout(n9_adj_1415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18557_4_lut_LC_17_16_3.C_ON=1'b0;
    defparam i18557_4_lut_LC_17_16_3.SEQ_MODE=4'b0000;
    defparam i18557_4_lut_LC_17_16_3.LUT_INIT=16'b1111110110101000;
    LogicCell40 i18557_4_lut_LC_17_16_3 (
            .in0(N__55189),
            .in1(N__57804),
            .in2(N__44394),
            .in3(N__44376),
            .lcout(),
            .ltout(n21167_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18460_3_lut_LC_17_16_4.C_ON=1'b0;
    defparam i18460_3_lut_LC_17_16_4.SEQ_MODE=4'b0000;
    defparam i18460_3_lut_LC_17_16_4.LUT_INIT=16'b1111001111000000;
    LogicCell40 i18460_3_lut_LC_17_16_4 (
            .in0(_gnd_net_),
            .in1(N__53761),
            .in2(N__44370),
            .in3(N__44367),
            .lcout(n21070),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19684_LC_17_16_7.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19684_LC_17_16_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19684_LC_17_16_7.LUT_INIT=16'b1111100001011000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19684_LC_17_16_7 (
            .in0(N__54696),
            .in1(N__44352),
            .in2(N__53796),
            .in3(N__44346),
            .lcout(n22309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i3_LC_17_17_0.C_ON=1'b0;
    defparam buf_dds0_i3_LC_17_17_0.SEQ_MODE=4'b1000;
    defparam buf_dds0_i3_LC_17_17_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i3_LC_17_17_0 (
            .in0(N__56179),
            .in1(N__46915),
            .in2(N__51021),
            .in3(N__48026),
            .lcout(buf_dds0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54423),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i7_LC_17_17_1.C_ON=1'b0;
    defparam acadc_skipCount_i7_LC_17_17_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i7_LC_17_17_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i7_LC_17_17_1 (
            .in0(N__56220),
            .in1(N__44317),
            .in2(N__50322),
            .in3(N__46976),
            .lcout(acadc_skipCount_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54423),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i4_LC_17_17_2.C_ON=1'b0;
    defparam buf_device_acadc_i4_LC_17_17_2.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i4_LC_17_17_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i4_LC_17_17_2 (
            .in0(N__56180),
            .in1(N__44820),
            .in2(N__44197),
            .in3(N__44104),
            .lcout(IAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54423),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds1_305_LC_17_17_3.C_ON=1'b0;
    defparam trig_dds1_305_LC_17_17_3.SEQ_MODE=4'b1000;
    defparam trig_dds1_305_LC_17_17_3.LUT_INIT=16'b0101000110100000;
    LogicCell40 trig_dds1_305_LC_17_17_3 (
            .in0(N__56221),
            .in1(N__44085),
            .in2(N__44032),
            .in3(N__57092),
            .lcout(trig_dds1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54423),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_17_17_4.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_17_17_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_17_17_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_17_17_4 (
            .in0(N__57091),
            .in1(N__45099),
            .in2(N__56292),
            .in3(N__45092),
            .lcout(data_index_9_N_216_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i3_LC_17_18_1.C_ON=1'b0;
    defparam buf_dds1_i3_LC_17_18_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i3_LC_17_18_1.LUT_INIT=16'b1100111110101010;
    LogicCell40 buf_dds1_i3_LC_17_18_1 (
            .in0(N__46945),
            .in1(N__47092),
            .in2(N__57143),
            .in3(N__44970),
            .lcout(buf_dds1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54430),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i3_LC_17_18_5.C_ON=1'b0;
    defparam buf_device_acadc_i3_LC_17_18_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i3_LC_17_18_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i3_LC_17_18_5 (
            .in0(N__56222),
            .in1(N__44819),
            .in2(N__44786),
            .in3(N__44668),
            .lcout(IAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54430),
            .ce(),
            .sr(_gnd_net_));
    defparam i15107_2_lut_2_lut_LC_17_20_6.C_ON=1'b0;
    defparam i15107_2_lut_2_lut_LC_17_20_6.SEQ_MODE=4'b0000;
    defparam i15107_2_lut_2_lut_LC_17_20_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 i15107_2_lut_2_lut_LC_17_20_6 (
            .in0(N__44649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44612),
            .lcout(CONT_SD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_18_3_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_18_3_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_18_3_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_18_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_12182_12183_reset_LC_18_4_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12182_12183_reset_LC_18_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imosi_44_12182_12183_reset_LC_18_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_12182_12183_reset_LC_18_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55601),
            .lcout(\comm_spi.n14601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54283),
            .ce(),
            .sr(N__44577));
    defparam \comm_spi.data_tx_i5_12216_12217_set_LC_18_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12216_12217_set_LC_18_5_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i5_12216_12217_set_LC_18_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_12216_12217_set_LC_18_5_0  (
            .in0(N__44562),
            .in1(N__44535),
            .in2(_gnd_net_),
            .in3(N__44517),
            .lcout(\comm_spi.n14634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52587),
            .ce(),
            .sr(N__44499));
    defparam \comm_spi.data_tx_i6_12220_12221_set_LC_18_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12220_12221_set_LC_18_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i6_12220_12221_set_LC_18_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_12220_12221_set_LC_18_6_0  (
            .in0(N__44487),
            .in1(N__44468),
            .in2(_gnd_net_),
            .in3(N__44457),
            .lcout(\comm_spi.n14638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52531),
            .ce(),
            .sr(N__45375));
    defparam \ADC_VDC.genclk.i19300_4_lut_LC_18_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19300_4_lut_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19300_4_lut_LC_18_7_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i19300_4_lut_LC_18_7_0  (
            .in0(N__48098),
            .in1(N__48191),
            .in2(N__48144),
            .in3(N__48206),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n21446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19039_4_lut_LC_18_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19039_4_lut_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19039_4_lut_LC_18_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i19039_4_lut_LC_18_7_1  (
            .in0(N__45381),
            .in1(N__45393),
            .in2(N__45396),
            .in3(N__45387),
            .lcout(\ADC_VDC.genclk.n21444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_LC_18_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_18_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_LC_18_7_2  (
            .in0(N__48989),
            .in1(N__48902),
            .in2(N__48120),
            .in3(N__48158),
            .lcout(\ADC_VDC.genclk.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_LC_18_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_18_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_LC_18_7_3  (
            .in0(N__48173),
            .in1(N__48920),
            .in2(N__49008),
            .in3(N__48953),
            .lcout(\ADC_VDC.genclk.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_adj_8_LC_18_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_8_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_8_LC_18_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_adj_8_LC_18_7_4  (
            .in0(N__48935),
            .in1(N__49212),
            .in2(N__48974),
            .in3(N__48887),
            .lcout(\ADC_VDC.genclk.n28_adj_1397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_18_7_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_18_7_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_18_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_93_2_lut_LC_18_7_6  (
            .in0(_gnd_net_),
            .in1(N__45259),
            .in2(_gnd_net_),
            .in3(N__55778),
            .lcout(\comm_spi.data_tx_7__N_767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_6_i1_3_lut_LC_18_8_0.C_ON=1'b0;
    defparam mux_137_Mux_6_i1_3_lut_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_6_i1_3_lut_LC_18_8_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_137_Mux_6_i1_3_lut_LC_18_8_0 (
            .in0(N__45338),
            .in1(N__47878),
            .in2(_gnd_net_),
            .in3(N__50793),
            .lcout(),
            .ltout(n1_adj_1588_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i6_LC_18_8_1.C_ON=1'b0;
    defparam comm_tx_buf_i6_LC_18_8_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i6_LC_18_8_1.LUT_INIT=16'b1110111001010000;
    LogicCell40 comm_tx_buf_i6_LC_18_8_1 (
            .in0(N__50604),
            .in1(N__45105),
            .in2(N__45273),
            .in3(N__45570),
            .lcout(comm_tx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54324),
            .ce(N__45233),
            .sr(N__45177));
    defparam mux_137_Mux_6_i2_3_lut_LC_18_8_2.C_ON=1'b0;
    defparam mux_137_Mux_6_i2_3_lut_LC_18_8_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_6_i2_3_lut_LC_18_8_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_6_i2_3_lut_LC_18_8_2 (
            .in0(N__45474),
            .in1(N__45114),
            .in2(_gnd_net_),
            .in3(N__50792),
            .lcout(n2_adj_1589),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19276_2_lut_LC_18_8_4.C_ON=1'b0;
    defparam i19276_2_lut_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam i19276_2_lut_LC_18_8_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19276_2_lut_LC_18_8_4 (
            .in0(_gnd_net_),
            .in1(N__45600),
            .in2(_gnd_net_),
            .in3(N__50791),
            .lcout(),
            .ltout(n21539_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19724_LC_18_8_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19724_LC_18_8_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19724_LC_18_8_5.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_index_1__bdd_4_lut_19724_LC_18_8_5 (
            .in0(N__50603),
            .in1(N__45579),
            .in2(N__45573),
            .in3(N__52411),
            .lcout(n22339),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i0_LC_18_9_0.C_ON=1'b0;
    defparam comm_buf_3__i0_LC_18_9_0.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i0_LC_18_9_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_3__i0_LC_18_9_0 (
            .in0(N__45564),
            .in1(N__51950),
            .in2(_gnd_net_),
            .in3(N__53035),
            .lcout(comm_buf_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam comm_buf_3__i4_LC_18_9_1.C_ON=1'b0;
    defparam comm_buf_3__i4_LC_18_9_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i4_LC_18_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i4_LC_18_9_1 (
            .in0(N__51948),
            .in1(N__46772),
            .in2(_gnd_net_),
            .in3(N__45546),
            .lcout(comm_buf_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam comm_buf_3__i7_LC_18_9_2.C_ON=1'b0;
    defparam comm_buf_3__i7_LC_18_9_2.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i7_LC_18_9_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i7_LC_18_9_2 (
            .in0(N__50409),
            .in1(N__45519),
            .in2(_gnd_net_),
            .in3(N__51945),
            .lcout(comm_buf_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam comm_buf_3__i6_LC_18_9_3.C_ON=1'b0;
    defparam comm_buf_3__i6_LC_18_9_3.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i6_LC_18_9_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i6_LC_18_9_3 (
            .in0(N__51949),
            .in1(N__46461),
            .in2(_gnd_net_),
            .in3(N__45489),
            .lcout(comm_buf_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam comm_buf_3__i5_LC_18_9_4.C_ON=1'b0;
    defparam comm_buf_3__i5_LC_18_9_4.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i5_LC_18_9_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i5_LC_18_9_4 (
            .in0(N__52112),
            .in1(N__45465),
            .in2(_gnd_net_),
            .in3(N__51944),
            .lcout(comm_buf_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam comm_buf_3__i3_LC_18_9_5.C_ON=1'b0;
    defparam comm_buf_3__i3_LC_18_9_5.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i3_LC_18_9_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i3_LC_18_9_5 (
            .in0(N__51947),
            .in1(N__51108),
            .in2(_gnd_net_),
            .in3(N__45444),
            .lcout(comm_buf_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam comm_buf_3__i2_LC_18_9_6.C_ON=1'b0;
    defparam comm_buf_3__i2_LC_18_9_6.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i2_LC_18_9_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i2_LC_18_9_6 (
            .in0(N__47236),
            .in1(N__45420),
            .in2(_gnd_net_),
            .in3(N__51943),
            .lcout(comm_buf_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam comm_buf_3__i1_LC_18_9_7.C_ON=1'b0;
    defparam comm_buf_3__i1_LC_18_9_7.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i1_LC_18_9_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i1_LC_18_9_7 (
            .in0(N__51946),
            .in1(N__45795),
            .in2(_gnd_net_),
            .in3(N__45696),
            .lcout(comm_buf_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54336),
            .ce(N__45651),
            .sr(N__45642));
    defparam i2_3_lut_adj_78_LC_18_10_0.C_ON=1'b0;
    defparam i2_3_lut_adj_78_LC_18_10_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_78_LC_18_10_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 i2_3_lut_adj_78_LC_18_10_0 (
            .in0(N__49793),
            .in1(N__49748),
            .in2(_gnd_net_),
            .in3(N__49712),
            .lcout(n20878),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19274_2_lut_LC_18_10_1.C_ON=1'b0;
    defparam i19274_2_lut_LC_18_10_1.SEQ_MODE=4'b0000;
    defparam i19274_2_lut_LC_18_10_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19274_2_lut_LC_18_10_1 (
            .in0(_gnd_net_),
            .in1(N__45631),
            .in2(_gnd_net_),
            .in3(N__49800),
            .lcout(),
            .ltout(n21352_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_LC_18_10_2.C_ON=1'b0;
    defparam i19_4_lut_LC_18_10_2.SEQ_MODE=4'b0000;
    defparam i19_4_lut_LC_18_10_2.LUT_INIT=16'b1000000011010101;
    LogicCell40 i19_4_lut_LC_18_10_2 (
            .in0(N__51924),
            .in1(N__50752),
            .in2(N__45657),
            .in3(N__45954),
            .lcout(),
            .ltout(n12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_272_LC_18_10_3.C_ON=1'b0;
    defparam i1_3_lut_adj_272_LC_18_10_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_272_LC_18_10_3.LUT_INIT=16'b1100110011000000;
    LogicCell40 i1_3_lut_adj_272_LC_18_10_3 (
            .in0(_gnd_net_),
            .in1(N__45915),
            .in2(N__45654),
            .in3(N__45880),
            .lcout(n12136),
            .ltout(n12136_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12358_2_lut_LC_18_10_4.C_ON=1'b0;
    defparam i12358_2_lut_LC_18_10_4.SEQ_MODE=4'b0000;
    defparam i12358_2_lut_LC_18_10_4.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12358_2_lut_LC_18_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45645),
            .in3(N__56867),
            .lcout(n14771),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_50_LC_18_10_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_50_LC_18_10_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_50_LC_18_10_5.LUT_INIT=16'b0000000000010000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_50_LC_18_10_5 (
            .in0(N__50026),
            .in1(N__52388),
            .in2(N__49877),
            .in3(N__52243),
            .lcout(n18991),
            .ltout(n18991_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_265_LC_18_10_6.C_ON=1'b0;
    defparam i1_4_lut_adj_265_LC_18_10_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_265_LC_18_10_6.LUT_INIT=16'b0001000011111111;
    LogicCell40 i1_4_lut_adj_265_LC_18_10_6 (
            .in0(N__45632),
            .in1(N__50751),
            .in2(N__45606),
            .in3(N__51999),
            .lcout(),
            .ltout(n4_adj_1545_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_266_LC_18_10_7.C_ON=1'b0;
    defparam i1_4_lut_adj_266_LC_18_10_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_266_LC_18_10_7.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_266_LC_18_10_7 (
            .in0(N__49665),
            .in1(N__45914),
            .in2(N__45603),
            .in3(N__45879),
            .lcout(n11961),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_47_LC_18_11_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_47_LC_18_11_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_47_LC_18_11_0.LUT_INIT=16'b0010001000000000;
    LogicCell40 i1_2_lut_3_lut_adj_47_LC_18_11_0 (
            .in0(N__50584),
            .in1(N__49503),
            .in2(_gnd_net_),
            .in3(N__49292),
            .lcout(n18993),
            .ltout(n18993_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_276_LC_18_11_1.C_ON=1'b0;
    defparam i19_4_lut_adj_276_LC_18_11_1.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_276_LC_18_11_1.LUT_INIT=16'b1100000001010101;
    LogicCell40 i19_4_lut_adj_276_LC_18_11_1 (
            .in0(N__45953),
            .in1(N__50786),
            .in2(N__46095),
            .in3(N__51917),
            .lcout(n12_adj_1605),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_269_LC_18_11_2.C_ON=1'b0;
    defparam i1_3_lut_adj_269_LC_18_11_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_269_LC_18_11_2.LUT_INIT=16'b1111000010100000;
    LogicCell40 i1_3_lut_adj_269_LC_18_11_2 (
            .in0(N__45876),
            .in1(_gnd_net_),
            .in2(N__45920),
            .in3(N__49236),
            .lcout(n11991),
            .ltout(n11991_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12344_2_lut_LC_18_11_3.C_ON=1'b0;
    defparam i12344_2_lut_LC_18_11_3.SEQ_MODE=4'b0000;
    defparam i12344_2_lut_LC_18_11_3.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12344_2_lut_LC_18_11_3 (
            .in0(N__57066),
            .in1(_gnd_net_),
            .in2(N__46086),
            .in3(_gnd_net_),
            .lcout(n14757),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_48_LC_18_11_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_48_LC_18_11_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_48_LC_18_11_4.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_adj_48_LC_18_11_4 (
            .in0(N__49587),
            .in1(N__55408),
            .in2(_gnd_net_),
            .in3(N__57065),
            .lcout(n20843),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i7_LC_18_11_5.C_ON=1'b0;
    defparam comm_cmd_i7_LC_18_11_5.SEQ_MODE=4'b1000;
    defparam comm_cmd_i7_LC_18_11_5.LUT_INIT=16'b1010000011001100;
    LogicCell40 comm_cmd_i7_LC_18_11_5 (
            .in0(N__46083),
            .in1(N__52254),
            .in2(N__50412),
            .in3(N__46014),
            .lcout(comm_cmd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54364),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_273_LC_18_11_6.C_ON=1'b0;
    defparam i19_4_lut_adj_273_LC_18_11_6.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_273_LC_18_11_6.LUT_INIT=16'b0001101100010001;
    LogicCell40 i19_4_lut_adj_273_LC_18_11_6 (
            .in0(N__51916),
            .in1(N__45952),
            .in2(N__50798),
            .in3(N__45933),
            .lcout(),
            .ltout(n12_adj_1635_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_274_LC_18_11_7.C_ON=1'b0;
    defparam i1_3_lut_adj_274_LC_18_11_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_274_LC_18_11_7.LUT_INIT=16'b1100110011000000;
    LogicCell40 i1_3_lut_adj_274_LC_18_11_7 (
            .in0(_gnd_net_),
            .in1(N__45910),
            .in2(N__45885),
            .in3(N__45877),
            .lcout(n12178),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19639_LC_18_12_0.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19639_LC_18_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19639_LC_18_12_0.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_2__bdd_4_lut_19639_LC_18_12_0 (
            .in0(N__54757),
            .in1(N__53611),
            .in2(N__46557),
            .in3(N__46470),
            .lcout(),
            .ltout(n22225_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22225_bdd_4_lut_LC_18_12_1.C_ON=1'b0;
    defparam n22225_bdd_4_lut_LC_18_12_1.SEQ_MODE=4'b0000;
    defparam n22225_bdd_4_lut_LC_18_12_1.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22225_bdd_4_lut_LC_18_12_1 (
            .in0(N__47007),
            .in1(N__46287),
            .in2(N__46539),
            .in3(N__54758),
            .lcout(n22228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_6_i26_3_lut_LC_18_12_2.C_ON=1'b0;
    defparam mux_129_Mux_6_i26_3_lut_LC_18_12_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i26_3_lut_LC_18_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_6_i26_3_lut_LC_18_12_2 (
            .in0(N__46536),
            .in1(N__57805),
            .in2(_gnd_net_),
            .in3(N__46515),
            .lcout(),
            .ltout(n26_adj_1507_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18568_4_lut_LC_18_12_3.C_ON=1'b0;
    defparam i18568_4_lut_LC_18_12_3.SEQ_MODE=4'b0000;
    defparam i18568_4_lut_LC_18_12_3.LUT_INIT=16'b1110111011110000;
    LogicCell40 i18568_4_lut_LC_18_12_3 (
            .in0(N__57807),
            .in1(N__46485),
            .in2(N__46473),
            .in3(N__55153),
            .lcout(n21178),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i6_LC_18_12_4.C_ON=1'b0;
    defparam comm_buf_1__i6_LC_18_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i6_LC_18_12_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_1__i6_LC_18_12_4 (
            .in0(N__51860),
            .in1(N__46463),
            .in2(_gnd_net_),
            .in3(N__46383),
            .lcout(comm_buf_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54377),
            .ce(N__51356),
            .sr(N__51257));
    defparam mux_129_Mux_6_i19_3_lut_LC_18_12_5.C_ON=1'b0;
    defparam mux_129_Mux_6_i19_3_lut_LC_18_12_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i19_3_lut_LC_18_12_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_6_i19_3_lut_LC_18_12_5 (
            .in0(N__57806),
            .in1(N__46377),
            .in2(_gnd_net_),
            .in3(N__46349),
            .lcout(),
            .ltout(n19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18436_3_lut_LC_18_12_6.C_ON=1'b0;
    defparam i18436_3_lut_LC_18_12_6.SEQ_MODE=4'b0000;
    defparam i18436_3_lut_LC_18_12_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 i18436_3_lut_LC_18_12_6 (
            .in0(N__55154),
            .in1(_gnd_net_),
            .in2(N__46320),
            .in3(N__46317),
            .lcout(n21046),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22231_bdd_4_lut_LC_18_13_0.C_ON=1'b0;
    defparam n22231_bdd_4_lut_LC_18_13_0.SEQ_MODE=4'b0000;
    defparam n22231_bdd_4_lut_LC_18_13_0.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22231_bdd_4_lut_LC_18_13_0 (
            .in0(N__53791),
            .in1(N__46281),
            .in2(N__46269),
            .in3(N__46230),
            .lcout(n22234),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i26_3_lut_LC_18_13_2.C_ON=1'b0;
    defparam mux_129_Mux_4_i26_3_lut_LC_18_13_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i26_3_lut_LC_18_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_4_i26_3_lut_LC_18_13_2 (
            .in0(N__46218),
            .in1(N__57817),
            .in2(_gnd_net_),
            .in3(N__46197),
            .lcout(),
            .ltout(n26_adj_1512_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19714_LC_18_13_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19714_LC_18_13_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19714_LC_18_13_3.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19714_LC_18_13_3 (
            .in0(N__53883),
            .in1(N__55157),
            .in2(N__46854),
            .in3(N__53792),
            .lcout(),
            .ltout(n22351_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22351_bdd_4_lut_LC_18_13_4.C_ON=1'b0;
    defparam n22351_bdd_4_lut_LC_18_13_4.SEQ_MODE=4'b0000;
    defparam n22351_bdd_4_lut_LC_18_13_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22351_bdd_4_lut_LC_18_13_4 (
            .in0(N__53793),
            .in1(N__46851),
            .in2(N__46824),
            .in3(N__46821),
            .lcout(),
            .ltout(n22354_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1555570_i1_3_lut_LC_18_13_5.C_ON=1'b0;
    defparam i1555570_i1_3_lut_LC_18_13_5.SEQ_MODE=4'b0000;
    defparam i1555570_i1_3_lut_LC_18_13_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1555570_i1_3_lut_LC_18_13_5 (
            .in0(_gnd_net_),
            .in1(N__46797),
            .in2(N__46791),
            .in3(N__54744),
            .lcout(),
            .ltout(n30_adj_1513_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i4_LC_18_13_6.C_ON=1'b0;
    defparam comm_buf_1__i4_LC_18_13_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i4_LC_18_13_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i4_LC_18_13_6 (
            .in0(N__46788),
            .in1(_gnd_net_),
            .in2(N__46689),
            .in3(N__52008),
            .lcout(comm_buf_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54391),
            .ce(N__51384),
            .sr(N__51283));
    defparam comm_cmd_1__bdd_4_lut_19598_LC_18_14_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19598_LC_18_14_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19598_LC_18_14_1.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19598_LC_18_14_1 (
            .in0(N__46686),
            .in1(N__55155),
            .in2(N__46674),
            .in3(N__53787),
            .lcout(),
            .ltout(n22207_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22207_bdd_4_lut_LC_18_14_2.C_ON=1'b0;
    defparam n22207_bdd_4_lut_LC_18_14_2.SEQ_MODE=4'b0000;
    defparam n22207_bdd_4_lut_LC_18_14_2.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22207_bdd_4_lut_LC_18_14_2 (
            .in0(N__53788),
            .in1(N__46640),
            .in2(N__46617),
            .in3(N__46863),
            .lcout(n22210),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_LC_18_14_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_LC_18_14_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_LC_18_14_3.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_LC_18_14_3 (
            .in0(N__55156),
            .in1(N__47103),
            .in2(N__52722),
            .in3(N__53789),
            .lcout(),
            .ltout(n22429_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22429_bdd_4_lut_LC_18_14_4.C_ON=1'b0;
    defparam n22429_bdd_4_lut_LC_18_14_4.SEQ_MODE=4'b0000;
    defparam n22429_bdd_4_lut_LC_18_14_4.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22429_bdd_4_lut_LC_18_14_4 (
            .in0(N__53790),
            .in1(N__46614),
            .in2(N__46587),
            .in3(N__46584),
            .lcout(),
            .ltout(n22432_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1554364_i1_3_lut_LC_18_14_5.C_ON=1'b0;
    defparam i1554364_i1_3_lut_LC_18_14_5.SEQ_MODE=4'b0000;
    defparam i1554364_i1_3_lut_LC_18_14_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1554364_i1_3_lut_LC_18_14_5 (
            .in0(_gnd_net_),
            .in1(N__47253),
            .in2(N__47247),
            .in3(N__54764),
            .lcout(),
            .ltout(n30_adj_1520_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i2_LC_18_14_6.C_ON=1'b0;
    defparam comm_buf_1__i2_LC_18_14_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i2_LC_18_14_6.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_1__i2_LC_18_14_6 (
            .in0(N__51998),
            .in1(N__47243),
            .in2(N__47151),
            .in3(_gnd_net_),
            .lcout(comm_buf_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54403),
            .ce(N__51374),
            .sr(N__51300));
    defparam mux_129_Mux_2_i26_3_lut_LC_18_15_0.C_ON=1'b0;
    defparam mux_129_Mux_2_i26_3_lut_LC_18_15_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i26_3_lut_LC_18_15_0.LUT_INIT=16'b1010111110100000;
    LogicCell40 mux_129_Mux_2_i26_3_lut_LC_18_15_0 (
            .in0(N__47148),
            .in1(_gnd_net_),
            .in2(N__57819),
            .in3(N__47127),
            .lcout(n26_adj_1519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15326_2_lut_3_lut_LC_18_15_1.C_ON=1'b0;
    defparam i15326_2_lut_3_lut_LC_18_15_1.SEQ_MODE=4'b0000;
    defparam i15326_2_lut_3_lut_LC_18_15_1.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15326_2_lut_3_lut_LC_18_15_1 (
            .in0(N__50999),
            .in1(N__55480),
            .in2(_gnd_net_),
            .in3(N__52027),
            .lcout(n14_adj_1585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_18_15_3.C_ON=1'b0;
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_18_15_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_18_15_3.LUT_INIT=16'b1111111100110011;
    LogicCell40 comm_cmd_6__I_0_368_i8_2_lut_LC_18_15_3 (
            .in0(_gnd_net_),
            .in1(N__55148),
            .in2(_gnd_net_),
            .in3(N__53766),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18435_3_lut_LC_18_15_4.C_ON=1'b0;
    defparam i18435_3_lut_LC_18_15_4.SEQ_MODE=4'b0000;
    defparam i18435_3_lut_LC_18_15_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18435_3_lut_LC_18_15_4 (
            .in0(N__47039),
            .in1(N__47016),
            .in2(_gnd_net_),
            .in3(N__55150),
            .lcout(n21045),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18444_3_lut_LC_18_15_5.C_ON=1'b0;
    defparam i18444_3_lut_LC_18_15_5.SEQ_MODE=4'b0000;
    defparam i18444_3_lut_LC_18_15_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18444_3_lut_LC_18_15_5 (
            .in0(N__55149),
            .in1(N__46998),
            .in2(_gnd_net_),
            .in3(N__46977),
            .lcout(n21054),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_3_i16_3_lut_LC_18_15_7.C_ON=1'b0;
    defparam mux_129_Mux_3_i16_3_lut_LC_18_15_7.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i16_3_lut_LC_18_15_7.LUT_INIT=16'b1111001111000000;
    LogicCell40 mux_129_Mux_3_i16_3_lut_LC_18_15_7 (
            .in0(_gnd_net_),
            .in1(N__57763),
            .in2(N__46952),
            .in3(N__46916),
            .lcout(n16_adj_1514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i16_3_lut_LC_18_16_1.C_ON=1'b0;
    defparam mux_129_Mux_2_i16_3_lut_LC_18_16_1.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i16_3_lut_LC_18_16_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_2_i16_3_lut_LC_18_16_1 (
            .in0(N__46892),
            .in1(N__47914),
            .in2(_gnd_net_),
            .in3(N__57824),
            .lcout(n16_adj_1517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i2_LC_18_16_4.C_ON=1'b0;
    defparam buf_dds0_i2_LC_18_16_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i2_LC_18_16_4.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_dds0_i2_LC_18_16_4 (
            .in0(N__47915),
            .in1(N__56451),
            .in2(N__48067),
            .in3(N__48011),
            .lcout(buf_dds0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54424),
            .ce(),
            .sr(_gnd_net_));
    defparam i15342_2_lut_3_lut_LC_18_17_0.C_ON=1'b0;
    defparam i15342_2_lut_3_lut_LC_18_17_0.SEQ_MODE=4'b0000;
    defparam i15342_2_lut_3_lut_LC_18_17_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15342_2_lut_3_lut_LC_18_17_0 (
            .in0(N__47891),
            .in1(N__51997),
            .in2(_gnd_net_),
            .in3(N__55541),
            .lcout(n14_adj_1552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6419_3_lut_LC_18_18_2.C_ON=1'b0;
    defparam i6419_3_lut_LC_18_18_2.SEQ_MODE=4'b0000;
    defparam i6419_3_lut_LC_18_18_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6419_3_lut_LC_18_18_2 (
            .in0(N__47763),
            .in1(N__47727),
            .in2(_gnd_net_),
            .in3(N__47701),
            .lcout(n8_adj_1567),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_18_19_5.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_18_19_5.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_18_19_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_18_19_5 (
            .in0(N__57138),
            .in1(N__47633),
            .in2(N__56477),
            .in3(N__47621),
            .lcout(data_index_9_N_216_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19407_2_lut_4_lut_LC_19_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19407_2_lut_4_lut_LC_19_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19407_2_lut_4_lut_LC_19_5_0 .LUT_INIT=16'b0010011111111111;
    LogicCell40 \ADC_VDC.genclk.i19407_2_lut_4_lut_LC_19_5_0  (
            .in0(N__58010),
            .in1(N__53351),
            .in2(N__58160),
            .in3(N__52908),
            .lcout(\ADC_VDC.genclk.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19334_2_lut_LC_19_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19334_2_lut_LC_19_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19334_2_lut_LC_19_5_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ADC_VDC.genclk.i19334_2_lut_LC_19_5_4  (
            .in0(_gnd_net_),
            .in1(N__52907),
            .in2(_gnd_net_),
            .in3(N__58006),
            .lcout(\ADC_VDC.genclk.n11735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16159_4_lut_LC_19_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i16159_4_lut_LC_19_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16159_4_lut_LC_19_5_5 .LUT_INIT=16'b1001100010111010;
    LogicCell40 \ADC_VDC.i16159_4_lut_LC_19_5_5  (
            .in0(N__48786),
            .in1(N__48581),
            .in2(N__47262),
            .in3(N__48356),
            .lcout(\ADC_VDC.n11750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_LC_19_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_LC_19_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_LC_19_5_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_LC_19_5_6  (
            .in0(_gnd_net_),
            .in1(N__47493),
            .in2(_gnd_net_),
            .in3(N__47363),
            .lcout(\ADC_VDC.n62 ),
            .ltout(\ADC_VDC.n62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i24_4_lut_LC_19_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.i24_4_lut_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i24_4_lut_LC_19_5_7 .LUT_INIT=16'b1001100010111010;
    LogicCell40 \ADC_VDC.i24_4_lut_LC_19_5_7  (
            .in0(N__48785),
            .in1(N__48580),
            .in2(N__48360),
            .in3(N__48355),
            .lcout(\ADC_VDC.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12196_12197_set_LC_19_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12196_12197_set_LC_19_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_rx_i0_12196_12197_set_LC_19_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.data_rx_i0_12196_12197_set_LC_19_6_0  (
            .in0(N__52971),
            .in1(N__52948),
            .in2(_gnd_net_),
            .in3(N__55902),
            .lcout(\comm_spi.n14614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52570),
            .ce(),
            .sr(N__52920));
    defparam \ADC_VDC.genclk.t0off_i0_LC_19_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i0_LC_19_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i0_LC_19_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i0_LC_19_7_0  (
            .in0(_gnd_net_),
            .in1(N__48207),
            .in2(_gnd_net_),
            .in3(N__48195),
            .lcout(\ADC_VDC.genclk.t0off_0 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\ADC_VDC.genclk.n19709 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i1_LC_19_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i1_LC_19_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i1_LC_19_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i1_LC_19_7_1  (
            .in0(_gnd_net_),
            .in1(N__48192),
            .in2(N__58522),
            .in3(N__48180),
            .lcout(\ADC_VDC.genclk.t0off_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19709 ),
            .carryout(\ADC_VDC.genclk.n19710 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i2_LC_19_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i2_LC_19_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i2_LC_19_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i2_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(N__58447),
            .in2(N__48177),
            .in3(N__48162),
            .lcout(\ADC_VDC.genclk.t0off_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19710 ),
            .carryout(\ADC_VDC.genclk.n19711 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i3_LC_19_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i3_LC_19_7_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0off_i3_LC_19_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i3_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(N__48159),
            .in2(N__58523),
            .in3(N__48147),
            .lcout(\ADC_VDC.genclk.t0off_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19711 ),
            .carryout(\ADC_VDC.genclk.n19712 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i4_LC_19_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i4_LC_19_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i4_LC_19_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i4_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(N__58451),
            .in2(N__48143),
            .in3(N__48123),
            .lcout(\ADC_VDC.genclk.t0off_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19712 ),
            .carryout(\ADC_VDC.genclk.n19713 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i5_LC_19_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i5_LC_19_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i5_LC_19_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i5_LC_19_7_5  (
            .in0(_gnd_net_),
            .in1(N__48119),
            .in2(N__58524),
            .in3(N__48105),
            .lcout(\ADC_VDC.genclk.t0off_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19713 ),
            .carryout(\ADC_VDC.genclk.n19714 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i6_LC_19_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i6_LC_19_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i6_LC_19_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i6_LC_19_7_6  (
            .in0(_gnd_net_),
            .in1(N__58455),
            .in2(N__48102),
            .in3(N__48087),
            .lcout(\ADC_VDC.genclk.t0off_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19714 ),
            .carryout(\ADC_VDC.genclk.n19715 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i7_LC_19_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i7_LC_19_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i7_LC_19_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i7_LC_19_7_7  (
            .in0(_gnd_net_),
            .in1(N__49007),
            .in2(N__58525),
            .in3(N__48993),
            .lcout(\ADC_VDC.genclk.t0off_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19715 ),
            .carryout(\ADC_VDC.genclk.n19716 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__49197),
            .sr(N__58243));
    defparam \ADC_VDC.genclk.t0off_i8_LC_19_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i8_LC_19_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i8_LC_19_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i8_LC_19_8_0  (
            .in0(_gnd_net_),
            .in1(N__48990),
            .in2(N__58576),
            .in3(N__48978),
            .lcout(\ADC_VDC.genclk.t0off_8 ),
            .ltout(),
            .carryin(bfn_19_8_0_),
            .carryout(\ADC_VDC.genclk.n19717 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam \ADC_VDC.genclk.t0off_i9_LC_19_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i9_LC_19_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i9_LC_19_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i9_LC_19_8_1  (
            .in0(_gnd_net_),
            .in1(N__58541),
            .in2(N__48975),
            .in3(N__48957),
            .lcout(\ADC_VDC.genclk.t0off_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19717 ),
            .carryout(\ADC_VDC.genclk.n19718 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam \ADC_VDC.genclk.t0off_i10_LC_19_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i10_LC_19_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i10_LC_19_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i10_LC_19_8_2  (
            .in0(_gnd_net_),
            .in1(N__48954),
            .in2(N__58573),
            .in3(N__48942),
            .lcout(\ADC_VDC.genclk.t0off_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19718 ),
            .carryout(\ADC_VDC.genclk.n19719 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam \ADC_VDC.genclk.t0off_i11_LC_19_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i11_LC_19_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i11_LC_19_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i11_LC_19_8_3  (
            .in0(_gnd_net_),
            .in1(N__58529),
            .in2(N__48939),
            .in3(N__48924),
            .lcout(\ADC_VDC.genclk.t0off_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19719 ),
            .carryout(\ADC_VDC.genclk.n19720 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam \ADC_VDC.genclk.t0off_i12_LC_19_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i12_LC_19_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i12_LC_19_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i12_LC_19_8_4  (
            .in0(_gnd_net_),
            .in1(N__48921),
            .in2(N__58574),
            .in3(N__48909),
            .lcout(\ADC_VDC.genclk.t0off_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19720 ),
            .carryout(\ADC_VDC.genclk.n19721 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam \ADC_VDC.genclk.t0off_i13_LC_19_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i13_LC_19_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i13_LC_19_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i13_LC_19_8_5  (
            .in0(_gnd_net_),
            .in1(N__58533),
            .in2(N__48906),
            .in3(N__48891),
            .lcout(\ADC_VDC.genclk.t0off_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19721 ),
            .carryout(\ADC_VDC.genclk.n19722 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam \ADC_VDC.genclk.t0off_i14_LC_19_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i14_LC_19_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i14_LC_19_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i14_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(N__48888),
            .in2(N__58575),
            .in3(N__48876),
            .lcout(\ADC_VDC.genclk.t0off_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19722 ),
            .carryout(\ADC_VDC.genclk.n19723 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam \ADC_VDC.genclk.t0off_i15_LC_19_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0off_i15_LC_19_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i15_LC_19_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0off_i15_LC_19_8_7  (
            .in0(N__49211),
            .in1(N__58537),
            .in2(_gnd_net_),
            .in3(N__49215),
            .lcout(\ADC_VDC.genclk.t0off_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__49196),
            .sr(N__58263));
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_19_9_0.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_19_9_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_19_9_0.LUT_INIT=16'b1111101011011000;
    LogicCell40 comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_19_9_0 (
            .in0(N__55350),
            .in1(N__49017),
            .in2(N__49026),
            .in3(N__49176),
            .lcout(n17815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_LC_19_9_1.C_ON=1'b0;
    defparam i1_4_lut_4_lut_LC_19_9_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_LC_19_9_1.LUT_INIT=16'b0010011000000000;
    LogicCell40 i1_4_lut_4_lut_LC_19_9_1 (
            .in0(N__51724),
            .in1(N__55351),
            .in2(N__50046),
            .in3(N__49881),
            .lcout(),
            .ltout(n21_adj_1598_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19391_4_lut_LC_19_9_2.C_ON=1'b0;
    defparam i19391_4_lut_LC_19_9_2.SEQ_MODE=4'b0000;
    defparam i19391_4_lut_LC_19_9_2.LUT_INIT=16'b0000101111111111;
    LogicCell40 i19391_4_lut_LC_19_9_2 (
            .in0(N__55352),
            .in1(N__49128),
            .in2(N__49113),
            .in3(N__49110),
            .lcout(n18_adj_1619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i32_4_lut_LC_19_9_3.C_ON=1'b0;
    defparam i32_4_lut_LC_19_9_3.SEQ_MODE=4'b0000;
    defparam i32_4_lut_LC_19_9_3.LUT_INIT=16'b1110101001000000;
    LogicCell40 i32_4_lut_LC_19_9_3 (
            .in0(N__51725),
            .in1(N__55353),
            .in2(N__49674),
            .in3(N__49092),
            .lcout(),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i2_LC_19_9_4.C_ON=1'b0;
    defparam comm_state_i2_LC_19_9_4.SEQ_MODE=4'b1000;
    defparam comm_state_i2_LC_19_9_4.LUT_INIT=16'b1000100011111000;
    LogicCell40 comm_state_i2_LC_19_9_4 (
            .in0(N__50058),
            .in1(N__49050),
            .in2(N__49035),
            .in3(N__49464),
            .lcout(comm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54350),
            .ce(N__49032),
            .sr(N__57118));
    defparam i11712_2_lut_LC_19_9_5.C_ON=1'b0;
    defparam i11712_2_lut_LC_19_9_5.SEQ_MODE=4'b0000;
    defparam i11712_2_lut_LC_19_9_5.LUT_INIT=16'b1111111111110000;
    LogicCell40 i11712_2_lut_LC_19_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49494),
            .in3(N__51721),
            .lcout(n14130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_318_LC_19_9_6.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_318_LC_19_9_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_318_LC_19_9_6.LUT_INIT=16'b1011111111111011;
    LogicCell40 i1_2_lut_4_lut_adj_318_LC_19_9_6 (
            .in0(N__52428),
            .in1(N__51723),
            .in2(N__54459),
            .in3(N__52410),
            .lcout(n20880),
            .ltout(n20880_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i33_3_lut_LC_19_9_7.C_ON=1'b0;
    defparam i33_3_lut_LC_19_9_7.SEQ_MODE=4'b0000;
    defparam i33_3_lut_LC_19_9_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 i33_3_lut_LC_19_9_7 (
            .in0(N__49463),
            .in1(_gnd_net_),
            .in2(N__49011),
            .in3(N__51722),
            .lcout(n12_adj_1548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_19_10_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_19_10_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_19_10_0.LUT_INIT=16'b0000001000000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_19_10_0 (
            .in0(N__52409),
            .in1(N__52244),
            .in2(N__50051),
            .in3(N__49867),
            .lcout(n18984),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19308_2_lut_3_lut_LC_19_10_1.C_ON=1'b0;
    defparam i19308_2_lut_3_lut_LC_19_10_1.SEQ_MODE=4'b0000;
    defparam i19308_2_lut_3_lut_LC_19_10_1.LUT_INIT=16'b0000000000100010;
    LogicCell40 i19308_2_lut_3_lut_LC_19_10_1 (
            .in0(N__49794),
            .in1(N__49749),
            .in2(_gnd_net_),
            .in3(N__49713),
            .lcout(n21546),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_19_10_2.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_19_10_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_19_10_2.LUT_INIT=16'b1111111111111101;
    LogicCell40 i1_3_lut_4_lut_LC_19_10_2 (
            .in0(N__55348),
            .in1(N__56852),
            .in2(N__51995),
            .in3(N__49279),
            .lcout(n12092),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_281_LC_19_10_4.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_281_LC_19_10_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_281_LC_19_10_4.LUT_INIT=16'b1101111111011101;
    LogicCell40 i1_3_lut_4_lut_adj_281_LC_19_10_4 (
            .in0(N__55349),
            .in1(N__56853),
            .in2(N__51996),
            .in3(N__49281),
            .lcout(),
            .ltout(n11853_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_121_LC_19_10_5.C_ON=1'b0;
    defparam i1_4_lut_adj_121_LC_19_10_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_121_LC_19_10_5.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_adj_121_LC_19_10_5 (
            .in0(N__49656),
            .in1(N__49623),
            .in2(N__49605),
            .in3(N__49585),
            .lcout(n11860),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19318_3_lut_4_lut_LC_19_10_6.C_ON=1'b0;
    defparam i19318_3_lut_4_lut_LC_19_10_6.SEQ_MODE=4'b0000;
    defparam i19318_3_lut_4_lut_LC_19_10_6.LUT_INIT=16'b0001000000000000;
    LogicCell40 i19318_3_lut_4_lut_LC_19_10_6 (
            .in0(N__50602),
            .in1(N__49492),
            .in2(N__50799),
            .in3(N__49293),
            .lcout(),
            .ltout(n21339_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i42_4_lut_LC_19_10_7.C_ON=1'b0;
    defparam i42_4_lut_LC_19_10_7.SEQ_MODE=4'b0000;
    defparam i42_4_lut_LC_19_10_7.LUT_INIT=16'b1111000010001000;
    LogicCell40 i42_4_lut_LC_19_10_7 (
            .in0(N__49280),
            .in1(N__49254),
            .in2(N__49239),
            .in3(N__51909),
            .lcout(n38_adj_1608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19674_LC_19_11_0.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19674_LC_19_11_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19674_LC_19_11_0.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_2__bdd_4_lut_19674_LC_19_11_0 (
            .in0(N__54759),
            .in1(N__53767),
            .in2(N__49230),
            .in3(N__50418),
            .lcout(),
            .ltout(n22267_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22267_bdd_4_lut_LC_19_11_1.C_ON=1'b0;
    defparam n22267_bdd_4_lut_LC_19_11_1.SEQ_MODE=4'b0000;
    defparam n22267_bdd_4_lut_LC_19_11_1.LUT_INIT=16'b1111000010101100;
    LogicCell40 n22267_bdd_4_lut_LC_19_11_1 (
            .in0(N__50160),
            .in1(N__52134),
            .in2(N__50481),
            .in3(N__54760),
            .lcout(n22270),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i26_3_lut_LC_19_11_2.C_ON=1'b0;
    defparam mux_129_Mux_7_i26_3_lut_LC_19_11_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i26_3_lut_LC_19_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_7_i26_3_lut_LC_19_11_2 (
            .in0(N__50478),
            .in1(N__50457),
            .in2(_gnd_net_),
            .in3(N__57651),
            .lcout(),
            .ltout(n26_adj_1502_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18445_4_lut_LC_19_11_3.C_ON=1'b0;
    defparam i18445_4_lut_LC_19_11_3.SEQ_MODE=4'b0000;
    defparam i18445_4_lut_LC_19_11_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18445_4_lut_LC_19_11_3 (
            .in0(N__57653),
            .in1(N__50433),
            .in2(N__50421),
            .in3(N__55233),
            .lcout(n21055),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i7_LC_19_11_4.C_ON=1'b0;
    defparam comm_buf_1__i7_LC_19_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i7_LC_19_11_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i7_LC_19_11_4 (
            .in0(N__50408),
            .in1(N__52007),
            .in2(_gnd_net_),
            .in3(N__50328),
            .lcout(comm_buf_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54378),
            .ce(N__51357),
            .sr(N__51306));
    defparam mux_129_Mux_7_i19_3_lut_LC_19_11_5.C_ON=1'b0;
    defparam mux_129_Mux_7_i19_3_lut_LC_19_11_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i19_3_lut_LC_19_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_7_i19_3_lut_LC_19_11_5 (
            .in0(N__57652),
            .in1(N__50238),
            .in2(_gnd_net_),
            .in3(N__50216),
            .lcout(),
            .ltout(n19_adj_1503_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18439_3_lut_LC_19_11_6.C_ON=1'b0;
    defparam i18439_3_lut_LC_19_11_6.SEQ_MODE=4'b0000;
    defparam i18439_3_lut_LC_19_11_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 i18439_3_lut_LC_19_11_6 (
            .in0(N__55234),
            .in1(_gnd_net_),
            .in2(N__50187),
            .in3(N__50184),
            .lcout(n21049),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18517_3_lut_LC_19_12_0.C_ON=1'b0;
    defparam i18517_3_lut_LC_19_12_0.SEQ_MODE=4'b0000;
    defparam i18517_3_lut_LC_19_12_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 i18517_3_lut_LC_19_12_0 (
            .in0(N__50154),
            .in1(N__50889),
            .in2(N__55212),
            .in3(_gnd_net_),
            .lcout(n21127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18522_3_lut_LC_19_12_1.C_ON=1'b0;
    defparam i18522_3_lut_LC_19_12_1.SEQ_MODE=4'b0000;
    defparam i18522_3_lut_LC_19_12_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 i18522_3_lut_LC_19_12_1 (
            .in0(N__50124),
            .in1(N__55145),
            .in2(_gnd_net_),
            .in3(N__50088),
            .lcout(),
            .ltout(n21132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19788_LC_19_12_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19788_LC_19_12_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19788_LC_19_12_2.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_2__bdd_4_lut_19788_LC_19_12_2 (
            .in0(N__54761),
            .in1(N__53612),
            .in2(N__51126),
            .in3(N__50817),
            .lcout(),
            .ltout(n22333_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22333_bdd_4_lut_LC_19_12_3.C_ON=1'b0;
    defparam n22333_bdd_4_lut_LC_19_12_3.SEQ_MODE=4'b0000;
    defparam n22333_bdd_4_lut_LC_19_12_3.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22333_bdd_4_lut_LC_19_12_3 (
            .in0(N__52746),
            .in1(N__51123),
            .in2(N__51117),
            .in3(N__54762),
            .lcout(),
            .ltout(n22336_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i3_LC_19_12_4.C_ON=1'b0;
    defparam comm_buf_1__i3_LC_19_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i3_LC_19_12_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i3_LC_19_12_4 (
            .in0(_gnd_net_),
            .in1(N__51109),
            .in2(N__51024),
            .in3(N__51925),
            .lcout(comm_buf_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54392),
            .ce(N__51358),
            .sr(N__51299));
    defparam mux_129_Mux_3_i19_3_lut_LC_19_12_5.C_ON=1'b0;
    defparam mux_129_Mux_3_i19_3_lut_LC_19_12_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i19_3_lut_LC_19_12_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_3_i19_3_lut_LC_19_12_5 (
            .in0(N__57812),
            .in1(N__50949),
            .in2(_gnd_net_),
            .in3(N__50922),
            .lcout(n19_adj_1515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_3_i26_3_lut_LC_19_12_6.C_ON=1'b0;
    defparam mux_129_Mux_3_i26_3_lut_LC_19_12_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i26_3_lut_LC_19_12_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_3_i26_3_lut_LC_19_12_6 (
            .in0(N__50883),
            .in1(N__57813),
            .in2(_gnd_net_),
            .in3(N__50861),
            .lcout(),
            .ltout(n26_adj_1516_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18523_4_lut_LC_19_12_7.C_ON=1'b0;
    defparam i18523_4_lut_LC_19_12_7.SEQ_MODE=4'b0000;
    defparam i18523_4_lut_LC_19_12_7.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18523_4_lut_LC_19_12_7 (
            .in0(N__57814),
            .in1(N__50835),
            .in2(N__50820),
            .in3(N__55141),
            .lcout(n21133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19098_4_lut_LC_19_13_0.C_ON=1'b0;
    defparam i19098_4_lut_LC_19_13_0.SEQ_MODE=4'b0000;
    defparam i19098_4_lut_LC_19_13_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 i19098_4_lut_LC_19_13_0 (
            .in0(N__57089),
            .in1(N__54653),
            .in2(N__52197),
            .in3(N__53794),
            .lcout(),
            .ltout(n21316_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i2_LC_19_13_1.C_ON=1'b0;
    defparam comm_length_i2_LC_19_13_1.SEQ_MODE=4'b1000;
    defparam comm_length_i2_LC_19_13_1.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_length_i2_LC_19_13_1 (
            .in0(N__53924),
            .in1(N__50808),
            .in2(N__50811),
            .in3(N__57754),
            .lcout(comm_length_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54404),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_315_LC_19_13_2.C_ON=1'b0;
    defparam i1_4_lut_adj_315_LC_19_13_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_315_LC_19_13_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_315_LC_19_13_2 (
            .in0(N__50807),
            .in1(N__50782),
            .in2(N__55248),
            .in3(N__50601),
            .lcout(n4_adj_1600),
            .ltout(n4_adj_1600_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_319_LC_19_13_3.C_ON=1'b0;
    defparam i2_3_lut_adj_319_LC_19_13_3.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_319_LC_19_13_3.LUT_INIT=16'b1111001111111100;
    LogicCell40 i2_3_lut_adj_319_LC_19_13_3 (
            .in0(_gnd_net_),
            .in1(N__54449),
            .in2(N__52416),
            .in3(N__52412),
            .lcout(),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19278_3_lut_LC_19_13_4.C_ON=1'b0;
    defparam i19278_3_lut_LC_19_13_4.SEQ_MODE=4'b0000;
    defparam i19278_3_lut_LC_19_13_4.LUT_INIT=16'b1100110011000000;
    LogicCell40 i19278_3_lut_LC_19_13_4 (
            .in0(_gnd_net_),
            .in1(N__52000),
            .in2(N__52269),
            .in3(N__52258),
            .lcout(n21888),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19194_2_lut_LC_19_13_5.C_ON=1'b0;
    defparam i19194_2_lut_LC_19_13_5.SEQ_MODE=4'b0000;
    defparam i19194_2_lut_LC_19_13_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 i19194_2_lut_LC_19_13_5 (
            .in0(N__55231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55421),
            .lcout(n21317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18438_3_lut_LC_19_13_6.C_ON=1'b0;
    defparam i18438_3_lut_LC_19_13_6.SEQ_MODE=4'b0000;
    defparam i18438_3_lut_LC_19_13_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18438_3_lut_LC_19_13_6 (
            .in0(N__52187),
            .in1(N__52146),
            .in2(_gnd_net_),
            .in3(N__55230),
            .lcout(n21048),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i5_LC_19_14_0.C_ON=1'b0;
    defparam comm_buf_1__i5_LC_19_14_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i5_LC_19_14_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i5_LC_19_14_0 (
            .in0(N__52124),
            .in1(N__52028),
            .in2(_gnd_net_),
            .in3(N__52794),
            .lcout(comm_buf_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54417),
            .ce(N__51382),
            .sr(N__51301));
    defparam comm_cmd_1__bdd_4_lut_19759_LC_19_14_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19759_LC_19_14_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19759_LC_19_14_2.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19759_LC_19_14_2 (
            .in0(N__51228),
            .in1(N__55218),
            .in2(N__51210),
            .in3(N__53782),
            .lcout(n22399),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i26_3_lut_LC_19_14_3.C_ON=1'b0;
    defparam mux_129_Mux_5_i26_3_lut_LC_19_14_3.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i26_3_lut_LC_19_14_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_5_i26_3_lut_LC_19_14_3 (
            .in0(N__51177),
            .in1(N__57750),
            .in2(_gnd_net_),
            .in3(N__51156),
            .lcout(),
            .ltout(n26_adj_1498_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19709_LC_19_14_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19709_LC_19_14_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19709_LC_19_14_4.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19709_LC_19_14_4 (
            .in0(N__57837),
            .in1(N__55219),
            .in2(N__51129),
            .in3(N__53783),
            .lcout(),
            .ltout(n22345_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22345_bdd_4_lut_LC_19_14_5.C_ON=1'b0;
    defparam n22345_bdd_4_lut_LC_19_14_5.SEQ_MODE=4'b0000;
    defparam n22345_bdd_4_lut_LC_19_14_5.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22345_bdd_4_lut_LC_19_14_5 (
            .in0(N__53784),
            .in1(N__52851),
            .in2(N__52824),
            .in3(N__52821),
            .lcout(),
            .ltout(n22348_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1556776_i1_3_lut_LC_19_14_6.C_ON=1'b0;
    defparam i1556776_i1_3_lut_LC_19_14_6.SEQ_MODE=4'b0000;
    defparam i1556776_i1_3_lut_LC_19_14_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1556776_i1_3_lut_LC_19_14_6 (
            .in0(_gnd_net_),
            .in1(N__53358),
            .in2(N__52797),
            .in3(N__54763),
            .lcout(n30_adj_1500),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18516_3_lut_LC_19_15_0.C_ON=1'b0;
    defparam i18516_3_lut_LC_19_15_0.SEQ_MODE=4'b0000;
    defparam i18516_3_lut_LC_19_15_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18516_3_lut_LC_19_15_0 (
            .in0(N__52787),
            .in1(N__52752),
            .in2(_gnd_net_),
            .in3(N__55232),
            .lcout(n21126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19322_2_lut_LC_19_17_3.C_ON=1'b0;
    defparam i19322_2_lut_LC_19_17_3.SEQ_MODE=4'b0000;
    defparam i19322_2_lut_LC_19_17_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19322_2_lut_LC_19_17_3 (
            .in0(_gnd_net_),
            .in1(N__52734),
            .in2(_gnd_net_),
            .in3(N__57749),
            .lcout(n21564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18970_2_lut_LC_19_18_2.C_ON=1'b0;
    defparam i18970_2_lut_LC_19_18_2.SEQ_MODE=4'b0000;
    defparam i18970_2_lut_LC_19_18_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18970_2_lut_LC_19_18_2 (
            .in0(_gnd_net_),
            .in1(N__52707),
            .in2(_gnd_net_),
            .in3(N__57748),
            .lcout(n21218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19053_2_lut_LC_20_3_2.C_ON=1'b0;
    defparam i19053_2_lut_LC_20_3_2.SEQ_MODE=4'b0000;
    defparam i19053_2_lut_LC_20_3_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 i19053_2_lut_LC_20_3_2 (
            .in0(N__52680),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57820),
            .lcout(n21364),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i1_LC_20_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i1_LC_20_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i1_LC_20_5_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ADC_VDC.genclk.div_state_i1_LC_20_5_4  (
            .in0(_gnd_net_),
            .in1(N__52906),
            .in2(_gnd_net_),
            .in3(N__58002),
            .lcout(\ADC_VDC.genclk.div_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i1C_net ),
            .ce(N__52650),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12196_12197_reset_LC_20_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12196_12197_reset_LC_20_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i0_12196_12197_reset_LC_20_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_12196_12197_reset_LC_20_6_0  (
            .in0(N__55901),
            .in1(N__52950),
            .in2(_gnd_net_),
            .in3(N__52970),
            .lcout(\comm_spi.n14615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52627),
            .ce(),
            .sr(N__53334));
    defparam \ADC_VDC.genclk.div_state_i0_LC_20_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i0_LC_20_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i0_LC_20_7_0 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \ADC_VDC.genclk.div_state_i0_LC_20_7_0  (
            .in0(N__58005),
            .in1(N__53352),
            .in2(N__58161),
            .in3(N__52894),
            .lcout(\ADC_VDC.genclk.div_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_20_7_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_20_7_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_87_2_lut_LC_20_7_1  (
            .in0(N__55765),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52875),
            .lcout(\comm_spi.DOUT_7__N_747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t_clk_24_LC_20_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t_clk_24_LC_20_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t_clk_24_LC_20_7_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ADC_VDC.genclk.t_clk_24_LC_20_7_2  (
            .in0(N__58004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(VDC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12198_3_lut_LC_20_7_3 .C_ON=1'b0;
    defparam \comm_spi.i12198_3_lut_LC_20_7_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12198_3_lut_LC_20_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i12198_3_lut_LC_20_7_3  (
            .in0(N__53067),
            .in1(N__53061),
            .in2(_gnd_net_),
            .in3(N__52862),
            .lcout(comm_rx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19420_4_lut_3_lut_LC_20_7_4 .C_ON=1'b0;
    defparam \comm_spi.i19420_4_lut_3_lut_LC_20_7_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19420_4_lut_3_lut_LC_20_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19420_4_lut_3_lut_LC_20_7_4  (
            .in0(N__55614),
            .in1(N__52969),
            .in2(_gnd_net_),
            .in3(N__55763),
            .lcout(\comm_spi.n22866 ),
            .ltout(\comm_spi.n22866_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12184_3_lut_LC_20_7_5 .C_ON=1'b0;
    defparam \comm_spi.i12184_3_lut_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12184_3_lut_LC_20_7_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.i12184_3_lut_LC_20_7_5  (
            .in0(_gnd_net_),
            .in1(N__55900),
            .in2(N__52953),
            .in3(N__52949),
            .lcout(\comm_spi.imosi ),
            .ltout(\comm_spi.imosi_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_20_7_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_20_7_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_20_7_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \comm_spi.RESET_I_0_86_2_lut_LC_20_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52923),
            .in3(N__55764),
            .lcout(\comm_spi.DOUT_7__N_746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12646_2_lut_2_lut_LC_20_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12646_2_lut_2_lut_LC_20_7_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12646_2_lut_2_lut_LC_20_7_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ADC_VDC.genclk.i12646_2_lut_2_lut_LC_20_7_7  (
            .in0(N__52893),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58003),
            .lcout(\ADC_VDC.genclk.n15051 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19435_4_lut_3_lut_LC_20_8_1 .C_ON=1'b0;
    defparam \comm_spi.i19435_4_lut_3_lut_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19435_4_lut_3_lut_LC_20_8_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.i19435_4_lut_3_lut_LC_20_8_1  (
            .in0(N__52863),
            .in1(N__55868),
            .in2(_gnd_net_),
            .in3(N__52874),
            .lcout(\comm_spi.n22863 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_12182_12183_set_LC_20_9_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12182_12183_set_LC_20_9_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imosi_44_12182_12183_set_LC_20_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_12182_12183_set_LC_20_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55636),
            .lcout(\comm_spi.n14600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54365),
            .ce(),
            .sr(N__55572));
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_20_10_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_20_10_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_88_2_lut_LC_20_10_3  (
            .in0(N__55867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55638),
            .lcout(\comm_spi.imosi_N_752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12237_3_lut_LC_20_11_5.C_ON=1'b0;
    defparam i12237_3_lut_LC_20_11_5.SEQ_MODE=4'b0000;
    defparam i12237_3_lut_LC_20_11_5.LUT_INIT=16'b1010101000100010;
    LogicCell40 i12237_3_lut_LC_20_11_5 (
            .in0(N__53917),
            .in1(N__55422),
            .in2(_gnd_net_),
            .in3(N__57000),
            .lcout(n14655),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i0_LC_20_12_0.C_ON=1'b0;
    defparam comm_length_i0_LC_20_12_0.SEQ_MODE=4'b1000;
    defparam comm_length_i0_LC_20_12_0.LUT_INIT=16'b0001010111000110;
    LogicCell40 comm_length_i0_LC_20_12_0 (
            .in0(N__54711),
            .in1(N__55235),
            .in2(N__57825),
            .in3(N__53614),
            .lcout(comm_length_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54405),
            .ce(N__53925),
            .sr(N__53901));
    defparam comm_length_i1_LC_20_12_1.C_ON=1'b0;
    defparam comm_length_i1_LC_20_12_1.SEQ_MODE=4'b1000;
    defparam comm_length_i1_LC_20_12_1.LUT_INIT=16'b1011111011001111;
    LogicCell40 comm_length_i1_LC_20_12_1 (
            .in0(N__53613),
            .in1(N__57808),
            .in2(N__55239),
            .in3(N__54712),
            .lcout(comm_length_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__54405),
            .ce(N__53925),
            .sr(N__53901));
    defparam i19319_2_lut_LC_20_13_0.C_ON=1'b0;
    defparam i19319_2_lut_LC_20_13_0.SEQ_MODE=4'b0000;
    defparam i19319_2_lut_LC_20_13_0.LUT_INIT=16'b1111101011111010;
    LogicCell40 i19319_2_lut_LC_20_13_0 (
            .in0(N__57779),
            .in1(_gnd_net_),
            .in2(N__53895),
            .in3(_gnd_net_),
            .lcout(n21451),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18978_2_lut_LC_20_13_3.C_ON=1'b0;
    defparam i18978_2_lut_LC_20_13_3.SEQ_MODE=4'b0000;
    defparam i18978_2_lut_LC_20_13_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 i18978_2_lut_LC_20_13_3 (
            .in0(_gnd_net_),
            .in1(N__53874),
            .in2(_gnd_net_),
            .in3(N__57778),
            .lcout(n21151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22399_bdd_4_lut_LC_20_14_0.C_ON=1'b0;
    defparam n22399_bdd_4_lut_LC_20_14_0.SEQ_MODE=4'b0000;
    defparam n22399_bdd_4_lut_LC_20_14_0.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22399_bdd_4_lut_LC_20_14_0 (
            .in0(N__53850),
            .in1(N__53838),
            .in2(N__53831),
            .in3(N__53785),
            .lcout(n22402),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19119_2_lut_LC_20_14_2.C_ON=1'b0;
    defparam i19119_2_lut_LC_20_14_2.SEQ_MODE=4'b0000;
    defparam i19119_2_lut_LC_20_14_2.LUT_INIT=16'b1111111110101010;
    LogicCell40 i19119_2_lut_LC_20_14_2 (
            .in0(N__57843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57780),
            .lcout(n21350),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19283_2_lut_LC_20_19_1.C_ON=1'b0;
    defparam i19283_2_lut_LC_20_19_1.SEQ_MODE=4'b0000;
    defparam i19283_2_lut_LC_20_19_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19283_2_lut_LC_20_19_1 (
            .in0(_gnd_net_),
            .in1(N__57831),
            .in2(_gnd_net_),
            .in3(N__57818),
            .lcout(n21529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15092_4_lut_LC_20_19_4.C_ON=1'b0;
    defparam i15092_4_lut_LC_20_19_4.SEQ_MODE=4'b0000;
    defparam i15092_4_lut_LC_20_19_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 i15092_4_lut_LC_20_19_4 (
            .in0(N__56999),
            .in1(N__56594),
            .in2(N__56518),
            .in3(N__56031),
            .lcout(data_index_9_N_216_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0on_i0_LC_22_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i0_LC_22_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i0_LC_22_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i0_LC_22_7_0  (
            .in0(_gnd_net_),
            .in1(N__58176),
            .in2(_gnd_net_),
            .in3(N__55917),
            .lcout(\ADC_VDC.genclk.t0on_0 ),
            .ltout(),
            .carryin(bfn_22_7_0_),
            .carryout(\ADC_VDC.genclk.n19724 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i1_LC_22_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i1_LC_22_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i1_LC_22_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i1_LC_22_7_1  (
            .in0(_gnd_net_),
            .in1(N__58206),
            .in2(N__58577),
            .in3(N__55914),
            .lcout(\ADC_VDC.genclk.t0on_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19724 ),
            .carryout(\ADC_VDC.genclk.n19725 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i2_LC_22_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i2_LC_22_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i2_LC_22_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i2_LC_22_7_2  (
            .in0(_gnd_net_),
            .in1(N__58545),
            .in2(N__58119),
            .in3(N__55911),
            .lcout(\ADC_VDC.genclk.t0on_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19725 ),
            .carryout(\ADC_VDC.genclk.n19726 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i3_LC_22_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i3_LC_22_7_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0on_i3_LC_22_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i3_LC_22_7_3  (
            .in0(_gnd_net_),
            .in1(N__58071),
            .in2(N__58578),
            .in3(N__55908),
            .lcout(\ADC_VDC.genclk.t0on_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19726 ),
            .carryout(\ADC_VDC.genclk.n19727 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i4_LC_22_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i4_LC_22_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i4_LC_22_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i4_LC_22_7_4  (
            .in0(_gnd_net_),
            .in1(N__58549),
            .in2(N__58194),
            .in3(N__55905),
            .lcout(\ADC_VDC.genclk.t0on_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19727 ),
            .carryout(\ADC_VDC.genclk.n19728 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i5_LC_22_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i5_LC_22_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i5_LC_22_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i5_LC_22_7_5  (
            .in0(_gnd_net_),
            .in1(N__58043),
            .in2(N__58579),
            .in3(N__57870),
            .lcout(\ADC_VDC.genclk.t0on_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19728 ),
            .carryout(\ADC_VDC.genclk.n19729 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i6_LC_22_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i6_LC_22_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i6_LC_22_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i6_LC_22_7_6  (
            .in0(_gnd_net_),
            .in1(N__58553),
            .in2(N__58221),
            .in3(N__57867),
            .lcout(\ADC_VDC.genclk.t0on_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19729 ),
            .carryout(\ADC_VDC.genclk.n19730 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i7_LC_22_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i7_LC_22_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i7_LC_22_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i7_LC_22_7_7  (
            .in0(_gnd_net_),
            .in1(N__58103),
            .in2(N__58580),
            .in3(N__57864),
            .lcout(\ADC_VDC.genclk.t0on_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19730 ),
            .carryout(\ADC_VDC.genclk.n19731 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57959),
            .sr(N__58259));
    defparam \ADC_VDC.genclk.t0on_i8_LC_22_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i8_LC_22_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i8_LC_22_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i8_LC_22_8_0  (
            .in0(_gnd_net_),
            .in1(N__58029),
            .in2(N__58503),
            .in3(N__57861),
            .lcout(\ADC_VDC.genclk.t0on_8 ),
            .ltout(),
            .carryin(bfn_22_8_0_),
            .carryout(\ADC_VDC.genclk.n19732 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.t0on_i9_LC_22_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i9_LC_22_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i9_LC_22_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i9_LC_22_8_1  (
            .in0(_gnd_net_),
            .in1(N__58420),
            .in2(N__57924),
            .in3(N__57858),
            .lcout(\ADC_VDC.genclk.t0on_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19732 ),
            .carryout(\ADC_VDC.genclk.n19733 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.t0on_i10_LC_22_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i10_LC_22_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i10_LC_22_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i10_LC_22_8_2  (
            .in0(_gnd_net_),
            .in1(N__58089),
            .in2(N__58500),
            .in3(N__57855),
            .lcout(\ADC_VDC.genclk.t0on_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19733 ),
            .carryout(\ADC_VDC.genclk.n19734 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.t0on_i11_LC_22_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i11_LC_22_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i11_LC_22_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i11_LC_22_8_3  (
            .in0(_gnd_net_),
            .in1(N__58408),
            .in2(N__57894),
            .in3(N__57852),
            .lcout(\ADC_VDC.genclk.t0on_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19734 ),
            .carryout(\ADC_VDC.genclk.n19735 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.t0on_i12_LC_22_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i12_LC_22_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i12_LC_22_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i12_LC_22_8_4  (
            .in0(_gnd_net_),
            .in1(N__58131),
            .in2(N__58501),
            .in3(N__57849),
            .lcout(\ADC_VDC.genclk.t0on_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19735 ),
            .carryout(\ADC_VDC.genclk.n19736 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.t0on_i13_LC_22_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i13_LC_22_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i13_LC_22_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i13_LC_22_8_5  (
            .in0(_gnd_net_),
            .in1(N__58412),
            .in2(N__58059),
            .in3(N__57846),
            .lcout(\ADC_VDC.genclk.t0on_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19736 ),
            .carryout(\ADC_VDC.genclk.n19737 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.t0on_i14_LC_22_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i14_LC_22_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i14_LC_22_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i14_LC_22_8_6  (
            .in0(_gnd_net_),
            .in1(N__57936),
            .in2(N__58502),
            .in3(N__58626),
            .lcout(\ADC_VDC.genclk.t0on_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19737 ),
            .carryout(\ADC_VDC.genclk.n19738 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.t0on_i15_LC_22_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0on_i15_LC_22_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i15_LC_22_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0on_i15_LC_22_8_7  (
            .in0(N__57908),
            .in1(N__58416),
            .in2(_gnd_net_),
            .in3(N__58266),
            .lcout(\ADC_VDC.genclk.t0on_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57963),
            .sr(N__58258));
    defparam \ADC_VDC.genclk.i19049_4_lut_LC_23_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19049_4_lut_LC_23_7_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19049_4_lut_LC_23_7_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i19049_4_lut_LC_23_7_0  (
            .in0(N__58217),
            .in1(N__58205),
            .in2(N__58193),
            .in3(N__58175),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n21449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19183_4_lut_LC_23_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19183_4_lut_LC_23_7_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19183_4_lut_LC_23_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i19183_4_lut_LC_23_7_1  (
            .in0(N__57879),
            .in1(N__58017),
            .in2(N__58164),
            .in3(N__58077),
            .lcout(\ADC_VDC.genclk.n21443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_adj_7_LC_23_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_7_LC_23_7_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_7_LC_23_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_adj_7_LC_23_7_2  (
            .in0(N__58130),
            .in1(N__58115),
            .in2(N__58104),
            .in3(N__58088),
            .lcout(\ADC_VDC.genclk.n27_adj_1396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_adj_6_LC_23_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_6_LC_23_7_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_6_LC_23_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_adj_6_LC_23_7_3  (
            .in0(N__58070),
            .in1(N__58055),
            .in2(N__58044),
            .in3(N__58028),
            .lcout(\ADC_VDC.genclk.n26_adj_1395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_23_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_23_7_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_23_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_23_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58011),
            .lcout(\ADC_VDC.genclk.div_state_1__N_1274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_LC_23_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_23_8_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_23_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_LC_23_8_3  (
            .in0(N__57935),
            .in1(N__57920),
            .in2(N__57909),
            .in3(N__57890),
            .lcout(\ADC_VDC.genclk.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // zim
