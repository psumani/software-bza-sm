// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 1 2024 11:48:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "zimaux" view "INTERFACE"

module zimaux (
    M_CS1,
    ICE_SYSCLK,
    M_MOSI1,
    M_DRDY1,
    M_CLK2,
    M_SCLK1,
    M_FLT0,
    M_CS3,
    ICE_CHKCABLE,
    M_OSR1,
    ICE_GPMO_1,
    EIS_SYNCCLK,
    M_SCLK3,
    M_OSR0,
    M_MISO4,
    M_DRDY4,
    ICE_SPI_MOSI,
    ICE_GPMO_0,
    DDS_MOSI1,
    M_SCLK4,
    M_MISO3,
    M_CS4,
    ICE_SPI_SCLK,
    M_MOSI4,
    M_MISO2,
    M_DRDY2,
    M_CLK1,
    ICE_SPI_MISO,
    ICE_GPMO_2,
    ICE_GPMI_0,
    TEST_LED,
    M_POW,
    M_MOSI3,
    M_MISO1,
    M_DRDY3,
    M_DCSEL,
    M_START,
    M_MOSI2,
    M_CLK3,
    DDS_CS1,
    M_FLT1,
    DISP_COMM,
    DDS_MCLK1,
    ICE_SPI_CE0,
    M_SCLK2,
    M_CS2,
    M_CLK4,
    DDS_SCK1);

    output M_CS1;
    input ICE_SYSCLK;
    output M_MOSI1;
    input M_DRDY1;
    output M_CLK2;
    output M_SCLK1;
    output M_FLT0;
    output M_CS3;
    input ICE_CHKCABLE;
    output M_OSR1;
    input ICE_GPMO_1;
    input EIS_SYNCCLK;
    output M_SCLK3;
    output M_OSR0;
    input M_MISO4;
    input M_DRDY4;
    input ICE_SPI_MOSI;
    input ICE_GPMO_0;
    output DDS_MOSI1;
    output M_SCLK4;
    input M_MISO3;
    output M_CS4;
    input ICE_SPI_SCLK;
    output M_MOSI4;
    input M_MISO2;
    input M_DRDY2;
    output M_CLK1;
    output ICE_SPI_MISO;
    input ICE_GPMO_2;
    output ICE_GPMI_0;
    output TEST_LED;
    output M_POW;
    output M_MOSI3;
    input M_MISO1;
    input M_DRDY3;
    output M_DCSEL;
    output M_START;
    output M_MOSI2;
    output M_CLK3;
    output DDS_CS1;
    output M_FLT1;
    output DISP_COMM;
    output DDS_MCLK1;
    input ICE_SPI_CE0;
    output M_SCLK2;
    output M_CS2;
    output M_CLK4;
    output DDS_SCK1;

    wire N__54255;
    wire N__54254;
    wire N__54253;
    wire N__54246;
    wire N__54245;
    wire N__54244;
    wire N__54237;
    wire N__54236;
    wire N__54235;
    wire N__54228;
    wire N__54227;
    wire N__54226;
    wire N__54219;
    wire N__54218;
    wire N__54217;
    wire N__54210;
    wire N__54209;
    wire N__54208;
    wire N__54201;
    wire N__54200;
    wire N__54199;
    wire N__54192;
    wire N__54191;
    wire N__54190;
    wire N__54183;
    wire N__54182;
    wire N__54181;
    wire N__54174;
    wire N__54173;
    wire N__54172;
    wire N__54165;
    wire N__54164;
    wire N__54163;
    wire N__54156;
    wire N__54155;
    wire N__54154;
    wire N__54147;
    wire N__54146;
    wire N__54145;
    wire N__54138;
    wire N__54137;
    wire N__54136;
    wire N__54129;
    wire N__54128;
    wire N__54127;
    wire N__54120;
    wire N__54119;
    wire N__54118;
    wire N__54111;
    wire N__54110;
    wire N__54109;
    wire N__54102;
    wire N__54101;
    wire N__54100;
    wire N__54093;
    wire N__54092;
    wire N__54091;
    wire N__54084;
    wire N__54083;
    wire N__54082;
    wire N__54075;
    wire N__54074;
    wire N__54073;
    wire N__54066;
    wire N__54065;
    wire N__54064;
    wire N__54057;
    wire N__54056;
    wire N__54055;
    wire N__54048;
    wire N__54047;
    wire N__54046;
    wire N__54039;
    wire N__54038;
    wire N__54037;
    wire N__54030;
    wire N__54029;
    wire N__54028;
    wire N__54021;
    wire N__54020;
    wire N__54019;
    wire N__54012;
    wire N__54011;
    wire N__54010;
    wire N__54003;
    wire N__54002;
    wire N__54001;
    wire N__53994;
    wire N__53993;
    wire N__53992;
    wire N__53985;
    wire N__53984;
    wire N__53983;
    wire N__53976;
    wire N__53975;
    wire N__53974;
    wire N__53967;
    wire N__53966;
    wire N__53965;
    wire N__53958;
    wire N__53957;
    wire N__53956;
    wire N__53949;
    wire N__53948;
    wire N__53947;
    wire N__53940;
    wire N__53939;
    wire N__53938;
    wire N__53931;
    wire N__53930;
    wire N__53929;
    wire N__53922;
    wire N__53921;
    wire N__53920;
    wire N__53913;
    wire N__53912;
    wire N__53911;
    wire N__53904;
    wire N__53903;
    wire N__53902;
    wire N__53895;
    wire N__53894;
    wire N__53893;
    wire N__53886;
    wire N__53885;
    wire N__53884;
    wire N__53877;
    wire N__53876;
    wire N__53875;
    wire N__53868;
    wire N__53867;
    wire N__53866;
    wire N__53859;
    wire N__53858;
    wire N__53857;
    wire N__53850;
    wire N__53849;
    wire N__53848;
    wire N__53841;
    wire N__53840;
    wire N__53839;
    wire N__53832;
    wire N__53831;
    wire N__53830;
    wire N__53813;
    wire N__53812;
    wire N__53811;
    wire N__53810;
    wire N__53809;
    wire N__53806;
    wire N__53803;
    wire N__53800;
    wire N__53799;
    wire N__53798;
    wire N__53795;
    wire N__53792;
    wire N__53785;
    wire N__53782;
    wire N__53779;
    wire N__53776;
    wire N__53775;
    wire N__53774;
    wire N__53771;
    wire N__53766;
    wire N__53761;
    wire N__53758;
    wire N__53755;
    wire N__53754;
    wire N__53753;
    wire N__53752;
    wire N__53751;
    wire N__53740;
    wire N__53735;
    wire N__53734;
    wire N__53733;
    wire N__53730;
    wire N__53727;
    wire N__53722;
    wire N__53717;
    wire N__53716;
    wire N__53713;
    wire N__53710;
    wire N__53705;
    wire N__53704;
    wire N__53703;
    wire N__53702;
    wire N__53699;
    wire N__53698;
    wire N__53697;
    wire N__53696;
    wire N__53695;
    wire N__53692;
    wire N__53689;
    wire N__53686;
    wire N__53685;
    wire N__53678;
    wire N__53675;
    wire N__53672;
    wire N__53669;
    wire N__53664;
    wire N__53661;
    wire N__53656;
    wire N__53653;
    wire N__53650;
    wire N__53647;
    wire N__53642;
    wire N__53639;
    wire N__53636;
    wire N__53633;
    wire N__53626;
    wire N__53619;
    wire N__53616;
    wire N__53609;
    wire N__53606;
    wire N__53605;
    wire N__53602;
    wire N__53599;
    wire N__53596;
    wire N__53593;
    wire N__53592;
    wire N__53589;
    wire N__53586;
    wire N__53583;
    wire N__53576;
    wire N__53575;
    wire N__53574;
    wire N__53573;
    wire N__53572;
    wire N__53571;
    wire N__53570;
    wire N__53569;
    wire N__53566;
    wire N__53561;
    wire N__53552;
    wire N__53549;
    wire N__53546;
    wire N__53543;
    wire N__53540;
    wire N__53539;
    wire N__53538;
    wire N__53537;
    wire N__53536;
    wire N__53535;
    wire N__53534;
    wire N__53533;
    wire N__53532;
    wire N__53531;
    wire N__53528;
    wire N__53527;
    wire N__53526;
    wire N__53525;
    wire N__53524;
    wire N__53523;
    wire N__53522;
    wire N__53521;
    wire N__53520;
    wire N__53519;
    wire N__53518;
    wire N__53517;
    wire N__53516;
    wire N__53515;
    wire N__53510;
    wire N__53507;
    wire N__53494;
    wire N__53493;
    wire N__53492;
    wire N__53489;
    wire N__53484;
    wire N__53483;
    wire N__53482;
    wire N__53481;
    wire N__53478;
    wire N__53475;
    wire N__53474;
    wire N__53471;
    wire N__53468;
    wire N__53457;
    wire N__53446;
    wire N__53439;
    wire N__53438;
    wire N__53437;
    wire N__53436;
    wire N__53435;
    wire N__53434;
    wire N__53433;
    wire N__53430;
    wire N__53427;
    wire N__53422;
    wire N__53417;
    wire N__53414;
    wire N__53409;
    wire N__53408;
    wire N__53407;
    wire N__53406;
    wire N__53405;
    wire N__53404;
    wire N__53403;
    wire N__53402;
    wire N__53399;
    wire N__53394;
    wire N__53393;
    wire N__53392;
    wire N__53391;
    wire N__53390;
    wire N__53385;
    wire N__53382;
    wire N__53379;
    wire N__53370;
    wire N__53367;
    wire N__53362;
    wire N__53357;
    wire N__53356;
    wire N__53355;
    wire N__53354;
    wire N__53349;
    wire N__53336;
    wire N__53335;
    wire N__53332;
    wire N__53329;
    wire N__53326;
    wire N__53325;
    wire N__53316;
    wire N__53313;
    wire N__53310;
    wire N__53307;
    wire N__53304;
    wire N__53301;
    wire N__53298;
    wire N__53295;
    wire N__53294;
    wire N__53293;
    wire N__53290;
    wire N__53285;
    wire N__53282;
    wire N__53279;
    wire N__53278;
    wire N__53277;
    wire N__53276;
    wire N__53275;
    wire N__53272;
    wire N__53269;
    wire N__53264;
    wire N__53261;
    wire N__53258;
    wire N__53253;
    wire N__53248;
    wire N__53243;
    wire N__53240;
    wire N__53237;
    wire N__53234;
    wire N__53229;
    wire N__53224;
    wire N__53223;
    wire N__53222;
    wire N__53221;
    wire N__53220;
    wire N__53219;
    wire N__53216;
    wire N__53213;
    wire N__53210;
    wire N__53207;
    wire N__53204;
    wire N__53199;
    wire N__53192;
    wire N__53185;
    wire N__53176;
    wire N__53165;
    wire N__53144;
    wire N__53143;
    wire N__53140;
    wire N__53137;
    wire N__53134;
    wire N__53129;
    wire N__53128;
    wire N__53127;
    wire N__53126;
    wire N__53125;
    wire N__53124;
    wire N__53123;
    wire N__53118;
    wire N__53117;
    wire N__53116;
    wire N__53115;
    wire N__53114;
    wire N__53107;
    wire N__53102;
    wire N__53101;
    wire N__53098;
    wire N__53095;
    wire N__53092;
    wire N__53089;
    wire N__53086;
    wire N__53085;
    wire N__53084;
    wire N__53079;
    wire N__53078;
    wire N__53077;
    wire N__53076;
    wire N__53075;
    wire N__53072;
    wire N__53065;
    wire N__53064;
    wire N__53063;
    wire N__53060;
    wire N__53057;
    wire N__53052;
    wire N__53051;
    wire N__53050;
    wire N__53049;
    wire N__53046;
    wire N__53037;
    wire N__53034;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53022;
    wire N__53019;
    wire N__53016;
    wire N__53015;
    wire N__53012;
    wire N__53009;
    wire N__53006;
    wire N__53001;
    wire N__52998;
    wire N__52995;
    wire N__52990;
    wire N__52987;
    wire N__52984;
    wire N__52981;
    wire N__52978;
    wire N__52969;
    wire N__52966;
    wire N__52963;
    wire N__52956;
    wire N__52953;
    wire N__52944;
    wire N__52941;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52925;
    wire N__52922;
    wire N__52921;
    wire N__52918;
    wire N__52917;
    wire N__52914;
    wire N__52911;
    wire N__52908;
    wire N__52905;
    wire N__52898;
    wire N__52897;
    wire N__52896;
    wire N__52895;
    wire N__52894;
    wire N__52893;
    wire N__52892;
    wire N__52891;
    wire N__52890;
    wire N__52889;
    wire N__52888;
    wire N__52885;
    wire N__52884;
    wire N__52883;
    wire N__52882;
    wire N__52881;
    wire N__52880;
    wire N__52879;
    wire N__52878;
    wire N__52877;
    wire N__52876;
    wire N__52875;
    wire N__52874;
    wire N__52871;
    wire N__52868;
    wire N__52863;
    wire N__52860;
    wire N__52857;
    wire N__52854;
    wire N__52853;
    wire N__52852;
    wire N__52851;
    wire N__52850;
    wire N__52849;
    wire N__52848;
    wire N__52847;
    wire N__52846;
    wire N__52845;
    wire N__52844;
    wire N__52841;
    wire N__52838;
    wire N__52837;
    wire N__52836;
    wire N__52835;
    wire N__52834;
    wire N__52833;
    wire N__52832;
    wire N__52831;
    wire N__52814;
    wire N__52813;
    wire N__52810;
    wire N__52809;
    wire N__52806;
    wire N__52799;
    wire N__52798;
    wire N__52797;
    wire N__52796;
    wire N__52795;
    wire N__52794;
    wire N__52793;
    wire N__52790;
    wire N__52785;
    wire N__52782;
    wire N__52779;
    wire N__52778;
    wire N__52775;
    wire N__52774;
    wire N__52763;
    wire N__52760;
    wire N__52757;
    wire N__52754;
    wire N__52751;
    wire N__52748;
    wire N__52745;
    wire N__52742;
    wire N__52739;
    wire N__52736;
    wire N__52725;
    wire N__52722;
    wire N__52719;
    wire N__52714;
    wire N__52711;
    wire N__52708;
    wire N__52699;
    wire N__52696;
    wire N__52693;
    wire N__52690;
    wire N__52683;
    wire N__52680;
    wire N__52679;
    wire N__52678;
    wire N__52677;
    wire N__52676;
    wire N__52675;
    wire N__52674;
    wire N__52673;
    wire N__52672;
    wire N__52671;
    wire N__52670;
    wire N__52667;
    wire N__52664;
    wire N__52659;
    wire N__52656;
    wire N__52653;
    wire N__52650;
    wire N__52645;
    wire N__52636;
    wire N__52631;
    wire N__52628;
    wire N__52621;
    wire N__52620;
    wire N__52619;
    wire N__52618;
    wire N__52617;
    wire N__52616;
    wire N__52607;
    wire N__52606;
    wire N__52605;
    wire N__52604;
    wire N__52603;
    wire N__52598;
    wire N__52595;
    wire N__52578;
    wire N__52571;
    wire N__52564;
    wire N__52559;
    wire N__52552;
    wire N__52545;
    wire N__52540;
    wire N__52537;
    wire N__52528;
    wire N__52505;
    wire N__52504;
    wire N__52501;
    wire N__52498;
    wire N__52495;
    wire N__52490;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52469;
    wire N__52468;
    wire N__52467;
    wire N__52466;
    wire N__52463;
    wire N__52462;
    wire N__52461;
    wire N__52460;
    wire N__52459;
    wire N__52458;
    wire N__52457;
    wire N__52456;
    wire N__52455;
    wire N__52454;
    wire N__52453;
    wire N__52452;
    wire N__52451;
    wire N__52450;
    wire N__52449;
    wire N__52448;
    wire N__52447;
    wire N__52446;
    wire N__52445;
    wire N__52444;
    wire N__52443;
    wire N__52442;
    wire N__52439;
    wire N__52436;
    wire N__52435;
    wire N__52434;
    wire N__52433;
    wire N__52432;
    wire N__52431;
    wire N__52430;
    wire N__52427;
    wire N__52426;
    wire N__52425;
    wire N__52424;
    wire N__52423;
    wire N__52420;
    wire N__52419;
    wire N__52418;
    wire N__52415;
    wire N__52414;
    wire N__52411;
    wire N__52410;
    wire N__52407;
    wire N__52406;
    wire N__52403;
    wire N__52402;
    wire N__52399;
    wire N__52398;
    wire N__52395;
    wire N__52394;
    wire N__52391;
    wire N__52390;
    wire N__52387;
    wire N__52386;
    wire N__52385;
    wire N__52384;
    wire N__52381;
    wire N__52380;
    wire N__52377;
    wire N__52376;
    wire N__52369;
    wire N__52364;
    wire N__52361;
    wire N__52360;
    wire N__52357;
    wire N__52356;
    wire N__52351;
    wire N__52350;
    wire N__52349;
    wire N__52346;
    wire N__52345;
    wire N__52342;
    wire N__52337;
    wire N__52332;
    wire N__52327;
    wire N__52322;
    wire N__52319;
    wire N__52314;
    wire N__52313;
    wire N__52312;
    wire N__52311;
    wire N__52310;
    wire N__52309;
    wire N__52306;
    wire N__52303;
    wire N__52302;
    wire N__52301;
    wire N__52300;
    wire N__52297;
    wire N__52280;
    wire N__52265;
    wire N__52262;
    wire N__52259;
    wire N__52254;
    wire N__52247;
    wire N__52244;
    wire N__52241;
    wire N__52240;
    wire N__52239;
    wire N__52238;
    wire N__52233;
    wire N__52230;
    wire N__52225;
    wire N__52222;
    wire N__52221;
    wire N__52220;
    wire N__52219;
    wire N__52218;
    wire N__52217;
    wire N__52214;
    wire N__52211;
    wire N__52208;
    wire N__52205;
    wire N__52202;
    wire N__52187;
    wire N__52186;
    wire N__52185;
    wire N__52184;
    wire N__52183;
    wire N__52172;
    wire N__52169;
    wire N__52166;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52156;
    wire N__52149;
    wire N__52146;
    wire N__52143;
    wire N__52140;
    wire N__52133;
    wire N__52126;
    wire N__52119;
    wire N__52110;
    wire N__52105;
    wire N__52102;
    wire N__52091;
    wire N__52086;
    wire N__52083;
    wire N__52082;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52074;
    wire N__52073;
    wire N__52070;
    wire N__52067;
    wire N__52066;
    wire N__52063;
    wire N__52062;
    wire N__52061;
    wire N__52058;
    wire N__52051;
    wire N__52046;
    wire N__52039;
    wire N__52034;
    wire N__52033;
    wire N__52032;
    wire N__52025;
    wire N__52022;
    wire N__52019;
    wire N__52016;
    wire N__52013;
    wire N__52010;
    wire N__52007;
    wire N__52004;
    wire N__52001;
    wire N__51996;
    wire N__51991;
    wire N__51986;
    wire N__51977;
    wire N__51974;
    wire N__51969;
    wire N__51964;
    wire N__51953;
    wire N__51932;
    wire N__51931;
    wire N__51930;
    wire N__51929;
    wire N__51928;
    wire N__51927;
    wire N__51924;
    wire N__51923;
    wire N__51922;
    wire N__51919;
    wire N__51918;
    wire N__51917;
    wire N__51916;
    wire N__51915;
    wire N__51914;
    wire N__51913;
    wire N__51910;
    wire N__51909;
    wire N__51906;
    wire N__51903;
    wire N__51900;
    wire N__51899;
    wire N__51898;
    wire N__51897;
    wire N__51896;
    wire N__51895;
    wire N__51894;
    wire N__51893;
    wire N__51890;
    wire N__51887;
    wire N__51884;
    wire N__51881;
    wire N__51880;
    wire N__51879;
    wire N__51876;
    wire N__51873;
    wire N__51870;
    wire N__51869;
    wire N__51868;
    wire N__51867;
    wire N__51866;
    wire N__51863;
    wire N__51860;
    wire N__51857;
    wire N__51854;
    wire N__51853;
    wire N__51852;
    wire N__51851;
    wire N__51848;
    wire N__51845;
    wire N__51844;
    wire N__51843;
    wire N__51842;
    wire N__51841;
    wire N__51838;
    wire N__51835;
    wire N__51830;
    wire N__51829;
    wire N__51826;
    wire N__51825;
    wire N__51822;
    wire N__51817;
    wire N__51814;
    wire N__51811;
    wire N__51808;
    wire N__51805;
    wire N__51802;
    wire N__51797;
    wire N__51794;
    wire N__51787;
    wire N__51784;
    wire N__51779;
    wire N__51776;
    wire N__51771;
    wire N__51770;
    wire N__51769;
    wire N__51768;
    wire N__51767;
    wire N__51766;
    wire N__51763;
    wire N__51758;
    wire N__51753;
    wire N__51750;
    wire N__51749;
    wire N__51746;
    wire N__51743;
    wire N__51740;
    wire N__51739;
    wire N__51738;
    wire N__51737;
    wire N__51734;
    wire N__51731;
    wire N__51726;
    wire N__51725;
    wire N__51722;
    wire N__51719;
    wire N__51716;
    wire N__51711;
    wire N__51708;
    wire N__51705;
    wire N__51700;
    wire N__51683;
    wire N__51680;
    wire N__51679;
    wire N__51676;
    wire N__51675;
    wire N__51672;
    wire N__51669;
    wire N__51668;
    wire N__51665;
    wire N__51664;
    wire N__51663;
    wire N__51658;
    wire N__51655;
    wire N__51652;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51636;
    wire N__51633;
    wire N__51630;
    wire N__51625;
    wire N__51620;
    wire N__51617;
    wire N__51614;
    wire N__51607;
    wire N__51602;
    wire N__51599;
    wire N__51594;
    wire N__51583;
    wire N__51578;
    wire N__51569;
    wire N__51566;
    wire N__51561;
    wire N__51558;
    wire N__51555;
    wire N__51550;
    wire N__51541;
    wire N__51530;
    wire N__51515;
    wire N__51512;
    wire N__51509;
    wire N__51508;
    wire N__51505;
    wire N__51502;
    wire N__51499;
    wire N__51494;
    wire N__51491;
    wire N__51488;
    wire N__51485;
    wire N__51482;
    wire N__51479;
    wire N__51476;
    wire N__51473;
    wire N__51470;
    wire N__51467;
    wire N__51464;
    wire N__51461;
    wire N__51460;
    wire N__51457;
    wire N__51454;
    wire N__51451;
    wire N__51448;
    wire N__51445;
    wire N__51442;
    wire N__51439;
    wire N__51436;
    wire N__51433;
    wire N__51430;
    wire N__51427;
    wire N__51424;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51404;
    wire N__51401;
    wire N__51398;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51390;
    wire N__51385;
    wire N__51382;
    wire N__51379;
    wire N__51376;
    wire N__51375;
    wire N__51374;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51354;
    wire N__51351;
    wire N__51346;
    wire N__51343;
    wire N__51340;
    wire N__51335;
    wire N__51332;
    wire N__51329;
    wire N__51326;
    wire N__51323;
    wire N__51320;
    wire N__51319;
    wire N__51318;
    wire N__51317;
    wire N__51316;
    wire N__51315;
    wire N__51314;
    wire N__51313;
    wire N__51312;
    wire N__51311;
    wire N__51310;
    wire N__51309;
    wire N__51308;
    wire N__51307;
    wire N__51306;
    wire N__51305;
    wire N__51304;
    wire N__51303;
    wire N__51302;
    wire N__51301;
    wire N__51300;
    wire N__51299;
    wire N__51298;
    wire N__51297;
    wire N__51296;
    wire N__51295;
    wire N__51294;
    wire N__51293;
    wire N__51292;
    wire N__51291;
    wire N__51290;
    wire N__51289;
    wire N__51288;
    wire N__51287;
    wire N__51286;
    wire N__51285;
    wire N__51284;
    wire N__51283;
    wire N__51282;
    wire N__51281;
    wire N__51280;
    wire N__51279;
    wire N__51278;
    wire N__51277;
    wire N__51276;
    wire N__51275;
    wire N__51274;
    wire N__51273;
    wire N__51272;
    wire N__51271;
    wire N__51270;
    wire N__51269;
    wire N__51268;
    wire N__51267;
    wire N__51266;
    wire N__51265;
    wire N__51264;
    wire N__51263;
    wire N__51262;
    wire N__51261;
    wire N__51260;
    wire N__51259;
    wire N__51258;
    wire N__51257;
    wire N__51256;
    wire N__51255;
    wire N__51254;
    wire N__51253;
    wire N__51252;
    wire N__51251;
    wire N__51250;
    wire N__51249;
    wire N__51248;
    wire N__51247;
    wire N__51246;
    wire N__51245;
    wire N__51244;
    wire N__51243;
    wire N__51242;
    wire N__51241;
    wire N__51240;
    wire N__51239;
    wire N__51238;
    wire N__51237;
    wire N__51236;
    wire N__51235;
    wire N__51234;
    wire N__51233;
    wire N__51232;
    wire N__51231;
    wire N__51230;
    wire N__51229;
    wire N__51228;
    wire N__51227;
    wire N__51226;
    wire N__51225;
    wire N__51224;
    wire N__51223;
    wire N__51222;
    wire N__51221;
    wire N__51220;
    wire N__51219;
    wire N__51218;
    wire N__51217;
    wire N__51216;
    wire N__51215;
    wire N__51214;
    wire N__51213;
    wire N__51212;
    wire N__51211;
    wire N__51210;
    wire N__51209;
    wire N__51208;
    wire N__51207;
    wire N__51206;
    wire N__51205;
    wire N__51204;
    wire N__51203;
    wire N__51202;
    wire N__51201;
    wire N__51200;
    wire N__51199;
    wire N__51198;
    wire N__51197;
    wire N__51196;
    wire N__51195;
    wire N__51194;
    wire N__51193;
    wire N__51192;
    wire N__51191;
    wire N__51190;
    wire N__51189;
    wire N__51188;
    wire N__51187;
    wire N__51186;
    wire N__51185;
    wire N__51184;
    wire N__51183;
    wire N__51182;
    wire N__51181;
    wire N__51180;
    wire N__51179;
    wire N__51178;
    wire N__51177;
    wire N__51176;
    wire N__51175;
    wire N__51174;
    wire N__51173;
    wire N__51172;
    wire N__51171;
    wire N__51170;
    wire N__51169;
    wire N__51168;
    wire N__51167;
    wire N__51166;
    wire N__51165;
    wire N__51164;
    wire N__51163;
    wire N__51162;
    wire N__51161;
    wire N__51160;
    wire N__51159;
    wire N__51158;
    wire N__51157;
    wire N__51156;
    wire N__51155;
    wire N__51154;
    wire N__51153;
    wire N__51152;
    wire N__51151;
    wire N__51150;
    wire N__51149;
    wire N__51148;
    wire N__51147;
    wire N__51146;
    wire N__51145;
    wire N__51144;
    wire N__51143;
    wire N__51142;
    wire N__51141;
    wire N__51140;
    wire N__51139;
    wire N__51138;
    wire N__51137;
    wire N__51136;
    wire N__51135;
    wire N__51134;
    wire N__51133;
    wire N__51132;
    wire N__51131;
    wire N__51130;
    wire N__51129;
    wire N__51128;
    wire N__51127;
    wire N__51126;
    wire N__51125;
    wire N__51124;
    wire N__51123;
    wire N__51122;
    wire N__51121;
    wire N__51120;
    wire N__51119;
    wire N__51118;
    wire N__51117;
    wire N__51116;
    wire N__51115;
    wire N__51114;
    wire N__51113;
    wire N__51112;
    wire N__51111;
    wire N__51110;
    wire N__51109;
    wire N__51108;
    wire N__51107;
    wire N__51106;
    wire N__50675;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50657;
    wire N__50656;
    wire N__50653;
    wire N__50650;
    wire N__50647;
    wire N__50644;
    wire N__50641;
    wire N__50638;
    wire N__50633;
    wire N__50630;
    wire N__50627;
    wire N__50624;
    wire N__50621;
    wire N__50618;
    wire N__50615;
    wire N__50612;
    wire N__50609;
    wire N__50606;
    wire N__50605;
    wire N__50604;
    wire N__50603;
    wire N__50602;
    wire N__50601;
    wire N__50600;
    wire N__50599;
    wire N__50598;
    wire N__50597;
    wire N__50596;
    wire N__50595;
    wire N__50594;
    wire N__50593;
    wire N__50590;
    wire N__50583;
    wire N__50582;
    wire N__50581;
    wire N__50580;
    wire N__50575;
    wire N__50570;
    wire N__50565;
    wire N__50562;
    wire N__50561;
    wire N__50560;
    wire N__50559;
    wire N__50558;
    wire N__50555;
    wire N__50554;
    wire N__50553;
    wire N__50552;
    wire N__50551;
    wire N__50550;
    wire N__50547;
    wire N__50544;
    wire N__50541;
    wire N__50538;
    wire N__50537;
    wire N__50536;
    wire N__50533;
    wire N__50528;
    wire N__50525;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50513;
    wire N__50512;
    wire N__50511;
    wire N__50510;
    wire N__50509;
    wire N__50508;
    wire N__50507;
    wire N__50506;
    wire N__50505;
    wire N__50504;
    wire N__50503;
    wire N__50502;
    wire N__50501;
    wire N__50500;
    wire N__50499;
    wire N__50498;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50478;
    wire N__50477;
    wire N__50476;
    wire N__50473;
    wire N__50468;
    wire N__50465;
    wire N__50462;
    wire N__50459;
    wire N__50456;
    wire N__50447;
    wire N__50442;
    wire N__50439;
    wire N__50428;
    wire N__50421;
    wire N__50416;
    wire N__50413;
    wire N__50408;
    wire N__50403;
    wire N__50394;
    wire N__50387;
    wire N__50384;
    wire N__50377;
    wire N__50370;
    wire N__50345;
    wire N__50344;
    wire N__50343;
    wire N__50342;
    wire N__50341;
    wire N__50340;
    wire N__50339;
    wire N__50338;
    wire N__50337;
    wire N__50334;
    wire N__50331;
    wire N__50330;
    wire N__50329;
    wire N__50328;
    wire N__50327;
    wire N__50326;
    wire N__50325;
    wire N__50324;
    wire N__50323;
    wire N__50322;
    wire N__50321;
    wire N__50320;
    wire N__50319;
    wire N__50318;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50313;
    wire N__50312;
    wire N__50311;
    wire N__50310;
    wire N__50309;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50297;
    wire N__50294;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50289;
    wire N__50288;
    wire N__50287;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50280;
    wire N__50279;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50275;
    wire N__50274;
    wire N__50273;
    wire N__50272;
    wire N__50271;
    wire N__50270;
    wire N__50269;
    wire N__50268;
    wire N__50267;
    wire N__50266;
    wire N__50265;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50258;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50254;
    wire N__50253;
    wire N__50252;
    wire N__50247;
    wire N__50240;
    wire N__50235;
    wire N__50230;
    wire N__50221;
    wire N__50220;
    wire N__50219;
    wire N__50216;
    wire N__50215;
    wire N__50212;
    wire N__50211;
    wire N__50210;
    wire N__50207;
    wire N__50204;
    wire N__50203;
    wire N__50202;
    wire N__50201;
    wire N__50200;
    wire N__50183;
    wire N__50178;
    wire N__50167;
    wire N__50164;
    wire N__50153;
    wire N__50152;
    wire N__50151;
    wire N__50150;
    wire N__50149;
    wire N__50144;
    wire N__50143;
    wire N__50142;
    wire N__50141;
    wire N__50138;
    wire N__50135;
    wire N__50132;
    wire N__50131;
    wire N__50128;
    wire N__50127;
    wire N__50124;
    wire N__50123;
    wire N__50122;
    wire N__50121;
    wire N__50120;
    wire N__50115;
    wire N__50114;
    wire N__50113;
    wire N__50112;
    wire N__50111;
    wire N__50110;
    wire N__50109;
    wire N__50108;
    wire N__50107;
    wire N__50106;
    wire N__50099;
    wire N__50094;
    wire N__50093;
    wire N__50092;
    wire N__50091;
    wire N__50090;
    wire N__50089;
    wire N__50088;
    wire N__50085;
    wire N__50078;
    wire N__50069;
    wire N__50060;
    wire N__50057;
    wire N__50054;
    wire N__50051;
    wire N__50048;
    wire N__50031;
    wire N__50018;
    wire N__50015;
    wire N__50012;
    wire N__50005;
    wire N__50004;
    wire N__50001;
    wire N__50000;
    wire N__49997;
    wire N__49996;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49980;
    wire N__49977;
    wire N__49972;
    wire N__49967;
    wire N__49966;
    wire N__49965;
    wire N__49962;
    wire N__49957;
    wire N__49952;
    wire N__49943;
    wire N__49940;
    wire N__49939;
    wire N__49938;
    wire N__49935;
    wire N__49932;
    wire N__49929;
    wire N__49924;
    wire N__49921;
    wire N__49914;
    wire N__49911;
    wire N__49902;
    wire N__49899;
    wire N__49898;
    wire N__49897;
    wire N__49896;
    wire N__49895;
    wire N__49894;
    wire N__49893;
    wire N__49892;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49882;
    wire N__49881;
    wire N__49880;
    wire N__49879;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49871;
    wire N__49870;
    wire N__49869;
    wire N__49868;
    wire N__49865;
    wire N__49862;
    wire N__49859;
    wire N__49856;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49836;
    wire N__49831;
    wire N__49820;
    wire N__49819;
    wire N__49806;
    wire N__49795;
    wire N__49792;
    wire N__49779;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49770;
    wire N__49763;
    wire N__49758;
    wire N__49753;
    wire N__49750;
    wire N__49747;
    wire N__49742;
    wire N__49741;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49733;
    wire N__49726;
    wire N__49721;
    wire N__49716;
    wire N__49703;
    wire N__49700;
    wire N__49695;
    wire N__49688;
    wire N__49685;
    wire N__49682;
    wire N__49675;
    wire N__49660;
    wire N__49653;
    wire N__49650;
    wire N__49645;
    wire N__49638;
    wire N__49631;
    wire N__49628;
    wire N__49615;
    wire N__49612;
    wire N__49609;
    wire N__49602;
    wire N__49599;
    wire N__49576;
    wire N__49569;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49547;
    wire N__49546;
    wire N__49545;
    wire N__49544;
    wire N__49543;
    wire N__49542;
    wire N__49541;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49532;
    wire N__49531;
    wire N__49528;
    wire N__49521;
    wire N__49514;
    wire N__49509;
    wire N__49508;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49499;
    wire N__49496;
    wire N__49493;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49481;
    wire N__49480;
    wire N__49479;
    wire N__49474;
    wire N__49473;
    wire N__49472;
    wire N__49471;
    wire N__49470;
    wire N__49469;
    wire N__49464;
    wire N__49453;
    wire N__49450;
    wire N__49447;
    wire N__49446;
    wire N__49445;
    wire N__49442;
    wire N__49439;
    wire N__49438;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49427;
    wire N__49422;
    wire N__49419;
    wire N__49416;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49404;
    wire N__49403;
    wire N__49402;
    wire N__49399;
    wire N__49394;
    wire N__49389;
    wire N__49386;
    wire N__49383;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49360;
    wire N__49357;
    wire N__49348;
    wire N__49343;
    wire N__49338;
    wire N__49335;
    wire N__49328;
    wire N__49321;
    wire N__49298;
    wire N__49295;
    wire N__49292;
    wire N__49289;
    wire N__49286;
    wire N__49285;
    wire N__49282;
    wire N__49281;
    wire N__49278;
    wire N__49273;
    wire N__49268;
    wire N__49267;
    wire N__49266;
    wire N__49265;
    wire N__49264;
    wire N__49263;
    wire N__49262;
    wire N__49257;
    wire N__49256;
    wire N__49253;
    wire N__49244;
    wire N__49243;
    wire N__49242;
    wire N__49241;
    wire N__49240;
    wire N__49239;
    wire N__49238;
    wire N__49237;
    wire N__49234;
    wire N__49233;
    wire N__49232;
    wire N__49231;
    wire N__49228;
    wire N__49227;
    wire N__49226;
    wire N__49225;
    wire N__49222;
    wire N__49221;
    wire N__49220;
    wire N__49217;
    wire N__49214;
    wire N__49213;
    wire N__49212;
    wire N__49209;
    wire N__49206;
    wire N__49205;
    wire N__49204;
    wire N__49203;
    wire N__49202;
    wire N__49201;
    wire N__49200;
    wire N__49199;
    wire N__49198;
    wire N__49197;
    wire N__49196;
    wire N__49195;
    wire N__49194;
    wire N__49193;
    wire N__49192;
    wire N__49191;
    wire N__49190;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49178;
    wire N__49175;
    wire N__49170;
    wire N__49167;
    wire N__49158;
    wire N__49155;
    wire N__49150;
    wire N__49145;
    wire N__49142;
    wire N__49139;
    wire N__49136;
    wire N__49131;
    wire N__49130;
    wire N__49129;
    wire N__49128;
    wire N__49125;
    wire N__49124;
    wire N__49123;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49118;
    wire N__49115;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49108;
    wire N__49107;
    wire N__49102;
    wire N__49095;
    wire N__49090;
    wire N__49079;
    wire N__49078;
    wire N__49077;
    wire N__49074;
    wire N__49071;
    wire N__49066;
    wire N__49061;
    wire N__49056;
    wire N__49049;
    wire N__49046;
    wire N__49043;
    wire N__49040;
    wire N__49037;
    wire N__49030;
    wire N__49029;
    wire N__49024;
    wire N__49021;
    wire N__49020;
    wire N__49013;
    wire N__49012;
    wire N__49011;
    wire N__49008;
    wire N__49007;
    wire N__49004;
    wire N__48993;
    wire N__48988;
    wire N__48979;
    wire N__48978;
    wire N__48977;
    wire N__48972;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48950;
    wire N__48947;
    wire N__48944;
    wire N__48943;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48933;
    wire N__48930;
    wire N__48927;
    wire N__48924;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48905;
    wire N__48900;
    wire N__48889;
    wire N__48884;
    wire N__48879;
    wire N__48868;
    wire N__48845;
    wire N__48842;
    wire N__48841;
    wire N__48840;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48832;
    wire N__48831;
    wire N__48830;
    wire N__48825;
    wire N__48824;
    wire N__48819;
    wire N__48818;
    wire N__48817;
    wire N__48816;
    wire N__48815;
    wire N__48814;
    wire N__48811;
    wire N__48810;
    wire N__48809;
    wire N__48806;
    wire N__48805;
    wire N__48804;
    wire N__48803;
    wire N__48800;
    wire N__48797;
    wire N__48794;
    wire N__48791;
    wire N__48786;
    wire N__48785;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48777;
    wire N__48776;
    wire N__48773;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48763;
    wire N__48758;
    wire N__48757;
    wire N__48756;
    wire N__48755;
    wire N__48752;
    wire N__48749;
    wire N__48746;
    wire N__48741;
    wire N__48736;
    wire N__48735;
    wire N__48734;
    wire N__48733;
    wire N__48728;
    wire N__48723;
    wire N__48718;
    wire N__48715;
    wire N__48712;
    wire N__48707;
    wire N__48704;
    wire N__48701;
    wire N__48698;
    wire N__48693;
    wire N__48686;
    wire N__48681;
    wire N__48680;
    wire N__48679;
    wire N__48678;
    wire N__48671;
    wire N__48668;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48640;
    wire N__48637;
    wire N__48632;
    wire N__48627;
    wire N__48624;
    wire N__48619;
    wire N__48612;
    wire N__48599;
    wire N__48598;
    wire N__48595;
    wire N__48590;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48563;
    wire N__48560;
    wire N__48557;
    wire N__48554;
    wire N__48551;
    wire N__48548;
    wire N__48547;
    wire N__48546;
    wire N__48545;
    wire N__48544;
    wire N__48543;
    wire N__48542;
    wire N__48539;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48533;
    wire N__48530;
    wire N__48529;
    wire N__48528;
    wire N__48527;
    wire N__48526;
    wire N__48525;
    wire N__48524;
    wire N__48523;
    wire N__48522;
    wire N__48521;
    wire N__48520;
    wire N__48519;
    wire N__48518;
    wire N__48517;
    wire N__48510;
    wire N__48507;
    wire N__48506;
    wire N__48505;
    wire N__48504;
    wire N__48503;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48477;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48431;
    wire N__48424;
    wire N__48421;
    wire N__48420;
    wire N__48413;
    wire N__48410;
    wire N__48407;
    wire N__48404;
    wire N__48401;
    wire N__48398;
    wire N__48389;
    wire N__48388;
    wire N__48387;
    wire N__48384;
    wire N__48383;
    wire N__48382;
    wire N__48381;
    wire N__48380;
    wire N__48377;
    wire N__48374;
    wire N__48367;
    wire N__48364;
    wire N__48363;
    wire N__48360;
    wire N__48357;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48335;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48316;
    wire N__48311;
    wire N__48308;
    wire N__48299;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48263;
    wire N__48260;
    wire N__48259;
    wire N__48256;
    wire N__48253;
    wire N__48252;
    wire N__48249;
    wire N__48246;
    wire N__48243;
    wire N__48240;
    wire N__48237;
    wire N__48234;
    wire N__48227;
    wire N__48226;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48212;
    wire N__48209;
    wire N__48206;
    wire N__48203;
    wire N__48202;
    wire N__48201;
    wire N__48198;
    wire N__48195;
    wire N__48192;
    wire N__48189;
    wire N__48186;
    wire N__48179;
    wire N__48176;
    wire N__48173;
    wire N__48172;
    wire N__48169;
    wire N__48166;
    wire N__48163;
    wire N__48158;
    wire N__48155;
    wire N__48152;
    wire N__48149;
    wire N__48146;
    wire N__48143;
    wire N__48140;
    wire N__48139;
    wire N__48136;
    wire N__48133;
    wire N__48130;
    wire N__48127;
    wire N__48122;
    wire N__48119;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48104;
    wire N__48101;
    wire N__48098;
    wire N__48095;
    wire N__48092;
    wire N__48091;
    wire N__48088;
    wire N__48087;
    wire N__48086;
    wire N__48085;
    wire N__48084;
    wire N__48083;
    wire N__48080;
    wire N__48075;
    wire N__48074;
    wire N__48073;
    wire N__48072;
    wire N__48071;
    wire N__48070;
    wire N__48069;
    wire N__48068;
    wire N__48067;
    wire N__48064;
    wire N__48061;
    wire N__48060;
    wire N__48057;
    wire N__48054;
    wire N__48049;
    wire N__48048;
    wire N__48047;
    wire N__48046;
    wire N__48043;
    wire N__48042;
    wire N__48041;
    wire N__48040;
    wire N__48039;
    wire N__48038;
    wire N__48037;
    wire N__48036;
    wire N__48035;
    wire N__48030;
    wire N__48023;
    wire N__48020;
    wire N__48015;
    wire N__48014;
    wire N__48013;
    wire N__48012;
    wire N__48007;
    wire N__48006;
    wire N__48005;
    wire N__48004;
    wire N__48001;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47989;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47983;
    wire N__47980;
    wire N__47977;
    wire N__47974;
    wire N__47971;
    wire N__47966;
    wire N__47963;
    wire N__47958;
    wire N__47955;
    wire N__47948;
    wire N__47945;
    wire N__47944;
    wire N__47941;
    wire N__47938;
    wire N__47935;
    wire N__47930;
    wire N__47929;
    wire N__47928;
    wire N__47925;
    wire N__47924;
    wire N__47923;
    wire N__47922;
    wire N__47921;
    wire N__47920;
    wire N__47919;
    wire N__47918;
    wire N__47917;
    wire N__47916;
    wire N__47915;
    wire N__47914;
    wire N__47913;
    wire N__47912;
    wire N__47911;
    wire N__47910;
    wire N__47909;
    wire N__47902;
    wire N__47895;
    wire N__47888;
    wire N__47877;
    wire N__47866;
    wire N__47865;
    wire N__47864;
    wire N__47861;
    wire N__47860;
    wire N__47859;
    wire N__47856;
    wire N__47855;
    wire N__47854;
    wire N__47853;
    wire N__47852;
    wire N__47849;
    wire N__47844;
    wire N__47841;
    wire N__47838;
    wire N__47835;
    wire N__47828;
    wire N__47825;
    wire N__47824;
    wire N__47823;
    wire N__47822;
    wire N__47817;
    wire N__47816;
    wire N__47815;
    wire N__47812;
    wire N__47811;
    wire N__47810;
    wire N__47807;
    wire N__47806;
    wire N__47805;
    wire N__47804;
    wire N__47803;
    wire N__47802;
    wire N__47801;
    wire N__47800;
    wire N__47799;
    wire N__47798;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47794;
    wire N__47793;
    wire N__47792;
    wire N__47791;
    wire N__47790;
    wire N__47787;
    wire N__47776;
    wire N__47771;
    wire N__47764;
    wire N__47759;
    wire N__47754;
    wire N__47751;
    wire N__47746;
    wire N__47745;
    wire N__47744;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47727;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47711;
    wire N__47708;
    wire N__47703;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47671;
    wire N__47670;
    wire N__47667;
    wire N__47664;
    wire N__47659;
    wire N__47654;
    wire N__47647;
    wire N__47640;
    wire N__47637;
    wire N__47636;
    wire N__47633;
    wire N__47620;
    wire N__47615;
    wire N__47606;
    wire N__47605;
    wire N__47604;
    wire N__47603;
    wire N__47602;
    wire N__47601;
    wire N__47600;
    wire N__47599;
    wire N__47596;
    wire N__47595;
    wire N__47594;
    wire N__47593;
    wire N__47588;
    wire N__47585;
    wire N__47580;
    wire N__47577;
    wire N__47572;
    wire N__47567;
    wire N__47564;
    wire N__47559;
    wire N__47544;
    wire N__47543;
    wire N__47542;
    wire N__47541;
    wire N__47540;
    wire N__47537;
    wire N__47522;
    wire N__47517;
    wire N__47510;
    wire N__47509;
    wire N__47508;
    wire N__47507;
    wire N__47504;
    wire N__47497;
    wire N__47496;
    wire N__47495;
    wire N__47492;
    wire N__47491;
    wire N__47490;
    wire N__47489;
    wire N__47488;
    wire N__47485;
    wire N__47480;
    wire N__47473;
    wire N__47470;
    wire N__47459;
    wire N__47452;
    wire N__47447;
    wire N__47440;
    wire N__47433;
    wire N__47426;
    wire N__47421;
    wire N__47412;
    wire N__47405;
    wire N__47378;
    wire N__47375;
    wire N__47372;
    wire N__47371;
    wire N__47368;
    wire N__47365;
    wire N__47360;
    wire N__47359;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47344;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47336;
    wire N__47335;
    wire N__47330;
    wire N__47327;
    wire N__47326;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47316;
    wire N__47315;
    wire N__47312;
    wire N__47311;
    wire N__47310;
    wire N__47309;
    wire N__47308;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47294;
    wire N__47293;
    wire N__47292;
    wire N__47291;
    wire N__47290;
    wire N__47285;
    wire N__47278;
    wire N__47275;
    wire N__47274;
    wire N__47273;
    wire N__47272;
    wire N__47269;
    wire N__47268;
    wire N__47267;
    wire N__47266;
    wire N__47263;
    wire N__47262;
    wire N__47261;
    wire N__47260;
    wire N__47257;
    wire N__47256;
    wire N__47255;
    wire N__47254;
    wire N__47253;
    wire N__47252;
    wire N__47251;
    wire N__47250;
    wire N__47249;
    wire N__47248;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47244;
    wire N__47243;
    wire N__47240;
    wire N__47239;
    wire N__47238;
    wire N__47237;
    wire N__47236;
    wire N__47233;
    wire N__47232;
    wire N__47231;
    wire N__47230;
    wire N__47227;
    wire N__47224;
    wire N__47217;
    wire N__47214;
    wire N__47209;
    wire N__47206;
    wire N__47199;
    wire N__47196;
    wire N__47191;
    wire N__47188;
    wire N__47185;
    wire N__47184;
    wire N__47183;
    wire N__47182;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47174;
    wire N__47173;
    wire N__47170;
    wire N__47163;
    wire N__47160;
    wire N__47153;
    wire N__47152;
    wire N__47151;
    wire N__47150;
    wire N__47143;
    wire N__47142;
    wire N__47141;
    wire N__47140;
    wire N__47139;
    wire N__47138;
    wire N__47137;
    wire N__47134;
    wire N__47127;
    wire N__47124;
    wire N__47121;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47107;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47095;
    wire N__47094;
    wire N__47089;
    wire N__47088;
    wire N__47087;
    wire N__47086;
    wire N__47085;
    wire N__47084;
    wire N__47081;
    wire N__47078;
    wire N__47077;
    wire N__47072;
    wire N__47065;
    wire N__47060;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47048;
    wire N__47047;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47027;
    wire N__47018;
    wire N__47011;
    wire N__47008;
    wire N__47001;
    wire N__46994;
    wire N__46977;
    wire N__46972;
    wire N__46967;
    wire N__46966;
    wire N__46965;
    wire N__46964;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46952;
    wire N__46947;
    wire N__46946;
    wire N__46943;
    wire N__46938;
    wire N__46935;
    wire N__46932;
    wire N__46931;
    wire N__46924;
    wire N__46917;
    wire N__46912;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46908;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46898;
    wire N__46891;
    wire N__46888;
    wire N__46875;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46835;
    wire N__46834;
    wire N__46833;
    wire N__46830;
    wire N__46827;
    wire N__46820;
    wire N__46819;
    wire N__46818;
    wire N__46817;
    wire N__46814;
    wire N__46811;
    wire N__46806;
    wire N__46799;
    wire N__46796;
    wire N__46787;
    wire N__46772;
    wire N__46765;
    wire N__46758;
    wire N__46751;
    wire N__46748;
    wire N__46743;
    wire N__46718;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46700;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46667;
    wire N__46666;
    wire N__46663;
    wire N__46660;
    wire N__46655;
    wire N__46652;
    wire N__46649;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46639;
    wire N__46638;
    wire N__46635;
    wire N__46630;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46618;
    wire N__46615;
    wire N__46610;
    wire N__46609;
    wire N__46608;
    wire N__46607;
    wire N__46606;
    wire N__46605;
    wire N__46604;
    wire N__46603;
    wire N__46602;
    wire N__46601;
    wire N__46600;
    wire N__46599;
    wire N__46588;
    wire N__46585;
    wire N__46584;
    wire N__46583;
    wire N__46582;
    wire N__46581;
    wire N__46580;
    wire N__46579;
    wire N__46578;
    wire N__46577;
    wire N__46576;
    wire N__46575;
    wire N__46574;
    wire N__46571;
    wire N__46562;
    wire N__46561;
    wire N__46560;
    wire N__46557;
    wire N__46556;
    wire N__46555;
    wire N__46550;
    wire N__46547;
    wire N__46540;
    wire N__46537;
    wire N__46524;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46503;
    wire N__46502;
    wire N__46501;
    wire N__46498;
    wire N__46495;
    wire N__46490;
    wire N__46487;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46471;
    wire N__46470;
    wire N__46469;
    wire N__46466;
    wire N__46465;
    wire N__46464;
    wire N__46463;
    wire N__46462;
    wire N__46457;
    wire N__46450;
    wire N__46447;
    wire N__46442;
    wire N__46437;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46419;
    wire N__46412;
    wire N__46397;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46377;
    wire N__46374;
    wire N__46371;
    wire N__46368;
    wire N__46361;
    wire N__46358;
    wire N__46357;
    wire N__46354;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46338;
    wire N__46331;
    wire N__46328;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46313;
    wire N__46310;
    wire N__46307;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46289;
    wire N__46286;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46272;
    wire N__46269;
    wire N__46266;
    wire N__46263;
    wire N__46256;
    wire N__46253;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46228;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46202;
    wire N__46199;
    wire N__46196;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46181;
    wire N__46178;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46164;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46145;
    wire N__46142;
    wire N__46141;
    wire N__46138;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46126;
    wire N__46121;
    wire N__46120;
    wire N__46119;
    wire N__46118;
    wire N__46117;
    wire N__46116;
    wire N__46115;
    wire N__46112;
    wire N__46109;
    wire N__46108;
    wire N__46097;
    wire N__46090;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46082;
    wire N__46081;
    wire N__46080;
    wire N__46079;
    wire N__46078;
    wire N__46077;
    wire N__46076;
    wire N__46073;
    wire N__46072;
    wire N__46067;
    wire N__46064;
    wire N__46063;
    wire N__46062;
    wire N__46059;
    wire N__46058;
    wire N__46053;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46039;
    wire N__46038;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46028;
    wire N__46025;
    wire N__46022;
    wire N__46019;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46004;
    wire N__46003;
    wire N__46002;
    wire N__46001;
    wire N__45998;
    wire N__45997;
    wire N__45994;
    wire N__45993;
    wire N__45986;
    wire N__45983;
    wire N__45978;
    wire N__45975;
    wire N__45968;
    wire N__45959;
    wire N__45950;
    wire N__45949;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45934;
    wire N__45931;
    wire N__45928;
    wire N__45923;
    wire N__45908;
    wire N__45905;
    wire N__45904;
    wire N__45903;
    wire N__45900;
    wire N__45895;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45881;
    wire N__45878;
    wire N__45877;
    wire N__45874;
    wire N__45871;
    wire N__45868;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45814;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45797;
    wire N__45796;
    wire N__45795;
    wire N__45794;
    wire N__45789;
    wire N__45786;
    wire N__45783;
    wire N__45778;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45754;
    wire N__45751;
    wire N__45746;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45730;
    wire N__45727;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45715;
    wire N__45712;
    wire N__45707;
    wire N__45704;
    wire N__45703;
    wire N__45700;
    wire N__45697;
    wire N__45694;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45676;
    wire N__45673;
    wire N__45670;
    wire N__45667;
    wire N__45662;
    wire N__45661;
    wire N__45660;
    wire N__45659;
    wire N__45658;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45653;
    wire N__45652;
    wire N__45651;
    wire N__45650;
    wire N__45649;
    wire N__45648;
    wire N__45647;
    wire N__45646;
    wire N__45645;
    wire N__45640;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45622;
    wire N__45619;
    wire N__45616;
    wire N__45613;
    wire N__45608;
    wire N__45607;
    wire N__45606;
    wire N__45605;
    wire N__45604;
    wire N__45603;
    wire N__45602;
    wire N__45599;
    wire N__45598;
    wire N__45597;
    wire N__45592;
    wire N__45589;
    wire N__45586;
    wire N__45583;
    wire N__45580;
    wire N__45575;
    wire N__45572;
    wire N__45569;
    wire N__45566;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45546;
    wire N__45545;
    wire N__45544;
    wire N__45543;
    wire N__45542;
    wire N__45541;
    wire N__45540;
    wire N__45539;
    wire N__45538;
    wire N__45537;
    wire N__45536;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45506;
    wire N__45501;
    wire N__45500;
    wire N__45497;
    wire N__45488;
    wire N__45483;
    wire N__45478;
    wire N__45471;
    wire N__45466;
    wire N__45465;
    wire N__45464;
    wire N__45461;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45451;
    wire N__45446;
    wire N__45441;
    wire N__45438;
    wire N__45437;
    wire N__45436;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45416;
    wire N__45415;
    wire N__45414;
    wire N__45413;
    wire N__45412;
    wire N__45411;
    wire N__45410;
    wire N__45409;
    wire N__45406;
    wire N__45405;
    wire N__45402;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45382;
    wire N__45379;
    wire N__45374;
    wire N__45369;
    wire N__45366;
    wire N__45361;
    wire N__45352;
    wire N__45349;
    wire N__45344;
    wire N__45317;
    wire N__45314;
    wire N__45313;
    wire N__45310;
    wire N__45309;
    wire N__45308;
    wire N__45307;
    wire N__45306;
    wire N__45303;
    wire N__45302;
    wire N__45299;
    wire N__45298;
    wire N__45297;
    wire N__45296;
    wire N__45295;
    wire N__45294;
    wire N__45293;
    wire N__45290;
    wire N__45289;
    wire N__45286;
    wire N__45285;
    wire N__45280;
    wire N__45279;
    wire N__45278;
    wire N__45273;
    wire N__45270;
    wire N__45265;
    wire N__45264;
    wire N__45263;
    wire N__45262;
    wire N__45261;
    wire N__45256;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45240;
    wire N__45239;
    wire N__45238;
    wire N__45237;
    wire N__45236;
    wire N__45235;
    wire N__45234;
    wire N__45233;
    wire N__45232;
    wire N__45231;
    wire N__45230;
    wire N__45229;
    wire N__45226;
    wire N__45225;
    wire N__45224;
    wire N__45223;
    wire N__45222;
    wire N__45221;
    wire N__45220;
    wire N__45219;
    wire N__45218;
    wire N__45217;
    wire N__45216;
    wire N__45215;
    wire N__45212;
    wire N__45207;
    wire N__45200;
    wire N__45197;
    wire N__45190;
    wire N__45185;
    wire N__45184;
    wire N__45183;
    wire N__45182;
    wire N__45173;
    wire N__45170;
    wire N__45167;
    wire N__45160;
    wire N__45155;
    wire N__45154;
    wire N__45153;
    wire N__45152;
    wire N__45151;
    wire N__45142;
    wire N__45139;
    wire N__45136;
    wire N__45133;
    wire N__45128;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45109;
    wire N__45106;
    wire N__45105;
    wire N__45096;
    wire N__45091;
    wire N__45084;
    wire N__45079;
    wire N__45076;
    wire N__45071;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45059;
    wire N__45058;
    wire N__45055;
    wire N__45044;
    wire N__45043;
    wire N__45042;
    wire N__45041;
    wire N__45040;
    wire N__45031;
    wire N__45026;
    wire N__45019;
    wire N__45006;
    wire N__45001;
    wire N__44996;
    wire N__44991;
    wire N__44986;
    wire N__44969;
    wire N__44968;
    wire N__44967;
    wire N__44964;
    wire N__44963;
    wire N__44960;
    wire N__44957;
    wire N__44954;
    wire N__44951;
    wire N__44948;
    wire N__44945;
    wire N__44942;
    wire N__44939;
    wire N__44934;
    wire N__44931;
    wire N__44926;
    wire N__44921;
    wire N__44918;
    wire N__44917;
    wire N__44914;
    wire N__44911;
    wire N__44910;
    wire N__44909;
    wire N__44908;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44888;
    wire N__44887;
    wire N__44886;
    wire N__44885;
    wire N__44884;
    wire N__44883;
    wire N__44874;
    wire N__44869;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44839;
    wire N__44834;
    wire N__44831;
    wire N__44828;
    wire N__44825;
    wire N__44822;
    wire N__44813;
    wire N__44808;
    wire N__44807;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44786;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44776;
    wire N__44775;
    wire N__44774;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44732;
    wire N__44727;
    wire N__44722;
    wire N__44717;
    wire N__44716;
    wire N__44713;
    wire N__44712;
    wire N__44711;
    wire N__44708;
    wire N__44705;
    wire N__44702;
    wire N__44699;
    wire N__44698;
    wire N__44695;
    wire N__44690;
    wire N__44687;
    wire N__44684;
    wire N__44681;
    wire N__44678;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44657;
    wire N__44654;
    wire N__44653;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44645;
    wire N__44642;
    wire N__44641;
    wire N__44636;
    wire N__44633;
    wire N__44630;
    wire N__44627;
    wire N__44622;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44603;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44567;
    wire N__44564;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44510;
    wire N__44509;
    wire N__44508;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44494;
    wire N__44491;
    wire N__44486;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44471;
    wire N__44468;
    wire N__44465;
    wire N__44464;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44419;
    wire N__44416;
    wire N__44413;
    wire N__44410;
    wire N__44405;
    wire N__44404;
    wire N__44403;
    wire N__44402;
    wire N__44401;
    wire N__44400;
    wire N__44399;
    wire N__44398;
    wire N__44395;
    wire N__44390;
    wire N__44383;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44369;
    wire N__44368;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44360;
    wire N__44359;
    wire N__44358;
    wire N__44357;
    wire N__44356;
    wire N__44355;
    wire N__44354;
    wire N__44353;
    wire N__44352;
    wire N__44351;
    wire N__44348;
    wire N__44345;
    wire N__44340;
    wire N__44337;
    wire N__44332;
    wire N__44331;
    wire N__44326;
    wire N__44321;
    wire N__44314;
    wire N__44311;
    wire N__44308;
    wire N__44303;
    wire N__44302;
    wire N__44299;
    wire N__44294;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44255;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44225;
    wire N__44214;
    wire N__44207;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44180;
    wire N__44179;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44171;
    wire N__44168;
    wire N__44163;
    wire N__44160;
    wire N__44159;
    wire N__44158;
    wire N__44157;
    wire N__44156;
    wire N__44155;
    wire N__44152;
    wire N__44151;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44119;
    wire N__44116;
    wire N__44113;
    wire N__44108;
    wire N__44105;
    wire N__44100;
    wire N__44099;
    wire N__44098;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44081;
    wire N__44078;
    wire N__44075;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44056;
    wire N__44053;
    wire N__44042;
    wire N__44041;
    wire N__44040;
    wire N__44039;
    wire N__44036;
    wire N__44035;
    wire N__44034;
    wire N__44033;
    wire N__44032;
    wire N__44029;
    wire N__44024;
    wire N__44021;
    wire N__44012;
    wire N__44003;
    wire N__44002;
    wire N__44001;
    wire N__43998;
    wire N__43997;
    wire N__43996;
    wire N__43995;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43981;
    wire N__43974;
    wire N__43967;
    wire N__43966;
    wire N__43963;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43937;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43909;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43892;
    wire N__43891;
    wire N__43890;
    wire N__43887;
    wire N__43880;
    wire N__43877;
    wire N__43874;
    wire N__43873;
    wire N__43870;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43858;
    wire N__43853;
    wire N__43850;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43827;
    wire N__43822;
    wire N__43819;
    wire N__43814;
    wire N__43811;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43778;
    wire N__43775;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43753;
    wire N__43748;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43738;
    wire N__43735;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43723;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43709;
    wire N__43708;
    wire N__43707;
    wire N__43704;
    wire N__43699;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43681;
    wire N__43678;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43668;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43636;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43621;
    wire N__43616;
    wire N__43615;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43596;
    wire N__43593;
    wire N__43590;
    wire N__43585;
    wire N__43580;
    wire N__43577;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43562;
    wire N__43561;
    wire N__43560;
    wire N__43559;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43534;
    wire N__43533;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43502;
    wire N__43493;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43451;
    wire N__43450;
    wire N__43449;
    wire N__43448;
    wire N__43447;
    wire N__43446;
    wire N__43445;
    wire N__43442;
    wire N__43441;
    wire N__43440;
    wire N__43439;
    wire N__43438;
    wire N__43437;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43421;
    wire N__43418;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43406;
    wire N__43403;
    wire N__43402;
    wire N__43399;
    wire N__43398;
    wire N__43395;
    wire N__43394;
    wire N__43393;
    wire N__43392;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43380;
    wire N__43379;
    wire N__43376;
    wire N__43371;
    wire N__43362;
    wire N__43359;
    wire N__43350;
    wire N__43343;
    wire N__43340;
    wire N__43333;
    wire N__43330;
    wire N__43323;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43311;
    wire N__43304;
    wire N__43301;
    wire N__43300;
    wire N__43299;
    wire N__43298;
    wire N__43297;
    wire N__43290;
    wire N__43289;
    wire N__43288;
    wire N__43287;
    wire N__43282;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43268;
    wire N__43267;
    wire N__43266;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43256;
    wire N__43255;
    wire N__43248;
    wire N__43239;
    wire N__43238;
    wire N__43235;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43221;
    wire N__43218;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43198;
    wire N__43197;
    wire N__43194;
    wire N__43189;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43174;
    wire N__43171;
    wire N__43166;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43138;
    wire N__43135;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43127;
    wire N__43126;
    wire N__43123;
    wire N__43122;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43110;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43066;
    wire N__43063;
    wire N__43058;
    wire N__43051;
    wire N__43048;
    wire N__43045;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43017;
    wire N__43012;
    wire N__43009;
    wire N__43006;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42935;
    wire N__42932;
    wire N__42931;
    wire N__42928;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42916;
    wire N__42913;
    wire N__42908;
    wire N__42905;
    wire N__42904;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42890;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42862;
    wire N__42857;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42839;
    wire N__42838;
    wire N__42833;
    wire N__42830;
    wire N__42825;
    wire N__42820;
    wire N__42815;
    wire N__42812;
    wire N__42811;
    wire N__42808;
    wire N__42805;
    wire N__42800;
    wire N__42799;
    wire N__42798;
    wire N__42797;
    wire N__42796;
    wire N__42795;
    wire N__42788;
    wire N__42785;
    wire N__42780;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42748;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42731;
    wire N__42728;
    wire N__42727;
    wire N__42726;
    wire N__42723;
    wire N__42718;
    wire N__42713;
    wire N__42710;
    wire N__42707;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42653;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42632;
    wire N__42629;
    wire N__42626;
    wire N__42623;
    wire N__42620;
    wire N__42617;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42602;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42581;
    wire N__42580;
    wire N__42577;
    wire N__42574;
    wire N__42571;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42557;
    wire N__42554;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42539;
    wire N__42536;
    wire N__42533;
    wire N__42530;
    wire N__42527;
    wire N__42524;
    wire N__42523;
    wire N__42520;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42490;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42466;
    wire N__42465;
    wire N__42464;
    wire N__42463;
    wire N__42462;
    wire N__42461;
    wire N__42460;
    wire N__42459;
    wire N__42456;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42448;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42440;
    wire N__42439;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42424;
    wire N__42421;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42404;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42385;
    wire N__42382;
    wire N__42381;
    wire N__42376;
    wire N__42375;
    wire N__42372;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42353;
    wire N__42350;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42314;
    wire N__42307;
    wire N__42302;
    wire N__42299;
    wire N__42294;
    wire N__42285;
    wire N__42280;
    wire N__42277;
    wire N__42272;
    wire N__42269;
    wire N__42260;
    wire N__42257;
    wire N__42254;
    wire N__42253;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42236;
    wire N__42233;
    wire N__42232;
    wire N__42229;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42191;
    wire N__42188;
    wire N__42187;
    wire N__42184;
    wire N__42181;
    wire N__42178;
    wire N__42177;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42161;
    wire N__42160;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42150;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42124;
    wire N__42121;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42095;
    wire N__42092;
    wire N__42089;
    wire N__42088;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42073;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42059;
    wire N__42056;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42044;
    wire N__42041;
    wire N__42038;
    wire N__42035;
    wire N__42032;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42017;
    wire N__42016;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41969;
    wire N__41966;
    wire N__41963;
    wire N__41960;
    wire N__41957;
    wire N__41956;
    wire N__41953;
    wire N__41950;
    wire N__41949;
    wire N__41944;
    wire N__41941;
    wire N__41936;
    wire N__41935;
    wire N__41932;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41914;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41897;
    wire N__41896;
    wire N__41895;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41869;
    wire N__41864;
    wire N__41863;
    wire N__41860;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41846;
    wire N__41843;
    wire N__41838;
    wire N__41835;
    wire N__41828;
    wire N__41827;
    wire N__41826;
    wire N__41825;
    wire N__41824;
    wire N__41823;
    wire N__41822;
    wire N__41821;
    wire N__41820;
    wire N__41819;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41807;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41791;
    wire N__41790;
    wire N__41789;
    wire N__41786;
    wire N__41785;
    wire N__41782;
    wire N__41779;
    wire N__41776;
    wire N__41773;
    wire N__41766;
    wire N__41761;
    wire N__41758;
    wire N__41757;
    wire N__41756;
    wire N__41753;
    wire N__41746;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41719;
    wire N__41708;
    wire N__41705;
    wire N__41704;
    wire N__41701;
    wire N__41698;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41675;
    wire N__41674;
    wire N__41671;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41657;
    wire N__41656;
    wire N__41653;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41578;
    wire N__41575;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41558;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41550;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41528;
    wire N__41527;
    wire N__41526;
    wire N__41525;
    wire N__41524;
    wire N__41521;
    wire N__41520;
    wire N__41519;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41511;
    wire N__41510;
    wire N__41507;
    wire N__41506;
    wire N__41505;
    wire N__41502;
    wire N__41499;
    wire N__41498;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41429;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41404;
    wire N__41399;
    wire N__41396;
    wire N__41391;
    wire N__41388;
    wire N__41381;
    wire N__41380;
    wire N__41379;
    wire N__41378;
    wire N__41375;
    wire N__41374;
    wire N__41373;
    wire N__41370;
    wire N__41369;
    wire N__41368;
    wire N__41365;
    wire N__41362;
    wire N__41361;
    wire N__41360;
    wire N__41357;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41315;
    wire N__41314;
    wire N__41313;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41301;
    wire N__41288;
    wire N__41285;
    wire N__41280;
    wire N__41277;
    wire N__41272;
    wire N__41269;
    wire N__41258;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41227;
    wire N__41222;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41211;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41201;
    wire N__41200;
    wire N__41197;
    wire N__41190;
    wire N__41187;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41170;
    wire N__41169;
    wire N__41168;
    wire N__41167;
    wire N__41166;
    wire N__41161;
    wire N__41158;
    wire N__41155;
    wire N__41152;
    wire N__41151;
    wire N__41148;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41105;
    wire N__41102;
    wire N__41101;
    wire N__41098;
    wire N__41097;
    wire N__41096;
    wire N__41093;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41063;
    wire N__41060;
    wire N__41055;
    wire N__41052;
    wire N__41045;
    wire N__41044;
    wire N__41041;
    wire N__41040;
    wire N__41039;
    wire N__41038;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41021;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41003;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40990;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40969;
    wire N__40966;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40951;
    wire N__40946;
    wire N__40945;
    wire N__40944;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40930;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40907;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40889;
    wire N__40886;
    wire N__40885;
    wire N__40884;
    wire N__40881;
    wire N__40880;
    wire N__40879;
    wire N__40876;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40864;
    wire N__40863;
    wire N__40862;
    wire N__40861;
    wire N__40860;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40830;
    wire N__40827;
    wire N__40822;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40784;
    wire N__40783;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40759;
    wire N__40754;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40739;
    wire N__40736;
    wire N__40733;
    wire N__40732;
    wire N__40731;
    wire N__40730;
    wire N__40727;
    wire N__40724;
    wire N__40723;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40715;
    wire N__40710;
    wire N__40707;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40693;
    wire N__40692;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40657;
    wire N__40652;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40632;
    wire N__40629;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40595;
    wire N__40592;
    wire N__40589;
    wire N__40586;
    wire N__40583;
    wire N__40580;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40565;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40550;
    wire N__40547;
    wire N__40546;
    wire N__40545;
    wire N__40544;
    wire N__40543;
    wire N__40540;
    wire N__40535;
    wire N__40534;
    wire N__40533;
    wire N__40532;
    wire N__40529;
    wire N__40528;
    wire N__40525;
    wire N__40520;
    wire N__40517;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40505;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40477;
    wire N__40472;
    wire N__40471;
    wire N__40470;
    wire N__40465;
    wire N__40464;
    wire N__40463;
    wire N__40462;
    wire N__40461;
    wire N__40460;
    wire N__40459;
    wire N__40458;
    wire N__40457;
    wire N__40456;
    wire N__40455;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40438;
    wire N__40435;
    wire N__40434;
    wire N__40433;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40408;
    wire N__40405;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40368;
    wire N__40365;
    wire N__40358;
    wire N__40349;
    wire N__40346;
    wire N__40345;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40325;
    wire N__40324;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40314;
    wire N__40309;
    wire N__40304;
    wire N__40303;
    wire N__40302;
    wire N__40299;
    wire N__40294;
    wire N__40289;
    wire N__40288;
    wire N__40285;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40268;
    wire N__40267;
    wire N__40266;
    wire N__40263;
    wire N__40258;
    wire N__40253;
    wire N__40252;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40241;
    wire N__40240;
    wire N__40239;
    wire N__40238;
    wire N__40237;
    wire N__40234;
    wire N__40229;
    wire N__40226;
    wire N__40225;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40213;
    wire N__40212;
    wire N__40211;
    wire N__40210;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40196;
    wire N__40195;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40165;
    wire N__40164;
    wire N__40161;
    wire N__40156;
    wire N__40151;
    wire N__40148;
    wire N__40143;
    wire N__40140;
    wire N__40135;
    wire N__40124;
    wire N__40123;
    wire N__40122;
    wire N__40121;
    wire N__40120;
    wire N__40119;
    wire N__40118;
    wire N__40117;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40082;
    wire N__40077;
    wire N__40076;
    wire N__40075;
    wire N__40068;
    wire N__40065;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40040;
    wire N__40037;
    wire N__40036;
    wire N__40033;
    wire N__40028;
    wire N__40025;
    wire N__40022;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40010;
    wire N__40007;
    wire N__39998;
    wire N__39997;
    wire N__39996;
    wire N__39995;
    wire N__39992;
    wire N__39989;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39970;
    wire N__39965;
    wire N__39960;
    wire N__39957;
    wire N__39952;
    wire N__39947;
    wire N__39944;
    wire N__39941;
    wire N__39940;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39932;
    wire N__39929;
    wire N__39928;
    wire N__39923;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39915;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39905;
    wire N__39904;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39887;
    wire N__39882;
    wire N__39879;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39863;
    wire N__39860;
    wire N__39859;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39841;
    wire N__39838;
    wire N__39833;
    wire N__39832;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39812;
    wire N__39809;
    wire N__39808;
    wire N__39805;
    wire N__39804;
    wire N__39803;
    wire N__39802;
    wire N__39799;
    wire N__39798;
    wire N__39797;
    wire N__39796;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39766;
    wire N__39765;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39746;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39731;
    wire N__39728;
    wire N__39723;
    wire N__39720;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39700;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39688;
    wire N__39685;
    wire N__39682;
    wire N__39677;
    wire N__39674;
    wire N__39665;
    wire N__39664;
    wire N__39663;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39655;
    wire N__39654;
    wire N__39651;
    wire N__39650;
    wire N__39647;
    wire N__39644;
    wire N__39641;
    wire N__39640;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39622;
    wire N__39619;
    wire N__39614;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39581;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39570;
    wire N__39569;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39557;
    wire N__39556;
    wire N__39553;
    wire N__39552;
    wire N__39549;
    wire N__39544;
    wire N__39543;
    wire N__39542;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39476;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39397;
    wire N__39396;
    wire N__39395;
    wire N__39394;
    wire N__39391;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39361;
    wire N__39360;
    wire N__39355;
    wire N__39350;
    wire N__39347;
    wire N__39342;
    wire N__39339;
    wire N__39338;
    wire N__39335;
    wire N__39334;
    wire N__39333;
    wire N__39328;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39256;
    wire N__39255;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39239;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39227;
    wire N__39224;
    wire N__39215;
    wire N__39214;
    wire N__39213;
    wire N__39210;
    wire N__39209;
    wire N__39206;
    wire N__39205;
    wire N__39202;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39188;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39180;
    wire N__39179;
    wire N__39178;
    wire N__39177;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39142;
    wire N__39135;
    wire N__39132;
    wire N__39119;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39092;
    wire N__39083;
    wire N__39082;
    wire N__39077;
    wire N__39074;
    wire N__39073;
    wire N__39068;
    wire N__39065;
    wire N__39062;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39044;
    wire N__39041;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38996;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38977;
    wire N__38976;
    wire N__38973;
    wire N__38972;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38939;
    wire N__38936;
    wire N__38927;
    wire N__38926;
    wire N__38925;
    wire N__38924;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38904;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38854;
    wire N__38849;
    wire N__38848;
    wire N__38847;
    wire N__38846;
    wire N__38845;
    wire N__38844;
    wire N__38843;
    wire N__38842;
    wire N__38841;
    wire N__38840;
    wire N__38839;
    wire N__38838;
    wire N__38837;
    wire N__38836;
    wire N__38835;
    wire N__38834;
    wire N__38833;
    wire N__38832;
    wire N__38831;
    wire N__38830;
    wire N__38829;
    wire N__38828;
    wire N__38827;
    wire N__38826;
    wire N__38825;
    wire N__38824;
    wire N__38823;
    wire N__38822;
    wire N__38821;
    wire N__38816;
    wire N__38811;
    wire N__38810;
    wire N__38809;
    wire N__38802;
    wire N__38795;
    wire N__38790;
    wire N__38789;
    wire N__38788;
    wire N__38787;
    wire N__38786;
    wire N__38785;
    wire N__38784;
    wire N__38783;
    wire N__38782;
    wire N__38781;
    wire N__38780;
    wire N__38779;
    wire N__38776;
    wire N__38767;
    wire N__38766;
    wire N__38765;
    wire N__38764;
    wire N__38763;
    wire N__38760;
    wire N__38753;
    wire N__38746;
    wire N__38735;
    wire N__38730;
    wire N__38725;
    wire N__38718;
    wire N__38711;
    wire N__38704;
    wire N__38699;
    wire N__38694;
    wire N__38693;
    wire N__38690;
    wire N__38689;
    wire N__38686;
    wire N__38683;
    wire N__38680;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38655;
    wire N__38646;
    wire N__38643;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38631;
    wire N__38630;
    wire N__38619;
    wire N__38614;
    wire N__38609;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38564;
    wire N__38561;
    wire N__38560;
    wire N__38559;
    wire N__38558;
    wire N__38555;
    wire N__38552;
    wire N__38549;
    wire N__38548;
    wire N__38545;
    wire N__38538;
    wire N__38535;
    wire N__38534;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38511;
    wire N__38508;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38485;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38420;
    wire N__38419;
    wire N__38418;
    wire N__38417;
    wire N__38416;
    wire N__38415;
    wire N__38414;
    wire N__38413;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38391;
    wire N__38384;
    wire N__38381;
    wire N__38378;
    wire N__38377;
    wire N__38376;
    wire N__38375;
    wire N__38374;
    wire N__38373;
    wire N__38372;
    wire N__38371;
    wire N__38368;
    wire N__38353;
    wire N__38348;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38333;
    wire N__38332;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38284;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38269;
    wire N__38266;
    wire N__38261;
    wire N__38258;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38243;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38228;
    wire N__38227;
    wire N__38224;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38193;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38174;
    wire N__38171;
    wire N__38170;
    wire N__38167;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38150;
    wire N__38147;
    wire N__38146;
    wire N__38145;
    wire N__38142;
    wire N__38137;
    wire N__38132;
    wire N__38131;
    wire N__38128;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38108;
    wire N__38103;
    wire N__38098;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38090;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38074;
    wire N__38071;
    wire N__38064;
    wire N__38061;
    wire N__38048;
    wire N__38047;
    wire N__38044;
    wire N__38043;
    wire N__38042;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38016;
    wire N__38011;
    wire N__38006;
    wire N__38005;
    wire N__38002;
    wire N__37999;
    wire N__37996;
    wire N__37995;
    wire N__37994;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37949;
    wire N__37946;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37921;
    wire N__37918;
    wire N__37917;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37882;
    wire N__37879;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37871;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37829;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37811;
    wire N__37810;
    wire N__37807;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37778;
    wire N__37775;
    wire N__37772;
    wire N__37771;
    wire N__37768;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37758;
    wire N__37755;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37741;
    wire N__37740;
    wire N__37737;
    wire N__37732;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37693;
    wire N__37688;
    wire N__37687;
    wire N__37684;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37649;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37634;
    wire N__37631;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37615;
    wire N__37610;
    wire N__37607;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37586;
    wire N__37583;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37520;
    wire N__37517;
    wire N__37516;
    wire N__37513;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37496;
    wire N__37493;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37462;
    wire N__37461;
    wire N__37458;
    wire N__37453;
    wire N__37450;
    wire N__37445;
    wire N__37442;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37432;
    wire N__37427;
    wire N__37424;
    wire N__37423;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37408;
    wire N__37403;
    wire N__37400;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37387;
    wire N__37384;
    wire N__37381;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37349;
    wire N__37346;
    wire N__37345;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37318;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37285;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37273;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37241;
    wire N__37238;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37193;
    wire N__37190;
    wire N__37189;
    wire N__37186;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37172;
    wire N__37169;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36994;
    wire N__36991;
    wire N__36990;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36973;
    wire N__36972;
    wire N__36969;
    wire N__36968;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36920;
    wire N__36915;
    wire N__36908;
    wire N__36903;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36852;
    wire N__36845;
    wire N__36844;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36793;
    wire N__36790;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36763;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36748;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36715;
    wire N__36714;
    wire N__36713;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36662;
    wire N__36653;
    wire N__36650;
    wire N__36649;
    wire N__36648;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36595;
    wire N__36590;
    wire N__36587;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36505;
    wire N__36502;
    wire N__36499;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36485;
    wire N__36484;
    wire N__36479;
    wire N__36476;
    wire N__36475;
    wire N__36474;
    wire N__36471;
    wire N__36470;
    wire N__36467;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36457;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36438;
    wire N__36435;
    wire N__36434;
    wire N__36433;
    wire N__36430;
    wire N__36429;
    wire N__36428;
    wire N__36425;
    wire N__36416;
    wire N__36411;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36393;
    wire N__36390;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36358;
    wire N__36357;
    wire N__36352;
    wire N__36349;
    wire N__36344;
    wire N__36343;
    wire N__36342;
    wire N__36341;
    wire N__36334;
    wire N__36331;
    wire N__36326;
    wire N__36323;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36310;
    wire N__36307;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35873;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35787;
    wire N__35784;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35765;
    wire N__35764;
    wire N__35763;
    wire N__35760;
    wire N__35759;
    wire N__35756;
    wire N__35755;
    wire N__35754;
    wire N__35753;
    wire N__35752;
    wire N__35749;
    wire N__35748;
    wire N__35747;
    wire N__35746;
    wire N__35743;
    wire N__35742;
    wire N__35741;
    wire N__35738;
    wire N__35737;
    wire N__35736;
    wire N__35735;
    wire N__35734;
    wire N__35733;
    wire N__35732;
    wire N__35731;
    wire N__35730;
    wire N__35729;
    wire N__35728;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35688;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35670;
    wire N__35669;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35636;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35617;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35609;
    wire N__35608;
    wire N__35605;
    wire N__35600;
    wire N__35599;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35572;
    wire N__35569;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35517;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35193;
    wire N__35190;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35135;
    wire N__35132;
    wire N__35129;
    wire N__35126;
    wire N__35123;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34945;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34921;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34900;
    wire N__34897;
    wire N__34892;
    wire N__34889;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34859;
    wire N__34856;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34823;
    wire N__34820;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34790;
    wire N__34787;
    wire N__34786;
    wire N__34783;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34768;
    wire N__34763;
    wire N__34760;
    wire N__34759;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34661;
    wire N__34658;
    wire N__34657;
    wire N__34654;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34592;
    wire N__34591;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34560;
    wire N__34551;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34523;
    wire N__34520;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34503;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34480;
    wire N__34475;
    wire N__34474;
    wire N__34471;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34445;
    wire N__34442;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34427;
    wire N__34424;
    wire N__34423;
    wire N__34420;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34409;
    wire N__34408;
    wire N__34407;
    wire N__34400;
    wire N__34397;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34385;
    wire N__34382;
    wire N__34377;
    wire N__34374;
    wire N__34373;
    wire N__34370;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34352;
    wire N__34349;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34327;
    wire N__34322;
    wire N__34319;
    wire N__34318;
    wire N__34315;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34285;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34234;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34214;
    wire N__34211;
    wire N__34210;
    wire N__34207;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34190;
    wire N__34187;
    wire N__34186;
    wire N__34181;
    wire N__34178;
    wire N__34177;
    wire N__34176;
    wire N__34173;
    wire N__34168;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34142;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34134;
    wire N__34133;
    wire N__34130;
    wire N__34125;
    wire N__34124;
    wire N__34121;
    wire N__34120;
    wire N__34119;
    wire N__34118;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34102;
    wire N__34099;
    wire N__34094;
    wire N__34089;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34060;
    wire N__34059;
    wire N__34056;
    wire N__34051;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34030;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34015;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33970;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33962;
    wire N__33961;
    wire N__33958;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33907;
    wire N__33904;
    wire N__33903;
    wire N__33900;
    wire N__33897;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33882;
    wire N__33875;
    wire N__33872;
    wire N__33871;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33856;
    wire N__33851;
    wire N__33850;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33793;
    wire N__33790;
    wire N__33789;
    wire N__33786;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33775;
    wire N__33772;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33752;
    wire N__33749;
    wire N__33744;
    wire N__33741;
    wire N__33736;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33704;
    wire N__33701;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33669;
    wire N__33666;
    wire N__33661;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33649;
    wire N__33646;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33628;
    wire N__33627;
    wire N__33626;
    wire N__33625;
    wire N__33622;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33603;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33559;
    wire N__33556;
    wire N__33555;
    wire N__33552;
    wire N__33551;
    wire N__33548;
    wire N__33541;
    wire N__33536;
    wire N__33535;
    wire N__33534;
    wire N__33533;
    wire N__33532;
    wire N__33531;
    wire N__33526;
    wire N__33525;
    wire N__33524;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33520;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33502;
    wire N__33495;
    wire N__33492;
    wire N__33491;
    wire N__33490;
    wire N__33489;
    wire N__33488;
    wire N__33487;
    wire N__33486;
    wire N__33485;
    wire N__33484;
    wire N__33483;
    wire N__33480;
    wire N__33471;
    wire N__33468;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33449;
    wire N__33448;
    wire N__33441;
    wire N__33436;
    wire N__33431;
    wire N__33424;
    wire N__33419;
    wire N__33416;
    wire N__33415;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33389;
    wire N__33374;
    wire N__33373;
    wire N__33372;
    wire N__33371;
    wire N__33368;
    wire N__33363;
    wire N__33358;
    wire N__33353;
    wire N__33352;
    wire N__33351;
    wire N__33350;
    wire N__33349;
    wire N__33348;
    wire N__33347;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33332;
    wire N__33331;
    wire N__33330;
    wire N__33329;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33317;
    wire N__33312;
    wire N__33307;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33272;
    wire N__33269;
    wire N__33262;
    wire N__33255;
    wire N__33252;
    wire N__33251;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33239;
    wire N__33234;
    wire N__33229;
    wire N__33226;
    wire N__33215;
    wire N__33212;
    wire N__33211;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33207;
    wire N__33206;
    wire N__33205;
    wire N__33202;
    wire N__33195;
    wire N__33188;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33180;
    wire N__33179;
    wire N__33178;
    wire N__33177;
    wire N__33176;
    wire N__33175;
    wire N__33174;
    wire N__33173;
    wire N__33172;
    wire N__33171;
    wire N__33170;
    wire N__33169;
    wire N__33168;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33146;
    wire N__33141;
    wire N__33138;
    wire N__33133;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33121;
    wire N__33118;
    wire N__33117;
    wire N__33116;
    wire N__33113;
    wire N__33112;
    wire N__33111;
    wire N__33110;
    wire N__33107;
    wire N__33106;
    wire N__33105;
    wire N__33104;
    wire N__33103;
    wire N__33102;
    wire N__33101;
    wire N__33100;
    wire N__33099;
    wire N__33098;
    wire N__33097;
    wire N__33096;
    wire N__33091;
    wire N__33086;
    wire N__33085;
    wire N__33080;
    wire N__33077;
    wire N__33070;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33052;
    wire N__33041;
    wire N__33038;
    wire N__33031;
    wire N__33028;
    wire N__33021;
    wire N__33020;
    wire N__33015;
    wire N__33012;
    wire N__33007;
    wire N__33002;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32964;
    wire N__32959;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32938;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32926;
    wire N__32925;
    wire N__32924;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32916;
    wire N__32913;
    wire N__32912;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32900;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32889;
    wire N__32882;
    wire N__32879;
    wire N__32878;
    wire N__32877;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32858;
    wire N__32853;
    wire N__32840;
    wire N__32837;
    wire N__32836;
    wire N__32835;
    wire N__32834;
    wire N__32833;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32815;
    wire N__32814;
    wire N__32813;
    wire N__32812;
    wire N__32811;
    wire N__32810;
    wire N__32809;
    wire N__32808;
    wire N__32803;
    wire N__32798;
    wire N__32795;
    wire N__32790;
    wire N__32785;
    wire N__32782;
    wire N__32771;
    wire N__32768;
    wire N__32767;
    wire N__32764;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32737;
    wire N__32736;
    wire N__32735;
    wire N__32730;
    wire N__32729;
    wire N__32728;
    wire N__32725;
    wire N__32722;
    wire N__32715;
    wire N__32712;
    wire N__32707;
    wire N__32704;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32688;
    wire N__32685;
    wire N__32682;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32662;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32652;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32623;
    wire N__32620;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32590;
    wire N__32587;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32559;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32543;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32501;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32489;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32440;
    wire N__32437;
    wire N__32434;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32383;
    wire N__32378;
    wire N__32375;
    wire N__32372;
    wire N__32371;
    wire N__32368;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32333;
    wire N__32324;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32291;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32276;
    wire N__32273;
    wire N__32272;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32216;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32166;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32140;
    wire N__32137;
    wire N__32134;
    wire N__32131;
    wire N__32126;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32108;
    wire N__32105;
    wire N__32104;
    wire N__32101;
    wire N__32098;
    wire N__32095;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32081;
    wire N__32078;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32056;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32039;
    wire N__32038;
    wire N__32035;
    wire N__32032;
    wire N__32031;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32009;
    wire N__32006;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31991;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31972;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31946;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31912;
    wire N__31911;
    wire N__31908;
    wire N__31903;
    wire N__31900;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31885;
    wire N__31884;
    wire N__31881;
    wire N__31876;
    wire N__31871;
    wire N__31870;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31849;
    wire N__31848;
    wire N__31847;
    wire N__31846;
    wire N__31843;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31824;
    wire N__31819;
    wire N__31816;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31784;
    wire N__31783;
    wire N__31782;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31745;
    wire N__31742;
    wire N__31739;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31729;
    wire N__31728;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31705;
    wire N__31704;
    wire N__31703;
    wire N__31702;
    wire N__31701;
    wire N__31700;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31674;
    wire N__31673;
    wire N__31670;
    wire N__31663;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31641;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31598;
    wire N__31597;
    wire N__31594;
    wire N__31589;
    wire N__31584;
    wire N__31577;
    wire N__31576;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31553;
    wire N__31550;
    wire N__31549;
    wire N__31546;
    wire N__31543;
    wire N__31540;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31498;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31457;
    wire N__31456;
    wire N__31453;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31423;
    wire N__31422;
    wire N__31419;
    wire N__31414;
    wire N__31409;
    wire N__31408;
    wire N__31407;
    wire N__31404;
    wire N__31399;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31336;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31210;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31193;
    wire N__31190;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31144;
    wire N__31143;
    wire N__31142;
    wire N__31139;
    wire N__31132;
    wire N__31129;
    wire N__31124;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31112;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31075;
    wire N__31074;
    wire N__31073;
    wire N__31070;
    wire N__31065;
    wire N__31062;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__31000;
    wire N__30997;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30979;
    wire N__30976;
    wire N__30971;
    wire N__30968;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30887;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30845;
    wire N__30844;
    wire N__30843;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30835;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30800;
    wire N__30795;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30751;
    wire N__30748;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30707;
    wire N__30704;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30656;
    wire N__30655;
    wire N__30654;
    wire N__30649;
    wire N__30648;
    wire N__30647;
    wire N__30642;
    wire N__30637;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30622;
    wire N__30619;
    wire N__30618;
    wire N__30615;
    wire N__30610;
    wire N__30605;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30578;
    wire N__30577;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30542;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30497;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30385;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30259;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30249;
    wire N__30244;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30232;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30215;
    wire N__30214;
    wire N__30213;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30186;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30151;
    wire N__30148;
    wire N__30143;
    wire N__30140;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30125;
    wire N__30122;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30107;
    wire N__30106;
    wire N__30105;
    wire N__30102;
    wire N__30097;
    wire N__30094;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30062;
    wire N__30059;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30032;
    wire N__30029;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30004;
    wire N__30003;
    wire N__30000;
    wire N__29995;
    wire N__29992;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29977;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29960;
    wire N__29959;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29947;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29932;
    wire N__29927;
    wire N__29926;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29904;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29888;
    wire N__29887;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29759;
    wire N__29756;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29741;
    wire N__29738;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29710;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29692;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29585;
    wire N__29582;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29546;
    wire N__29545;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29512;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29489;
    wire N__29488;
    wire N__29485;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29428;
    wire N__29425;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29228;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29061;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29029;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28949;
    wire N__28946;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28897;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28849;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28838;
    wire N__28837;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28823;
    wire N__28822;
    wire N__28821;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28807;
    wire N__28806;
    wire N__28803;
    wire N__28802;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28782;
    wire N__28775;
    wire N__28774;
    wire N__28773;
    wire N__28772;
    wire N__28771;
    wire N__28770;
    wire N__28769;
    wire N__28768;
    wire N__28767;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28752;
    wire N__28751;
    wire N__28744;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28699;
    wire N__28696;
    wire N__28691;
    wire N__28686;
    wire N__28679;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28615;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28558;
    wire N__28555;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28501;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28489;
    wire N__28484;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28364;
    wire N__28363;
    wire N__28360;
    wire N__28359;
    wire N__28358;
    wire N__28355;
    wire N__28354;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28346;
    wire N__28345;
    wire N__28344;
    wire N__28341;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28326;
    wire N__28323;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28305;
    wire N__28302;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28273;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28226;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28066;
    wire N__28065;
    wire N__28062;
    wire N__28057;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27955;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27939;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27866;
    wire N__27863;
    wire N__27862;
    wire N__27861;
    wire N__27860;
    wire N__27857;
    wire N__27856;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27842;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27688;
    wire N__27687;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27658;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27575;
    wire N__27572;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27527;
    wire N__27526;
    wire N__27525;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27517;
    wire N__27516;
    wire N__27515;
    wire N__27514;
    wire N__27513;
    wire N__27512;
    wire N__27511;
    wire N__27506;
    wire N__27503;
    wire N__27490;
    wire N__27489;
    wire N__27486;
    wire N__27485;
    wire N__27484;
    wire N__27483;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27472;
    wire N__27471;
    wire N__27470;
    wire N__27469;
    wire N__27468;
    wire N__27467;
    wire N__27466;
    wire N__27465;
    wire N__27464;
    wire N__27461;
    wire N__27460;
    wire N__27459;
    wire N__27454;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27450;
    wire N__27449;
    wire N__27448;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27429;
    wire N__27416;
    wire N__27415;
    wire N__27412;
    wire N__27411;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27403;
    wire N__27400;
    wire N__27399;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27380;
    wire N__27379;
    wire N__27378;
    wire N__27377;
    wire N__27376;
    wire N__27375;
    wire N__27374;
    wire N__27373;
    wire N__27372;
    wire N__27369;
    wire N__27354;
    wire N__27353;
    wire N__27352;
    wire N__27347;
    wire N__27340;
    wire N__27337;
    wire N__27336;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27294;
    wire N__27289;
    wire N__27288;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27253;
    wire N__27252;
    wire N__27251;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27239;
    wire N__27238;
    wire N__27237;
    wire N__27236;
    wire N__27235;
    wire N__27234;
    wire N__27231;
    wire N__27230;
    wire N__27229;
    wire N__27222;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27202;
    wire N__27199;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27183;
    wire N__27180;
    wire N__27175;
    wire N__27172;
    wire N__27161;
    wire N__27156;
    wire N__27151;
    wire N__27144;
    wire N__27137;
    wire N__27116;
    wire N__27115;
    wire N__27114;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27109;
    wire N__27106;
    wire N__27105;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27097;
    wire N__27096;
    wire N__27095;
    wire N__27092;
    wire N__27087;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27060;
    wire N__27053;
    wire N__27048;
    wire N__27035;
    wire N__27034;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27023;
    wire N__27022;
    wire N__27019;
    wire N__27018;
    wire N__27017;
    wire N__27016;
    wire N__27011;
    wire N__27010;
    wire N__27009;
    wire N__27008;
    wire N__27007;
    wire N__27002;
    wire N__26999;
    wire N__26992;
    wire N__26989;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26963;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26927;
    wire N__26924;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26853;
    wire N__26852;
    wire N__26851;
    wire N__26850;
    wire N__26849;
    wire N__26848;
    wire N__26847;
    wire N__26846;
    wire N__26845;
    wire N__26844;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26840;
    wire N__26839;
    wire N__26838;
    wire N__26837;
    wire N__26836;
    wire N__26835;
    wire N__26834;
    wire N__26833;
    wire N__26832;
    wire N__26829;
    wire N__26820;
    wire N__26813;
    wire N__26812;
    wire N__26811;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26782;
    wire N__26775;
    wire N__26762;
    wire N__26757;
    wire N__26754;
    wire N__26753;
    wire N__26746;
    wire N__26743;
    wire N__26736;
    wire N__26733;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26705;
    wire N__26700;
    wire N__26695;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26665;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26643;
    wire N__26638;
    wire N__26637;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26625;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26437;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26405;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26393;
    wire N__26392;
    wire N__26389;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26363;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26326;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26314;
    wire N__26309;
    wire N__26308;
    wire N__26307;
    wire N__26304;
    wire N__26299;
    wire N__26294;
    wire N__26293;
    wire N__26290;
    wire N__26289;
    wire N__26286;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26212;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26185;
    wire N__26184;
    wire N__26183;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26177;
    wire N__26172;
    wire N__26167;
    wire N__26164;
    wire N__26163;
    wire N__26162;
    wire N__26161;
    wire N__26160;
    wire N__26159;
    wire N__26158;
    wire N__26157;
    wire N__26154;
    wire N__26149;
    wire N__26144;
    wire N__26139;
    wire N__26136;
    wire N__26131;
    wire N__26128;
    wire N__26127;
    wire N__26126;
    wire N__26117;
    wire N__26116;
    wire N__26115;
    wire N__26114;
    wire N__26113;
    wire N__26110;
    wire N__26105;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26089;
    wire N__26088;
    wire N__26085;
    wire N__26076;
    wire N__26075;
    wire N__26074;
    wire N__26073;
    wire N__26072;
    wire N__26071;
    wire N__26070;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26058;
    wire N__26055;
    wire N__26050;
    wire N__26045;
    wire N__26030;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25972;
    wire N__25967;
    wire N__25966;
    wire N__25963;
    wire N__25962;
    wire N__25961;
    wire N__25960;
    wire N__25957;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25945;
    wire N__25944;
    wire N__25943;
    wire N__25942;
    wire N__25941;
    wire N__25940;
    wire N__25939;
    wire N__25938;
    wire N__25937;
    wire N__25932;
    wire N__25927;
    wire N__25926;
    wire N__25925;
    wire N__25924;
    wire N__25923;
    wire N__25922;
    wire N__25921;
    wire N__25920;
    wire N__25917;
    wire N__25910;
    wire N__25905;
    wire N__25898;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25884;
    wire N__25883;
    wire N__25882;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25861;
    wire N__25858;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25825;
    wire N__25822;
    wire N__25811;
    wire N__25806;
    wire N__25799;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25708;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25690;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25669;
    wire N__25668;
    wire N__25665;
    wire N__25660;
    wire N__25655;
    wire N__25652;
    wire N__25651;
    wire N__25648;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25625;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25588;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25576;
    wire N__25573;
    wire N__25572;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25525;
    wire N__25520;
    wire N__25517;
    wire N__25516;
    wire N__25515;
    wire N__25508;
    wire N__25505;
    wire N__25504;
    wire N__25501;
    wire N__25500;
    wire N__25499;
    wire N__25496;
    wire N__25495;
    wire N__25490;
    wire N__25485;
    wire N__25482;
    wire N__25477;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25450;
    wire N__25449;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25399;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25357;
    wire N__25356;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25326;
    wire N__25319;
    wire N__25318;
    wire N__25317;
    wire N__25314;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25284;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25270;
    wire N__25269;
    wire N__25268;
    wire N__25267;
    wire N__25266;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25239;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25196;
    wire N__25193;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25030;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25013;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24935;
    wire N__24934;
    wire N__24929;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24862;
    wire N__24859;
    wire N__24854;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24575;
    wire N__24574;
    wire N__24573;
    wire N__24570;
    wire N__24565;
    wire N__24562;
    wire N__24557;
    wire N__24556;
    wire N__24553;
    wire N__24552;
    wire N__24547;
    wire N__24544;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24512;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24479;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24467;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24455;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24440;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24428;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24413;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24401;
    wire N__24398;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24194;
    wire N__24193;
    wire N__24192;
    wire N__24189;
    wire N__24188;
    wire N__24187;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24155;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24128;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24074;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24025;
    wire N__24022;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24010;
    wire N__24009;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23744;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23434;
    wire N__23431;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23419;
    wire N__23414;
    wire N__23413;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23236;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23219;
    wire N__23216;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23204;
    wire N__23201;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23144;
    wire N__23141;
    wire N__23140;
    wire N__23139;
    wire N__23132;
    wire N__23129;
    wire N__23128;
    wire N__23125;
    wire N__23124;
    wire N__23123;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23080;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23068;
    wire N__23067;
    wire N__23066;
    wire N__23063;
    wire N__23062;
    wire N__23059;
    wire N__23058;
    wire N__23057;
    wire N__23050;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23042;
    wire N__23041;
    wire N__23040;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23011;
    wire N__23004;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22984;
    wire N__22983;
    wire N__22982;
    wire N__22981;
    wire N__22980;
    wire N__22979;
    wire N__22978;
    wire N__22973;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22956;
    wire N__22955;
    wire N__22954;
    wire N__22953;
    wire N__22948;
    wire N__22945;
    wire N__22940;
    wire N__22937;
    wire N__22930;
    wire N__22927;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22871;
    wire N__22868;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22853;
    wire N__22850;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22838;
    wire N__22835;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22823;
    wire N__22820;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22808;
    wire N__22805;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22793;
    wire N__22790;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22715;
    wire N__22712;
    wire N__22711;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22693;
    wire N__22688;
    wire N__22685;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22670;
    wire N__22667;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22640;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22628;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22616;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22601;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22501;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22483;
    wire N__22478;
    wire N__22477;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22456;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22385;
    wire N__22384;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22348;
    wire N__22343;
    wire N__22340;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21712;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21680;
    wire N__21677;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21663;
    wire N__21658;
    wire N__21655;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21594;
    wire N__21589;
    wire N__21586;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21521;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21503;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21482;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21470;
    wire N__21469;
    wire N__21464;
    wire N__21461;
    wire N__21460;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21428;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21383;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21290;
    wire N__21289;
    wire N__21288;
    wire N__21283;
    wire N__21280;
    wire N__21275;
    wire N__21274;
    wire N__21273;
    wire N__21270;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20912;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20869;
    wire N__20868;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20797;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20758;
    wire N__20753;
    wire N__20750;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20678;
    wire N__20675;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20657;
    wire N__20656;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20644;
    wire N__20643;
    wire N__20642;
    wire N__20639;
    wire N__20638;
    wire N__20637;
    wire N__20636;
    wire N__20633;
    wire N__20632;
    wire N__20631;
    wire N__20628;
    wire N__20627;
    wire N__20624;
    wire N__20623;
    wire N__20622;
    wire N__20619;
    wire N__20612;
    wire N__20605;
    wire N__20594;
    wire N__20585;
    wire N__20582;
    wire N__20581;
    wire N__20580;
    wire N__20577;
    wire N__20576;
    wire N__20575;
    wire N__20574;
    wire N__20573;
    wire N__20570;
    wire N__20569;
    wire N__20568;
    wire N__20567;
    wire N__20566;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20552;
    wire N__20547;
    wire N__20536;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20518;
    wire N__20515;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20495;
    wire N__20492;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20396;
    wire N__20393;
    wire N__20392;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20375;
    wire N__20374;
    wire N__20371;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20359;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20330;
    wire N__20327;
    wire N__20326;
    wire N__20323;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20297;
    wire N__20296;
    wire N__20293;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20281;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20248;
    wire N__20247;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20207;
    wire N__20206;
    wire N__20203;
    wire N__20202;
    wire N__20199;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20088;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20042;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20021;
    wire N__20020;
    wire N__20019;
    wire N__20016;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19783;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19726;
    wire N__19723;
    wire N__19722;
    wire N__19719;
    wire N__19712;
    wire N__19709;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19657;
    wire N__19654;
    wire N__19649;
    wire N__19648;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19615;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19591;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19565;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19529;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19493;
    wire N__19492;
    wire N__19489;
    wire N__19488;
    wire N__19485;
    wire N__19480;
    wire N__19477;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19456;
    wire N__19453;
    wire N__19448;
    wire N__19447;
    wire N__19442;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19424;
    wire N__19423;
    wire N__19422;
    wire N__19419;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19264;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19028;
    wire N__19025;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19010;
    wire N__19007;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18995;
    wire N__18992;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18980;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18965;
    wire N__18962;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18947;
    wire N__18944;
    wire N__18943;
    wire N__18940;
    wire N__18937;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18845;
    wire N__18844;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18832;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18820;
    wire N__18815;
    wire N__18812;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18793;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18764;
    wire N__18761;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18739;
    wire N__18734;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18664;
    wire N__18659;
    wire N__18656;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18648;
    wire N__18645;
    wire N__18640;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18614;
    wire N__18613;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18584;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18569;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18533;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18459;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18443;
    wire N__18442;
    wire N__18439;
    wire N__18438;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18376;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18302;
    wire N__18299;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18287;
    wire N__18284;
    wire N__18283;
    wire N__18278;
    wire N__18275;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18267;
    wire N__18262;
    wire N__18259;
    wire N__18254;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18242;
    wire N__18241;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18220;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18203;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18188;
    wire N__18187;
    wire N__18184;
    wire N__18179;
    wire N__18176;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18151;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18125;
    wire N__18122;
    wire N__18121;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18016;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17954;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17946;
    wire N__17939;
    wire N__17936;
    wire N__17935;
    wire N__17932;
    wire N__17931;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17914;
    wire N__17911;
    wire N__17910;
    wire N__17907;
    wire N__17904;
    wire N__17901;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17870;
    wire N__17869;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17851;
    wire N__17846;
    wire N__17845;
    wire N__17844;
    wire N__17839;
    wire N__17836;
    wire N__17831;
    wire N__17830;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17818;
    wire N__17813;
    wire N__17812;
    wire N__17809;
    wire N__17808;
    wire N__17805;
    wire N__17800;
    wire N__17797;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17774;
    wire N__17771;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17756;
    wire N__17753;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17745;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17729;
    wire N__17728;
    wire N__17727;
    wire N__17724;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17710;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17692;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17673;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17657;
    wire N__17654;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17639;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17618;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17597;
    wire N__17596;
    wire N__17595;
    wire N__17592;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17473;
    wire N__17472;
    wire N__17469;
    wire N__17464;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17422;
    wire N__17419;
    wire N__17414;
    wire N__17411;
    wire N__17410;
    wire N__17407;
    wire N__17402;
    wire N__17399;
    wire N__17398;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17360;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17309;
    wire N__17308;
    wire N__17303;
    wire N__17300;
    wire N__17299;
    wire N__17296;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17278;
    wire N__17277;
    wire N__17276;
    wire N__17275;
    wire N__17272;
    wire N__17261;
    wire N__17258;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17250;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17195;
    wire N__17194;
    wire N__17193;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17179;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17153;
    wire N__17150;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17135;
    wire N__17132;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17120;
    wire N__17117;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17105;
    wire N__17102;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17087;
    wire N__17084;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17072;
    wire N__17069;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17039;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17024;
    wire N__17021;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17009;
    wire N__17006;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16994;
    wire N__16991;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16979;
    wire N__16976;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16964;
    wire N__16961;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16949;
    wire N__16946;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16931;
    wire N__16928;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16862;
    wire N__16859;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16844;
    wire N__16841;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16829;
    wire N__16826;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16753;
    wire N__16750;
    wire N__16749;
    wire N__16746;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16678;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire ICE_GPMO_2;
    wire M_CLK4;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN_net;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN_net;
    wire ICE_SYSCLK;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN_net;
    wire VCCG0;
    wire INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN_net;
    wire n25_cascade_;
    wire n27_adj_1173;
    wire n14114_cascade_;
    wire n10522_cascade_;
    wire TEST_LED;
    wire n28;
    wire n26_adj_1180;
    wire n10;
    wire DDS_MCLK1;
    wire secclk_cnt_0;
    wire bfn_3_7_0_;
    wire secclk_cnt_1;
    wire n14009;
    wire secclk_cnt_2;
    wire n14010;
    wire secclk_cnt_3;
    wire n14011;
    wire secclk_cnt_4;
    wire n14012;
    wire secclk_cnt_5;
    wire n14013;
    wire secclk_cnt_6;
    wire n14014;
    wire secclk_cnt_7;
    wire n14015;
    wire n14016;
    wire secclk_cnt_8;
    wire bfn_3_8_0_;
    wire secclk_cnt_9;
    wire n14017;
    wire secclk_cnt_10;
    wire n14018;
    wire secclk_cnt_11;
    wire n14019;
    wire n14020;
    wire secclk_cnt_13;
    wire n14021;
    wire secclk_cnt_14;
    wire n14022;
    wire secclk_cnt_15;
    wire n14023;
    wire n14024;
    wire secclk_cnt_16;
    wire bfn_3_9_0_;
    wire secclk_cnt_17;
    wire n14025;
    wire secclk_cnt_18;
    wire n14026;
    wire n14027;
    wire secclk_cnt_20;
    wire n14028;
    wire n14029;
    wire n14030;
    wire clk_16MHz;
    wire n10522;
    wire buf_adcdata2_0;
    wire cmd_rdadctmp_8_adj_1068;
    wire cmd_rdadctmp_7_adj_1069;
    wire cmd_rdadctmp_6_adj_1070;
    wire cmd_rdadctmp_5_adj_1071;
    wire cmd_rdadctmp_3_adj_1073;
    wire cmd_rdadctmp_4_adj_1072;
    wire n14_adj_1035_cascade_;
    wire M_CS2;
    wire n15165;
    wire M_MISO2;
    wire n8302_cascade_;
    wire cmd_rdadctmp_2_adj_1074;
    wire cmd_rdadctmp_0_adj_1076;
    wire cmd_rdadctmp_1_adj_1075;
    wire buf_data2_6;
    wire buf_adcdata4_7;
    wire buf_data2_7;
    wire buf_data2_4;
    wire n4304_cascade_;
    wire buf_data2_5;
    wire n4303_cascade_;
    wire n4302;
    wire n4301;
    wire buf_data2_0;
    wire buf_data2_1;
    wire buf_data2_2;
    wire n4307;
    wire n4306;
    wire n4308;
    wire buf_adcdata2_5;
    wire buf_adcdata2_6;
    wire buf_adcdata2_7;
    wire cmd_rdadctmp_15_adj_1061;
    wire buf_adcdata2_3;
    wire buf_adcdata2_4;
    wire cmd_rdadctmp_13_adj_1063;
    wire cmd_rdadctmp_14_adj_1062;
    wire cmd_rdadctmp_11_adj_1065;
    wire cmd_rdadctmp_12_adj_1064;
    wire buf_adcdata1_5;
    wire buf_adcdata1_7;
    wire buf_adcdata4_5;
    wire cmd_rdadctmp_13_adj_1136;
    wire cmd_rdadctmp_14_adj_1135;
    wire buf_adcdata4_6;
    wire cmd_rdadctmp_15_adj_1134;
    wire buf_adcdata4_0;
    wire buf_adcdata4_1;
    wire cmd_rdadctmp_9_adj_1140;
    wire cmd_rdadctmp_10_adj_1139;
    wire buf_adcdata4_2;
    wire cmd_rdadctmp_7_adj_1142;
    wire cmd_rdadctmp_8_adj_1141;
    wire cmd_rdadctmp_5_adj_1144;
    wire cmd_rdadctmp_6_adj_1143;
    wire cmd_rdadctmp_11_adj_1138;
    wire cmd_rdadctmp_4_adj_1145;
    wire cmd_rdadctmp_3_adj_1146;
    wire cmd_rdadctmp_2_adj_1147;
    wire cmd_rdadctmp_12_adj_1137;
    wire buf_adcdata4_4;
    wire buf_data1_6;
    wire n4146;
    wire buf_data1_0;
    wire buf_data1_7;
    wire n4145;
    wire n4152;
    wire n15131_cascade_;
    wire n8738_cascade_;
    wire n8847;
    wire n8847_cascade_;
    wire n10611;
    wire n8787_cascade_;
    wire buf_data1_2;
    wire n4150_cascade_;
    wire buf_data1_4;
    wire n4148_cascade_;
    wire buf_data1_5;
    wire n4147_cascade_;
    wire n8738;
    wire n10590;
    wire secclk_cnt_21;
    wire secclk_cnt_19;
    wire secclk_cnt_12;
    wire secclk_cnt_22;
    wire n14_adj_1163;
    wire buf_data2_10;
    wire n4062_cascade_;
    wire buf_adcdata3_2;
    wire cmd_rdadctmp_11_adj_1101;
    wire buf_adcdata1_3;
    wire buf_adcdata3_4;
    wire cmd_rdadctmp_1;
    wire buf_adcdata3_7;
    wire M_MISO1;
    wire cmd_rdadctmp_0;
    wire cmd_rdadctmp_12_adj_1100;
    wire buf_adcdata1_4;
    wire cmd_rdadctmp_2;
    wire cmd_rdadctmp_7;
    wire cmd_rdadctmp_6;
    wire cmd_rdadctmp_5;
    wire cmd_rdadctmp_3;
    wire cmd_rdadctmp_4;
    wire n15168;
    wire n15168_cascade_;
    wire M_CS1;
    wire n14_adj_1039;
    wire M_SCLK1;
    wire \ADC_VAC1.n9312_cascade_ ;
    wire \ADC_VAC1.n15338_cascade_ ;
    wire \ADC_VAC1.n15360_cascade_ ;
    wire \ADC_VAC1.bit_cnt_0 ;
    wire bfn_6_16_0_;
    wire \ADC_VAC1.bit_cnt_1 ;
    wire \ADC_VAC1.n13981 ;
    wire \ADC_VAC1.bit_cnt_2 ;
    wire \ADC_VAC1.n13982 ;
    wire \ADC_VAC1.bit_cnt_3 ;
    wire \ADC_VAC1.n13983 ;
    wire \ADC_VAC1.bit_cnt_4 ;
    wire \ADC_VAC1.n13984 ;
    wire \ADC_VAC1.bit_cnt_5 ;
    wire \ADC_VAC1.n13985 ;
    wire \ADC_VAC1.bit_cnt_6 ;
    wire \ADC_VAC1.n13986 ;
    wire \ADC_VAC1.n13987 ;
    wire \ADC_VAC1.bit_cnt_7 ;
    wire \ADC_VAC1.n9312 ;
    wire \ADC_VAC1.n10667 ;
    wire n16470_cascade_;
    wire comm_buf_5_5;
    wire comm_buf_2_5;
    wire n16416_cascade_;
    wire n16473;
    wire n16419_cascade_;
    wire n7_adj_1238_cascade_;
    wire buf_data2_21;
    wire n4103_cascade_;
    wire comm_buf_3_5;
    wire buf_data2_17;
    wire n4107_cascade_;
    wire buf_data2_18;
    wire n8787;
    wire n10599;
    wire comm_buf_2_2;
    wire n15388_cascade_;
    wire n16389_cascade_;
    wire comm_buf_4_2;
    wire comm_buf_5_2;
    wire n15448;
    wire n15447_cascade_;
    wire n16386;
    wire buf_adcdata4_18;
    wire comm_buf_2_3;
    wire comm_buf_4_3;
    wire comm_buf_5_3;
    wire n16440_cascade_;
    wire n15423;
    wire n15397;
    wire n16392_cascade_;
    wire n16443;
    wire n16395_cascade_;
    wire M_SCLK2;
    wire buf_adcdata3_5;
    wire buf_adcdata3_6;
    wire cmd_rdadctmp_12;
    wire cmd_rdadctmp_10_adj_1102;
    wire cmd_rdadctmp_16_adj_1133;
    wire cmd_rdadctmp_17_adj_1132;
    wire cmd_rdadctmp_18_adj_1131;
    wire buf_adcdata4_10;
    wire \ADC_VAC1.n15263_cascade_ ;
    wire \ADC_VAC1.n15553 ;
    wire \ADC_VAC1.n15264 ;
    wire M_DRDY1;
    wire \ADC_VAC1.n17_cascade_ ;
    wire \ADC_VAC1.n12 ;
    wire cmd_rdadctmp_13;
    wire cmd_rdadctmp_1_adj_1148;
    wire M_MISO4;
    wire cmd_rdadctmp_0_adj_1149;
    wire cmd_rdadctmp_15;
    wire M_START;
    wire comm_buf_3_0;
    wire comm_buf_2_0;
    wire n16413_cascade_;
    wire comm_buf_5_6;
    wire n16518_cascade_;
    wire n13493;
    wire n16521_cascade_;
    wire comm_buf_2_6;
    wire comm_buf_3_6;
    wire n16410;
    wire n16491;
    wire comm_buf_2_1;
    wire comm_buf_3_1;
    wire n16404_cascade_;
    wire n16407_cascade_;
    wire comm_buf_5_1;
    wire comm_buf_4_1;
    wire n16515;
    wire n16512;
    wire n7_adj_1240;
    wire n16425_cascade_;
    wire buf_data2_12;
    wire n4060_cascade_;
    wire comm_buf_4_5;
    wire comm_buf_4_6;
    wire buf_data2_15;
    wire n4057_cascade_;
    wire n10604;
    wire buf_adcdata1_17;
    wire buf_adcdata1_18;
    wire cmd_rdadctmp_26;
    wire cmd_rdadctmp_27;
    wire buf_adcdata1_19;
    wire cmd_rdadctmp_25;
    wire buf_adcdata1_20;
    wire n84_cascade_;
    wire n15593_cascade_;
    wire n8045_cascade_;
    wire n15573;
    wire cmd_rdadctmp_11;
    wire buf_adcdata4_12;
    wire cmd_rdadctmp_16_adj_1060;
    wire buf_adcdata2_8;
    wire cmd_rdadctmp_9_adj_1103;
    wire cmd_rdadctmp_28;
    wire buf_adcdata2_17;
    wire cmd_rdadctmp_13_adj_1099;
    wire cmd_rdadctmp_14_adj_1098;
    wire buf_data2_14;
    wire n4058;
    wire n14_adj_1031_cascade_;
    wire M_CS3;
    wire M_SCLK3;
    wire cmd_rdadctmp_4_adj_1108;
    wire DTRIG_N_957;
    wire adc_state_1;
    wire M_MISO3;
    wire cmd_rdadctmp_0_adj_1112;
    wire cmd_rdadctmp_1_adj_1111;
    wire \ADC_VAC3.n12 ;
    wire n15162;
    wire n15162_cascade_;
    wire \comm_spi.n16911 ;
    wire \comm_spi.n10433 ;
    wire \comm_spi.n16911_cascade_ ;
    wire \comm_spi.data_tx_7__N_811 ;
    wire \comm_spi.data_tx_7__N_831 ;
    wire \comm_spi.data_tx_7__N_812 ;
    wire comm_tx_buf_1;
    wire n15411;
    wire n16446_cascade_;
    wire n15391;
    wire n16449;
    wire buf_data2_3;
    wire buf_adcdata4_3;
    wire n4305;
    wire n16431;
    wire comm_buf_4_0;
    wire n16506_cascade_;
    wire comm_buf_5_0;
    wire n16509;
    wire n15424;
    wire n15412;
    wire comm_buf_5_7;
    wire comm_buf_4_7;
    wire n16482_cascade_;
    wire n16485;
    wire \INVcomm_spi.imiso_83_7340_7341_resetC_net ;
    wire comm_buf_3_7_N_501_2;
    wire comm_buf_3_2;
    wire comm_buf_3_3;
    wire buf_data4_19;
    wire comm_buf_9_3;
    wire buf_data4_20;
    wire n66_adj_1153_cascade_;
    wire DDS_SCK1;
    wire DDS_MOSI1;
    wire n15522;
    wire n15523;
    wire n16398_cascade_;
    wire n16401_cascade_;
    wire n109_adj_1155_cascade_;
    wire n8048_cascade_;
    wire n15578;
    wire buf_adcdata1_21;
    wire buf_adcdata1_22;
    wire cmd_rdadctmp_24_adj_1052;
    wire buf_adcdata2_16;
    wire cmd_rdadctmp_29;
    wire cmd_rdadctmp_30;
    wire buf_adcdata1_1;
    wire bfn_9_13_0_;
    wire \ADC_VAC2.n13988 ;
    wire \ADC_VAC2.n13989 ;
    wire \ADC_VAC2.n13990 ;
    wire \ADC_VAC2.n13991 ;
    wire \ADC_VAC2.n13992 ;
    wire \ADC_VAC2.n13993 ;
    wire \ADC_VAC2.n13994 ;
    wire \ADC_VAC2.bit_cnt_1 ;
    wire \ADC_VAC2.bit_cnt_7 ;
    wire \ADC_VAC2.n15261_cascade_ ;
    wire \ADC_VAC2.n15595 ;
    wire \ADC_VAC2.n15262 ;
    wire \ADC_VAC2.bit_cnt_6 ;
    wire \ADC_VAC2.bit_cnt_0 ;
    wire \ADC_VAC2.n16 ;
    wire \ADC_VAC2.n17_cascade_ ;
    wire cmd_rdadctmp_2_adj_1110;
    wire cmd_rdadctmp_3_adj_1109;
    wire acadc_dtrig2;
    wire acadc_dtrig1;
    wire acadc_dtrig4;
    wire acadc_dtrig3;
    wire cmd_rdadctmp_14;
    wire buf_adcdata1_6;
    wire cmd_rdadctmp_15_adj_1097;
    wire M_SCLK4;
    wire \comm_spi.n10434 ;
    wire comm_tx_buf_0;
    wire \comm_spi.data_tx_7__N_834 ;
    wire n16428;
    wire buf_data2_20;
    wire n4104;
    wire comm_buf_3_7;
    wire comm_buf_2_7;
    wire n15382_cascade_;
    wire n16383_cascade_;
    wire n16494_cascade_;
    wire n16497;
    wire n15450;
    wire n15451_cascade_;
    wire n16380;
    wire buf_data4_1;
    wire buf_data4_2;
    wire comm_buf_11_2;
    wire buf_data4_3;
    wire comm_buf_11_3;
    wire buf_data4_4;
    wire buf_data4_5;
    wire comm_buf_11_5;
    wire buf_data4_6;
    wire buf_data4_7;
    wire comm_buf_11_7;
    wire buf_data4_0;
    wire comm_buf_11_0;
    wire buf_data3_15;
    wire comm_buf_7_7;
    wire buf_data3_8;
    wire comm_buf_7_0;
    wire buf_data3_14;
    wire comm_buf_7_6;
    wire buf_data3_13;
    wire comm_buf_7_5;
    wire buf_data3_12;
    wire buf_data3_11;
    wire comm_buf_7_3;
    wire buf_data3_10;
    wire comm_buf_7_2;
    wire buf_data3_9;
    wire comm_buf_7_1;
    wire comm_buf_3_4;
    wire comm_buf_2_4;
    wire n15403_cascade_;
    wire n16479_cascade_;
    wire n10660;
    wire comm_buf_7_4;
    wire comm_buf_11_4;
    wire comm_buf_9_4;
    wire n16452_cascade_;
    wire n16455;
    wire comm_buf_5_4;
    wire comm_buf_4_4;
    wire n15400;
    wire n15399_cascade_;
    wire n16476;
    wire n15633_cascade_;
    wire n16458_cascade_;
    wire n16461_cascade_;
    wire n76_cascade_;
    wire n4_adj_1195_cascade_;
    wire n15632;
    wire n15589;
    wire n87_adj_1165_cascade_;
    wire n69_adj_1161_cascade_;
    wire n130;
    wire n8050;
    wire n8089;
    wire n96_adj_1159;
    wire n130_adj_1156_cascade_;
    wire n15587;
    wire n8051_cascade_;
    wire cmd_rdadctmp_19_adj_1130;
    wire cmd_rdadctmp_8;
    wire buf_adcdata1_0;
    wire cmd_rdadctmp_23;
    wire buf_adcdata1_15;
    wire cmd_rdadctmp_20_adj_1129;
    wire \ADC_VAC2.bit_cnt_4 ;
    wire \ADC_VAC2.bit_cnt_3 ;
    wire \ADC_VAC2.bit_cnt_5 ;
    wire \ADC_VAC2.bit_cnt_2 ;
    wire \ADC_VAC2.n15596 ;
    wire \ADC_VAC3.n15334_cascade_ ;
    wire \ADC_VAC3.n15358_cascade_ ;
    wire \ADC_VAC3.n15602_cascade_ ;
    wire \ADC_VAC3.n15260 ;
    wire \ADC_VAC3.n15259 ;
    wire \ADC_VAC3.n17 ;
    wire \ADC_VAC3.bit_cnt_0 ;
    wire bfn_10_15_0_;
    wire \ADC_VAC3.bit_cnt_1 ;
    wire \ADC_VAC3.n13995 ;
    wire \ADC_VAC3.bit_cnt_2 ;
    wire \ADC_VAC3.n13996 ;
    wire \ADC_VAC3.bit_cnt_3 ;
    wire \ADC_VAC3.n13997 ;
    wire \ADC_VAC3.bit_cnt_4 ;
    wire \ADC_VAC3.n13998 ;
    wire \ADC_VAC3.bit_cnt_5 ;
    wire \ADC_VAC3.n13999 ;
    wire \ADC_VAC3.bit_cnt_6 ;
    wire \ADC_VAC3.n14000 ;
    wire \ADC_VAC3.n14001 ;
    wire \ADC_VAC3.bit_cnt_7 ;
    wire cmd_rdadctmp_31;
    wire buf_adcdata1_23;
    wire M_DRDY3;
    wire adc_state_1_adj_1079;
    wire \ADC_VAC3.n9514 ;
    wire DTRIG_N_957_adj_1114;
    wire \ADC_VAC3.n9514_cascade_ ;
    wire \ADC_VAC3.n10744 ;
    wire bfn_10_17_0_;
    wire \ADC_VAC4.n14002 ;
    wire \ADC_VAC4.n14003 ;
    wire \ADC_VAC4.n14004 ;
    wire \ADC_VAC4.n14005 ;
    wire \ADC_VAC4.n14006 ;
    wire \ADC_VAC4.n14007 ;
    wire \ADC_VAC4.n14008 ;
    wire \comm_spi.n16908 ;
    wire \comm_spi.n10459 ;
    wire \comm_spi.n10460 ;
    wire \comm_spi.data_tx_7__N_828 ;
    wire buf_adcdata4_21;
    wire cmd_rdadctmp_29_adj_1120;
    wire cmd_rdadctmp_30_adj_1119;
    wire cmd_rdadctmp_31_adj_1118;
    wire buf_data3_7;
    wire comm_buf_8_7;
    wire buf_data3_6;
    wire comm_buf_8_6;
    wire buf_data3_5;
    wire comm_buf_8_5;
    wire buf_data3_4;
    wire comm_buf_8_4;
    wire buf_data3_3;
    wire comm_buf_8_3;
    wire buf_data3_2;
    wire comm_buf_8_2;
    wire buf_data3_1;
    wire comm_buf_8_1;
    wire buf_data3_0;
    wire comm_buf_8_0;
    wire buf_data3_23;
    wire comm_buf_6_7;
    wire buf_data3_22;
    wire comm_buf_6_6;
    wire buf_data3_21;
    wire comm_buf_6_5;
    wire buf_data3_20;
    wire comm_buf_6_4;
    wire buf_data3_19;
    wire comm_buf_6_3;
    wire buf_data3_18;
    wire comm_buf_6_2;
    wire n8907_cascade_;
    wire n8943;
    wire n8943_cascade_;
    wire n10625;
    wire n9123;
    wire n9123_cascade_;
    wire n10653;
    wire buf_data3_16;
    wire comm_buf_6_0;
    wire buf_data3_17;
    wire comm_buf_6_1;
    wire n8907;
    wire n10618;
    wire buf_data4_10;
    wire comm_buf_10_2;
    wire buf_data4_11;
    wire comm_buf_10_3;
    wire buf_data4_12;
    wire comm_buf_10_4;
    wire buf_data4_15;
    wire comm_buf_10_7;
    wire buf_data4_8;
    wire comm_buf_10_0;
    wire n16434_cascade_;
    wire n16437_cascade_;
    wire n109;
    wire n8054_cascade_;
    wire n59;
    wire cmd_rdadctmp_25_adj_1087;
    wire cmd_rdadctmp_7_adj_1105;
    wire n16500_cascade_;
    wire n16503_cascade_;
    wire n4_adj_1280;
    wire n8047_cascade_;
    wire n10576;
    wire cmd_rdadctmp_9;
    wire buf_control_3;
    wire n69_adj_1029;
    wire buf_adcdata4_14;
    wire buf_adcdata3_20;
    wire n61;
    wire buf_control_4;
    wire n69;
    wire buf_control_0;
    wire buf_data2_8;
    wire buf_adcdata4_8;
    wire n4064;
    wire cmd_rdadctmp_5_adj_1107;
    wire cmd_rdadctmp_6_adj_1106;
    wire cmd_rdadctmp_28_adj_1084;
    wire buf_adcdata1_9;
    wire cmd_rdadctmp_17;
    wire cmd_rdadctmp_19;
    wire buf_adcdata1_11;
    wire buf_adcdata3_8;
    wire \ADC_VAC4.bit_cnt_4 ;
    wire \ADC_VAC4.bit_cnt_3 ;
    wire \ADC_VAC4.bit_cnt_1 ;
    wire \ADC_VAC4.bit_cnt_2 ;
    wire \ADC_VAC4.bit_cnt_6 ;
    wire \ADC_VAC4.bit_cnt_0 ;
    wire \ADC_VAC4.n15330_cascade_ ;
    wire \ADC_VAC4.bit_cnt_7 ;
    wire \ADC_VAC4.bit_cnt_5 ;
    wire \ADC_VAC4.n15354 ;
    wire \ADC_VAC4.n15619_cascade_ ;
    wire \ADC_VAC4.n9631 ;
    wire \ADC_VAC4.n9631_cascade_ ;
    wire \ADC_VAC4.n10783 ;
    wire buf_adcdata4_20;
    wire \comm_spi.n16905_cascade_ ;
    wire \comm_spi.data_tx_7__N_809 ;
    wire comm_tx_buf_2;
    wire \comm_spi.data_tx_7__N_810 ;
    wire \comm_spi.n16905 ;
    wire \comm_spi.n10463 ;
    wire \comm_spi.n10464 ;
    wire buf_data4_21;
    wire comm_buf_9_5;
    wire buf_data4_22;
    wire comm_buf_9_6;
    wire buf_data4_23;
    wire comm_buf_9_7;
    wire buf_data4_18;
    wire comm_buf_9_2;
    wire buf_data4_17;
    wire comm_buf_9_1;
    wire n15161_cascade_;
    wire n8997;
    wire n8997_cascade_;
    wire n10632;
    wire buf_data4_16;
    wire comm_buf_9_0;
    wire n9027;
    wire n10639;
    wire comm_buf_11_1;
    wire n16422;
    wire buf_data4_9;
    wire comm_buf_10_1;
    wire n8763;
    wire n13470;
    wire n13497;
    wire n13497_cascade_;
    wire n9045_cascade_;
    wire comm_buf_11_6;
    wire n16488;
    wire buf_data4_14;
    wire comm_buf_10_6;
    wire n13457_cascade_;
    wire n15565_cascade_;
    wire n13_adj_1257_cascade_;
    wire n8823;
    wire n41;
    wire n13457;
    wire n13458;
    wire buf_data4_13;
    wire comm_buf_10_5;
    wire n9045;
    wire n10646;
    wire n11_adj_1279_cascade_;
    wire n8654;
    wire n5;
    wire n15221;
    wire n17_cascade_;
    wire n8702_cascade_;
    wire bit_cnt_3;
    wire bit_cnt_2;
    wire bit_cnt_0;
    wire n16524_cascade_;
    wire n16527_cascade_;
    wire n4_adj_1264_cascade_;
    wire n8055;
    wire buf_adcdata4_15;
    wire n15144;
    wire buf_adcdata4_17;
    wire n71;
    wire cmd_rdadctmp_26_adj_1123;
    wire cmd_rdadctmp_27_adj_1085;
    wire buf_adcdata3_23;
    wire cmd_rdadctmp_27_adj_1122;
    wire cmd_rdadctmp_28_adj_1121;
    wire cmd_rdadctmp_23_adj_1126;
    wire cmd_rdadctmp_24_adj_1125;
    wire cmd_rdadctmp_25_adj_1124;
    wire M_POW;
    wire buf_adcdata3_19;
    wire n87;
    wire n8272;
    wire cmd_rdadctmp_26_adj_1086;
    wire buf_adcdata3_18;
    wire n15811;
    wire cmd_rdadctmp_21_adj_1128;
    wire cmd_rdadctmp_22_adj_1127;
    wire buf_adcdata3_16;
    wire n90;
    wire n15156_cascade_;
    wire n9694;
    wire \ADC_VAC4.n15257_cascade_ ;
    wire \ADC_VAC4.n15258 ;
    wire \ADC_VAC4.n15278 ;
    wire M_DRDY4;
    wire n14_cascade_;
    wire n15156;
    wire M_CS4;
    wire buf_data2_11;
    wire buf_adcdata4_11;
    wire n4061;
    wire \ADC_VAC4.n17 ;
    wire adc_state_0_adj_1117;
    wire DTRIG_N_957_adj_1150;
    wire adc_state_1_adj_1116;
    wire \ADC_VAC4.n12 ;
    wire \ADC_VAC4.n14930 ;
    wire \comm_spi.n10467 ;
    wire \comm_spi.n10468 ;
    wire \comm_spi.data_tx_7__N_822 ;
    wire DDS_CS1;
    wire comm_tx_buf_7;
    wire comm_tx_buf_6;
    wire \comm_spi.n16884 ;
    wire buf_data1_23;
    wire n18_cascade_;
    wire n15466_cascade_;
    wire n104;
    wire n56;
    wire buf_adcdata3_1;
    wire buf_data1_1;
    wire n4151;
    wire n15567_cascade_;
    wire n7_adj_1255;
    wire n6;
    wire n5_adj_1235_cascade_;
    wire n15535_cascade_;
    wire n15_cascade_;
    wire n9021;
    wire n4814;
    wire n4814_cascade_;
    wire n5_adj_1235;
    wire n13475_cascade_;
    wire n15802_cascade_;
    wire n10_adj_1249;
    wire n15657_cascade_;
    wire n13_adj_1042;
    wire \comm_spi.n10479 ;
    wire \comm_spi.data_tx_7__N_806 ;
    wire n15576;
    wire n15691;
    wire n15475;
    wire n15835;
    wire n15542;
    wire n15679;
    wire n15543;
    wire buf_adcdata3_17;
    wire M_DCSEL;
    wire n90_adj_1023_cascade_;
    wire n69_adj_1113;
    wire n96;
    wire buf_device_acadc_4;
    wire M_OSR0;
    wire n15555;
    wire n3_cascade_;
    wire n10_adj_1242_cascade_;
    wire n8_adj_1212;
    wire eis_end;
    wire INVeis_end_328C_net;
    wire n15171_cascade_;
    wire raw_buf1_N_775;
    wire n14087;
    wire n15356_cascade_;
    wire n15695_cascade_;
    wire n15696;
    wire n15700_cascade_;
    wire n3;
    wire INVeis_state_i0C_net;
    wire n8459;
    wire data_index_9_N_258_4;
    wire eis_end_N_773;
    wire eis_end_N_773_cascade_;
    wire n15510;
    wire n8_adj_1227;
    wire cmd_rdadctmp_24_adj_1088;
    wire data_index_9_N_258_1;
    wire buf_data2_13;
    wire buf_adcdata4_13;
    wire n4059;
    wire n8_adj_1233;
    wire n8_adj_1233_cascade_;
    wire M_FLT0;
    wire n66_adj_1166;
    wire bfn_13_16_0_;
    wire INVacadc_skipcnt_i0_i0C_net;
    wire n13966;
    wire n13966_THRU_CRY_0_THRU_CO;
    wire n13966_THRU_CRY_1_THRU_CO;
    wire n13966_THRU_CRY_2_THRU_CO;
    wire n13966_THRU_CRY_3_THRU_CO;
    wire n13966_THRU_CRY_4_THRU_CO;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire n13966_THRU_CRY_5_THRU_CO;
    wire n13966_THRU_CRY_6_THRU_CO;
    wire acadc_skipcnt_1;
    wire bfn_13_17_0_;
    wire n13967;
    wire n13968;
    wire acadc_skipcnt_4;
    wire n13969;
    wire n13970;
    wire n13971;
    wire n13972;
    wire n13973;
    wire n13974;
    wire INVacadc_skipcnt_i0_i1C_net;
    wire bfn_13_18_0_;
    wire n13975;
    wire n13976;
    wire n13977;
    wire n13978;
    wire n13979;
    wire n13980;
    wire INVacadc_skipcnt_i0_i9C_net;
    wire buf_data2_22;
    wire buf_adcdata4_22;
    wire n4102;
    wire \comm_spi.n16902 ;
    wire \comm_spi.n10476 ;
    wire \comm_spi.n10480 ;
    wire \comm_spi.data_tx_7__N_816 ;
    wire \comm_spi.n10472 ;
    wire \comm_spi.n10471 ;
    wire \comm_spi.n10475 ;
    wire \comm_spi.data_tx_7__N_807 ;
    wire \comm_spi.n16896 ;
    wire n15474;
    wire n15478;
    wire n15680;
    wire \INVcomm_spi.data_valid_85C_net ;
    wire \comm_spi.n10449 ;
    wire \comm_spi.n10448 ;
    wire \INVcomm_spi.imiso_83_7340_7341_setC_net ;
    wire n15387;
    wire n15390;
    wire \CLOCK_DDS.tmp_buf_10 ;
    wire \CLOCK_DDS.tmp_buf_11 ;
    wire \CLOCK_DDS.tmp_buf_12 ;
    wire \CLOCK_DDS.tmp_buf_13 ;
    wire \CLOCK_DDS.tmp_buf_14 ;
    wire buf_dds_9;
    wire \CLOCK_DDS.tmp_buf_9 ;
    wire \CLOCK_DDS.tmp_buf_8 ;
    wire n4260_cascade_;
    wire n15402;
    wire ICE_CHKCABLE;
    wire n90_adj_1154_cascade_;
    wire n72;
    wire M_OSR1;
    wire n15479;
    wire cmd_rdadctmp_31_adj_1081;
    wire n8_adj_1221_cascade_;
    wire n4205;
    wire buf_device_acadc_7;
    wire buf_dds_14;
    wire n4219;
    wire req_data_cnt_15;
    wire req_data_cnt_9;
    wire n22;
    wire n24_adj_1216_cascade_;
    wire n30_adj_1278;
    wire n6791_cascade_;
    wire n8_adj_1178_cascade_;
    wire n7_adj_1177;
    wire n7_adj_1177_cascade_;
    wire n8_adj_1178;
    wire data_index_9_N_258_0;
    wire acadc_skipcnt_0;
    wire acadc_skipcnt_6;
    wire n18_adj_1276;
    wire n17_adj_1277_cascade_;
    wire n31;
    wire n31_cascade_;
    wire n15187;
    wire n8_adj_1231;
    wire data_index_9_N_258_2;
    wire M_FLT1;
    wire acadc_skipcnt_14;
    wire acadc_skipcnt_11;
    wire acadc_skipCount_11;
    wire n23_adj_1199_cascade_;
    wire n30;
    wire acadc_skipcnt_10;
    wire acadc_skipCount_12;
    wire acadc_skipcnt_12;
    wire n21;
    wire data_index_0;
    wire data_index_9_N_647_0;
    wire bfn_14_16_0_;
    wire data_index_1;
    wire n7_adj_1232;
    wire n14031;
    wire data_index_2;
    wire n7_adj_1230;
    wire n14032;
    wire n14033;
    wire data_index_4;
    wire n7_adj_1226;
    wire n14034;
    wire n14035;
    wire n14036;
    wire data_index_7;
    wire n14037;
    wire n14038;
    wire bfn_14_17_0_;
    wire data_index_3;
    wire M_DRDY2;
    wire n10532;
    wire n15344;
    wire n15171;
    wire n15328_cascade_;
    wire acadc_trig;
    wire INVacadc_trig_329C_net;
    wire data_index_6;
    wire n8_adj_1221;
    wire n7_adj_1220;
    wire data_index_9_N_258_7;
    wire n7_adj_1222;
    wire n8_adj_1223;
    wire data_index_9_N_258_6;
    wire ICE_SPI_MISO;
    wire \comm_spi.n10446 ;
    wire \INVcomm_spi.MISO_48_7334_7335_resetC_net ;
    wire \comm_spi.data_tx_7__N_813 ;
    wire comm_tx_buf_3;
    wire \comm_spi.data_tx_7__N_825 ;
    wire buf_data1_22;
    wire n66;
    wire \comm_spi.n10452 ;
    wire \comm_spi.n10451 ;
    wire \comm_spi.n10444 ;
    wire \comm_spi.n10445 ;
    wire \INVcomm_spi.MISO_48_7334_7335_setC_net ;
    wire \comm_spi.data_tx_7__N_805 ;
    wire n10640;
    wire n15176;
    wire n15396;
    wire n15670;
    wire n13475;
    wire n15_adj_1203;
    wire tmp_buf_15;
    wire \CLOCK_DDS.tmp_buf_0 ;
    wire \CLOCK_DDS.tmp_buf_1 ;
    wire \CLOCK_DDS.tmp_buf_2 ;
    wire \CLOCK_DDS.tmp_buf_3 ;
    wire \CLOCK_DDS.tmp_buf_4 ;
    wire \CLOCK_DDS.tmp_buf_5 ;
    wire \CLOCK_DDS.tmp_buf_6 ;
    wire \CLOCK_DDS.tmp_buf_7 ;
    wire \CLOCK_DDS.n9759 ;
    wire n10823;
    wire \CLOCK_DDS.n9_adj_1021 ;
    wire bit_cnt_1;
    wire n15556;
    wire n60_adj_1157;
    wire n4252;
    wire n4202;
    wire n4247;
    wire buf_dds_15;
    wire req_data_cnt_13;
    wire req_data_cnt_8;
    wire n15812;
    wire buf_device_acadc_6;
    wire buf_data1_16;
    wire n99;
    wire req_data_cnt_7;
    wire n4214;
    wire buf_dds_7;
    wire n7567;
    wire n21_adj_1204;
    wire comm_buf_1_4;
    wire buf_dds_4;
    wire buf_control_5;
    wire buf_data1_10;
    wire n4195_cascade_;
    wire n4232;
    wire acadc_skipcnt_9;
    wire acadc_skipcnt_15;
    wire n24_adj_1174;
    wire req_data_cnt_14;
    wire n23_adj_1194;
    wire acadc_skipCount_4;
    wire n9224;
    wire buf_device_acadc_5;
    wire acadc_skipCount_9;
    wire n15834;
    wire n19_adj_1234;
    wire n20_adj_1253_cascade_;
    wire n29;
    wire n84;
    wire n15546;
    wire data_index_5;
    wire buf_dds_12;
    wire acadc_skipcnt_2;
    wire acadc_skipCount_7;
    wire acadc_skipcnt_7;
    wire acadc_skipCount_2;
    wire n22_adj_1170;
    wire n8_adj_1229;
    wire n7_adj_1228;
    wire data_index_9_N_258_3;
    wire n8456;
    wire acadc_skipcnt_3;
    wire acadc_skipcnt_5;
    wire acadc_skipcnt_8;
    wire acadc_skipCount_8;
    wire n20_cascade_;
    wire n26;
    wire acadc_skipcnt_13;
    wire acadc_skipCount_13;
    wire n14_adj_1160;
    wire cmd_rdadctmp_16;
    wire buf_adcdata1_8;
    wire eis_state_0;
    wire eis_end_N_770;
    wire ICE_GPMO_0;
    wire data_index_8;
    wire buf_data1_3;
    wire buf_adcdata3_3;
    wire n4149;
    wire comm_tx_buf_5;
    wire \comm_spi.data_tx_7__N_819 ;
    wire n8561;
    wire n15460_cascade_;
    wire n19_cascade_;
    wire n15463;
    wire n23;
    wire n19_adj_1151_cascade_;
    wire comm_length_2;
    wire comm_index_2;
    wire comm_length_3;
    wire comm_index_3;
    wire n6_adj_1281_cascade_;
    wire comm_index_1;
    wire n2;
    wire n15119_cascade_;
    wire comm_length_1;
    wire n13_cascade_;
    wire n6_adj_1273;
    wire n5_adj_1282;
    wire comm_length_0;
    wire n10566;
    wire n13;
    wire n12649;
    wire n8525_cascade_;
    wire n4075;
    wire n8133;
    wire trig_dds;
    wire buf_dds_0;
    wire buf_dds_8;
    wire buf_data1_15;
    wire n4190_cascade_;
    wire n4227;
    wire n4262;
    wire comm_buf_0_5;
    wire n14_adj_1202_cascade_;
    wire buf_dds_13;
    wire n15690;
    wire req_data_cnt_12;
    wire n13_adj_1026;
    wire buf_data1_17;
    wire n78_cascade_;
    wire n99_adj_1024;
    wire n4257;
    wire comm_buf_1_6;
    wire buf_data1_21;
    wire n66_adj_1158;
    wire buf_dds_5;
    wire acadc_skipCount_10;
    wire n7485_cascade_;
    wire tacadc_rst;
    wire req_data_cnt_10;
    wire n90_adj_1167;
    wire n72_adj_1162;
    wire comm_buf_0_0;
    wire req_data_cnt_4;
    wire n18_adj_1217;
    wire buf_dds_6;
    wire comm_buf_0_1;
    wire n7485;
    wire eis_stop;
    wire cmd_rdadctmp_23_adj_1053;
    wire buf_adcdata2_15;
    wire comm_buf_0_2;
    wire buf_dds_10;
    wire acadc_skipCount_0;
    wire n17_adj_1214;
    wire req_data_cnt_0;
    wire acadc_skipCount_6;
    wire buf_data1_14;
    wire n4191_cascade_;
    wire n4215;
    wire n4228_cascade_;
    wire n4203;
    wire n4248_cascade_;
    wire n4258;
    wire bfn_16_16_0_;
    wire n13951;
    wire data_cntvec_2;
    wire n13952;
    wire n13953;
    wire n13954;
    wire n13955;
    wire data_cntvec_6;
    wire n13956;
    wire data_cntvec_7;
    wire n13957;
    wire n13958;
    wire INVdata_cntvec_i0_i0C_net;
    wire data_cntvec_8;
    wire bfn_16_17_0_;
    wire data_cntvec_9;
    wire n13959;
    wire data_cntvec_10;
    wire n13960;
    wire data_cntvec_11;
    wire n13961;
    wire data_cntvec_12;
    wire n13962;
    wire data_cntvec_13;
    wire n13963;
    wire data_cntvec_14;
    wire n13964;
    wire n13965;
    wire data_cntvec_15;
    wire INVdata_cntvec_i0_i8C_net;
    wire data_count_0;
    wire bfn_16_18_0_;
    wire data_count_1;
    wire n13942;
    wire data_count_2;
    wire n13943;
    wire data_count_3;
    wire n13944;
    wire data_count_4;
    wire n13945;
    wire data_count_5;
    wire n13946;
    wire data_count_6;
    wire n13947;
    wire data_count_7;
    wire n13948;
    wire n13949;
    wire INVdata_count_i0_i0C_net;
    wire bfn_16_19_0_;
    wire data_count_8;
    wire INVdata_count_i0_i8C_net;
    wire dds_state_2;
    wire \ADC_VAC2.n15280 ;
    wire adc_state_1_adj_1043;
    wire \ADC_VAC2.n12 ;
    wire \ADC_VAC2.n14926 ;
    wire \ADC_VAC2.n9413 ;
    wire DTRIG_N_957_adj_1077;
    wire \ADC_VAC2.n10706 ;
    wire \comm_spi.bit_cnt_2 ;
    wire \comm_spi.bit_cnt_1 ;
    wire \comm_spi.bit_cnt_0 ;
    wire \INVcomm_spi.bit_cnt_1603__i3C_net ;
    wire n15668_cascade_;
    wire n1523;
    wire n1523_cascade_;
    wire n2_adj_1200_cascade_;
    wire n16464;
    wire n16467_cascade_;
    wire n8_adj_1201;
    wire n15527;
    wire n14_adj_1189;
    wire n13_adj_1032;
    wire n13_adj_1032_cascade_;
    wire n8519;
    wire n22_adj_1115;
    wire n15651;
    wire n15526;
    wire buf_data1_20;
    wire n8058_cascade_;
    wire comm_buf_0_4;
    wire n15584;
    wire n83_cascade_;
    wire n15581;
    wire cmd_rdadctmp_29_adj_1083;
    wire buf_adcdata3_21;
    wire cmd_rdadctmp_23_adj_1089;
    wire buf_adcdata3_15;
    wire buf_data1_18;
    wire n75_adj_1164;
    wire comm_buf_1_0;
    wire data_cntvec_0;
    wire buf_data1_8;
    wire n4197_cascade_;
    wire n4221;
    wire n4234_cascade_;
    wire n4209;
    wire n4254_cascade_;
    wire n4264;
    wire n32_cascade_;
    wire n15557;
    wire data_idxvec_0;
    wire data_idxvec_15_N_673_0;
    wire bfn_17_12_0_;
    wire n14040;
    wire data_idxvec_2;
    wire n14041;
    wire n14042;
    wire n14_adj_1196;
    wire n14043;
    wire n14_adj_1213;
    wire n14044;
    wire data_idxvec_6;
    wire n14045;
    wire n14_adj_1168;
    wire data_idxvec_7;
    wire n14046;
    wire n14047;
    wire n14_adj_1211;
    wire bfn_17_13_0_;
    wire n14_adj_1210;
    wire data_idxvec_9;
    wire n14048;
    wire n14_adj_1209;
    wire data_idxvec_10;
    wire n14049;
    wire n14050;
    wire n14_adj_1207;
    wire data_idxvec_12;
    wire n14051;
    wire n14_adj_1202;
    wire data_idxvec_13;
    wire n14052;
    wire n14_adj_1206;
    wire data_idxvec_14;
    wire n14053;
    wire n14_adj_1205;
    wire n14054;
    wire n9187;
    wire buf_adcdata3_13;
    wire n14_adj_1198;
    wire cmd_rdadctmp_22;
    wire buf_adcdata1_14;
    wire req_data_cnt_11;
    wire n14_adj_1169;
    wire req_data_cnt_6;
    wire n4204;
    wire n4249_cascade_;
    wire n4259_cascade_;
    wire comm_buf_1_5;
    wire data_idxvec_4;
    wire data_cntvec_4;
    wire buf_data1_12;
    wire n4193_cascade_;
    wire req_data_cnt_5;
    wire acadc_skipCount_5;
    wire n4216;
    wire data_idxvec_5;
    wire data_cntvec_5;
    wire buf_data1_13;
    wire n4192_cascade_;
    wire n4229;
    wire cmd_rdadctmp_18_adj_1058;
    wire buf_adcdata2_10;
    wire data_idxvec_1;
    wire data_cntvec_1;
    wire cmd_rdadctmp_16_adj_1096;
    wire req_data_cnt_3;
    wire acadc_skipCount_3;
    wire eis_state_1;
    wire n9790;
    wire n10483;
    wire \comm_spi.n16887 ;
    wire \comm_spi.n10438 ;
    wire \comm_spi.iclk_N_802 ;
    wire \comm_spi.n16890 ;
    wire \comm_spi.n10455 ;
    wire \comm_spi.n16890_cascade_ ;
    wire \comm_spi.bit_cnt_3 ;
    wire \comm_spi.n12175 ;
    wire comm_buf_1_7;
    wire comm_buf_0_7;
    wire comm_index_0;
    wire n15381;
    wire n12846_cascade_;
    wire n4_adj_1179;
    wire n15204;
    wire n4_adj_1184_cascade_;
    wire n15290;
    wire n15241_cascade_;
    wire n15108;
    wire n15128;
    wire n8530;
    wire n15198;
    wire n15266;
    wire n15410_cascade_;
    wire n15130;
    wire n15408;
    wire n10394;
    wire n16190;
    wire n15635;
    wire n12_adj_1027;
    wire n12622;
    wire n14_adj_1152;
    wire n93;
    wire n27;
    wire n4;
    wire n15309_cascade_;
    wire comm_state_3_N_402_3;
    wire n15637;
    wire n13_adj_1040;
    wire n22_adj_1078;
    wire comm_rx_buf_7;
    wire comm_cmd_7;
    wire comm_rx_buf_0;
    wire comm_rx_buf_2;
    wire comm_buf_1_2;
    wire comm_rx_buf_4;
    wire n10363_cascade_;
    wire comm_rx_buf_5;
    wire n8062;
    wire n8085_cascade_;
    wire n24;
    wire comm_rx_buf_6;
    wire buf_data1_19;
    wire data_idxvec_11;
    wire n75;
    wire n12_cascade_;
    wire n6301;
    wire n8253;
    wire n14_adj_1197;
    wire req_data_cnt_2;
    wire comm_cmd_5;
    wire comm_cmd_4;
    wire comm_cmd_6;
    wire n8043;
    wire n7511;
    wire comm_buf_1_1;
    wire eis_start;
    wire data_idxvec_8;
    wire n78_adj_1022;
    wire buf_dds_3;
    wire n8;
    wire n15188;
    wire n12702;
    wire n15188_cascade_;
    wire n8085;
    wire n6_adj_1171_cascade_;
    wire n15190;
    wire buf_adcdata3_12;
    wire cmd_rdadctmp_21_adj_1091;
    wire n4_adj_1041;
    wire comm_buf_0_6;
    wire n8250;
    wire acadc_skipCount_14;
    wire data_idxvec_15;
    wire acadc_skipCount_15;
    wire n15468;
    wire n4217;
    wire n4230;
    wire n4250;
    wire cmd_rdadctmp_22_adj_1090;
    wire buf_adcdata3_14;
    wire n1;
    wire n8525;
    wire buf_dds_11;
    wire n12;
    wire n13_adj_1025;
    wire acadc_skipCount_1;
    wire req_data_cnt_1;
    wire n4220_cascade_;
    wire n4253_cascade_;
    wire n4263;
    wire buf_dds_1;
    wire buf_adcdata3_9;
    wire n4208;
    wire buf_data1_9;
    wire n4196;
    wire n4233;
    wire data_idxvec_3;
    wire data_cntvec_3;
    wire buf_data1_11;
    wire n4194_cascade_;
    wire n4218;
    wire n4231_cascade_;
    wire n4206;
    wire n4251_cascade_;
    wire buf_data2_9;
    wire buf_adcdata4_9;
    wire n4063;
    wire buf_adcdata2_11;
    wire n8_adj_1219;
    wire n7_adj_1218;
    wire data_index_9_N_258_8;
    wire \comm_spi.n10456 ;
    wire \comm_spi.iclk ;
    wire \comm_spi.n16893 ;
    wire \comm_spi.n10441 ;
    wire \comm_spi.n16893_cascade_ ;
    wire \comm_spi.imosi_cascade_ ;
    wire \comm_spi.DOUT_7__N_785 ;
    wire \comm_spi.imosi_N_791 ;
    wire cmd_rdadctmp_9_adj_1067;
    wire buf_adcdata2_1;
    wire \comm_spi.imosi ;
    wire \comm_spi.DOUT_7__N_786 ;
    wire n15131;
    wire n15241;
    wire n15191;
    wire n10148;
    wire n7;
    wire comm_state_3_N_418_1;
    wire n15711_cascade_;
    wire n8_adj_1193;
    wire n26_adj_1192_cascade_;
    wire n18_adj_1191;
    wire n15245;
    wire ICE_SPI_CE0;
    wire n15245_cascade_;
    wire comm_data_vld;
    wire n8544;
    wire n9_adj_1028;
    wire n9011;
    wire n9011_cascade_;
    wire n9215;
    wire buf_data2_19;
    wire buf_adcdata4_19;
    wire comm_buf_3_7_N_501_3;
    wire buf_control_6;
    wire n60;
    wire cmd_rdadctmp_8_adj_1104;
    wire buf_adcdata3_0;
    wire buf_adcdata3_11;
    wire cmd_rdadctmp_30_adj_1082;
    wire buf_adcdata3_22;
    wire n7_adj_1190;
    wire buf_dds_2;
    wire n4207;
    wire n8094;
    wire n729;
    wire buf_adcdata2_19;
    wire comm_buf_0_3;
    wire n14_adj_1208;
    wire cmd_rdadctmp_10;
    wire buf_adcdata1_2;
    wire n15147;
    wire buf_adcdata3_10;
    wire comm_rx_buf_1;
    wire n8618;
    wire n10363;
    wire cmd_rdadctmp_25_adj_1051;
    wire buf_adcdata2_18;
    wire n14_adj_1215;
    wire cmd_rdadctmp_26_adj_1050;
    wire cmd_rdadctmp_27_adj_1049;
    wire n4_adj_1250;
    wire buf_adcdata2_12;
    wire comm_cmd_2;
    wire comm_cmd_1;
    wire n9;
    wire comm_rx_buf_3;
    wire n4261;
    wire comm_buf_1_3;
    wire n8702;
    wire n10583;
    wire cmd_rdadctmp_21;
    wire buf_adcdata1_13;
    wire cmd_rdadctmp_17_adj_1095;
    wire cmd_rdadctmp_18_adj_1094;
    wire buf_adcdata2_13;
    wire cmd_rdadctmp_20;
    wire buf_adcdata1_12;
    wire cmd_rdadctmp_17_adj_1059;
    wire buf_adcdata2_9;
    wire cmd_rdadctmp_19_adj_1057;
    wire cmd_rdadctmp_20_adj_1056;
    wire n8302;
    wire cmd_rdadctmp_21_adj_1055;
    wire buf_data2_23;
    wire buf_adcdata4_23;
    wire n4101;
    wire \comm_spi.n10442 ;
    wire ICE_SPI_MOSI;
    wire \comm_spi.imosi_N_792 ;
    wire cmd_rdadctmp_28_adj_1048;
    wire buf_adcdata2_20;
    wire cmd_rdadctmp_31_adj_1045;
    wire buf_adcdata2_23;
    wire buf_data2_16;
    wire comm_cmd_0;
    wire buf_adcdata4_16;
    wire comm_cmd_3;
    wire n4108;
    wire cmd_rdadctmp_10_adj_1066;
    wire buf_adcdata2_2;
    wire \comm_spi.data_tx_7__N_808 ;
    wire comm_tx_buf_4;
    wire comm_clear;
    wire \comm_spi.n16899 ;
    wire cmd_rdadctmp_29_adj_1047;
    wire buf_adcdata2_21;
    wire ICE_GPMI_0;
    wire n8576;
    wire n8117;
    wire n6_adj_1175;
    wire comm_state_0;
    wire comm_state_1;
    wire comm_state_2;
    wire n8129;
    wire cmd_rdadctmp_19_adj_1093;
    wire adc_state_0_adj_1080;
    wire n8332;
    wire cmd_rdadctmp_20_adj_1092;
    wire n15640;
    wire n10_adj_1172;
    wire dds_state_1;
    wire dds_state_0;
    wire \CLOCK_DDS.n9 ;
    wire cmd_rdadctmp_24;
    wire buf_adcdata1_16;
    wire cmd_rdadctmp_30_adj_1046;
    wire buf_adcdata2_22;
    wire n15150;
    wire cmd_rdadctmp_22_adj_1054;
    wire adc_state_0_adj_1044;
    wire buf_adcdata2_14;
    wire n15153;
    wire cmd_rdadctmp_18;
    wire adc_state_0;
    wire buf_adcdata1_10;
    wire n8_adj_1225;
    wire comm_state_3;
    wire n6791;
    wire n7_adj_1224;
    wire data_index_9_N_258_5;
    wire ICE_SPI_SCLK;
    wire \comm_spi.n10437 ;
    wire _gnd_net_;
    wire clk_32MHz;
    wire \comm_spi.iclk_N_801 ;

    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_main.zim_pll_inst .TEST_MODE=1'b0;
    defparam \pll_main.zim_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll_main.zim_pll_inst .FILTER_RANGE=3'b011;
    defparam \pll_main.zim_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_main.zim_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_main.zim_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll_main.zim_pll_inst .DIVR=4'b0000;
    defparam \pll_main.zim_pll_inst .DIVQ=3'b101;
    defparam \pll_main.zim_pll_inst .DIVF=7'b0011111;
    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll_main.zim_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(),
            .REFERENCECLK(N__16769),
            .RESETB(N__28782),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(clk_16MHz),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(clk_32MHz),
            .SCLK(GNDG0));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical (
            .RDATA({dangling_wire_0,buf_data1_19,dangling_wire_1,buf_data4_19,dangling_wire_2,buf_data3_19,dangling_wire_3,buf_data2_19,dangling_wire_4,buf_data1_18,dangling_wire_5,buf_data4_18,dangling_wire_6,buf_data3_18,dangling_wire_7,buf_data2_18}),
            .RADDR({dangling_wire_8,dangling_wire_9,N__42539,N__30500,N__30356,N__51470,N__28157,N__32453,N__29660,N__28442,N__29840}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__35843,N__35951,N__36059,N__36167,N__36278,N__35039,N__35144,N__35249,N__35354}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,N__20237,dangling_wire_29,N__43031,dangling_wire_30,N__26225,dangling_wire_31,N__43580,dangling_wire_32,N__20042,dangling_wire_33,N__19295,dangling_wire_34,N__26465,dangling_wire_35,N__43937}),
            .RCLKE(),
            .RCLK(N__51259),
            .RE(N__28823),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN_net),
            .WE(N__28346));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical (
            .RDATA({dangling_wire_36,buf_data1_17,dangling_wire_37,buf_data4_17,dangling_wire_38,buf_data3_17,dangling_wire_39,buf_data2_17,dangling_wire_40,buf_data1_16,dangling_wire_41,buf_data4_16,dangling_wire_42,buf_data3_16,dangling_wire_43,buf_data2_16}),
            .RADDR({dangling_wire_44,dangling_wire_45,N__42533,N__30494,N__30350,N__51464,N__28151,N__32447,N__29654,N__28436,N__29834}),
            .WADDR({dangling_wire_46,dangling_wire_47,N__35837,N__35945,N__36053,N__36161,N__36272,N__35033,N__35138,N__35243,N__35348}),
            .MASK({dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63}),
            .WDATA({dangling_wire_64,N__20069,dangling_wire_65,N__25798,dangling_wire_66,N__27959,dangling_wire_67,N__20354,dangling_wire_68,N__48227,dangling_wire_69,N__47371,dangling_wire_70,N__26363,dangling_wire_71,N__21308}),
            .RCLKE(),
            .RCLK(N__51287),
            .RE(N__28837),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN_net),
            .WE(N__28272));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical (
            .RDATA({dangling_wire_72,buf_data1_7,dangling_wire_73,buf_data4_7,dangling_wire_74,buf_data3_7,dangling_wire_75,buf_data2_7,dangling_wire_76,buf_data1_6,dangling_wire_77,buf_data4_6,dangling_wire_78,buf_data3_6,dangling_wire_79,buf_data2_6}),
            .RADDR({dangling_wire_80,dangling_wire_81,N__42523,N__30481,N__30340,N__51460,N__28141,N__32440,N__29641,N__28426,N__29821}),
            .WADDR({dangling_wire_82,dangling_wire_83,N__35821,N__35929,N__36040,N__36148,N__36262,N__35020,N__35122,N__35227,N__35332}),
            .MASK({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99}),
            .WDATA({dangling_wire_100,N__17774,dangling_wire_101,N__17474,dangling_wire_102,N__18719,dangling_wire_103,N__17618,dangling_wire_104,N__21707,dangling_wire_105,N__17680,dangling_wire_106,N__19529,dangling_wire_107,N__17639}),
            .RCLKE(),
            .RCLK(N__51174),
            .RE(N__28802),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN_net),
            .WE(N__28345));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical (
            .RDATA({dangling_wire_108,buf_data1_15,dangling_wire_109,buf_data4_15,dangling_wire_110,buf_data3_15,dangling_wire_111,buf_data2_15,dangling_wire_112,buf_data1_14,dangling_wire_113,buf_data4_14,dangling_wire_114,buf_data3_14,dangling_wire_115,buf_data2_14}),
            .RADDR({dangling_wire_116,dangling_wire_117,N__42527,N__30488,N__30344,N__51457,N__28145,N__32441,N__29648,N__28430,N__29828}),
            .WADDR({dangling_wire_118,dangling_wire_119,N__35831,N__35939,N__36047,N__36155,N__36266,N__35027,N__35132,N__35237,N__35342}),
            .MASK({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .WDATA({dangling_wire_136,N__22688,dangling_wire_137,N__26002,dangling_wire_138,N__36770,dangling_wire_139,N__34445,dangling_wire_140,N__37445,dangling_wire_141,N__24107,dangling_wire_142,N__41558,dangling_wire_143,N__53144}),
            .RCLKE(),
            .RCLK(N__51305),
            .RE(N__28838),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN_net),
            .WE(N__28322));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical (
            .RDATA({dangling_wire_144,buf_data1_5,dangling_wire_145,buf_data4_5,dangling_wire_146,buf_data3_5,dangling_wire_147,buf_data2_5,dangling_wire_148,buf_data1_4,dangling_wire_149,buf_data4_4,dangling_wire_150,buf_data3_4,dangling_wire_151,buf_data2_4}),
            .RADDR({dangling_wire_152,dangling_wire_153,N__42511,N__30469,N__30328,N__51448,N__28129,N__32428,N__29629,N__28414,N__29809}),
            .WADDR({dangling_wire_154,dangling_wire_155,N__35809,N__35917,N__36028,N__36136,N__36250,N__35008,N__35110,N__35215,N__35320}),
            .MASK({dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171}),
            .WDATA({dangling_wire_172,N__17792,dangling_wire_173,N__17752,dangling_wire_174,N__19564,dangling_wire_175,N__17657,dangling_wire_176,N__18635,dangling_wire_177,N__18125,dangling_wire_178,N__18760,dangling_wire_179,N__17885}),
            .RCLKE(),
            .RCLK(N__51209),
            .RE(N__28821),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN_net),
            .WE(N__28344));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical (
            .RDATA({dangling_wire_180,buf_data1_1,dangling_wire_181,buf_data4_1,dangling_wire_182,buf_data3_1,dangling_wire_183,buf_data2_1,dangling_wire_184,buf_data1_0,dangling_wire_185,buf_data4_0,dangling_wire_186,buf_data3_0,dangling_wire_187,buf_data2_0}),
            .RADDR({dangling_wire_188,dangling_wire_189,N__42545,N__30506,N__30362,N__51476,N__28163,N__32459,N__29666,N__28448,N__29846}),
            .WADDR({dangling_wire_190,dangling_wire_191,N__35849,N__35957,N__36065,N__36173,N__36284,N__35045,N__35150,N__35255,N__35360}),
            .MASK({dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207}),
            .WDATA({dangling_wire_208,N__21260,dangling_wire_209,N__17993,dangling_wire_210,N__27593,dangling_wire_211,N__42908,dangling_wire_212,N__22451,dangling_wire_213,N__18029,dangling_wire_214,N__43810,dangling_wire_215,N__17225}),
            .RCLKE(),
            .RCLK(N__51226),
            .RE(N__28822),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN_net),
            .WE(N__28340));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical (
            .RDATA({dangling_wire_216,buf_data1_13,dangling_wire_217,buf_data4_13,dangling_wire_218,buf_data3_13,dangling_wire_219,buf_data2_13,dangling_wire_220,buf_data1_12,dangling_wire_221,buf_data4_12,dangling_wire_222,buf_data3_12,dangling_wire_223,buf_data2_12}),
            .RADDR({dangling_wire_224,dangling_wire_225,N__42520,N__30482,N__30337,N__51445,N__28138,N__32431,N__29642,N__28423,N__29822}),
            .WADDR({dangling_wire_226,dangling_wire_227,N__35825,N__35933,N__36041,N__36149,N__36259,N__35021,N__35126,N__35231,N__35336}),
            .MASK({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243}),
            .WDATA({dangling_wire_244,N__44563,dangling_wire_245,N__28615,dangling_wire_246,N__37520,dangling_wire_247,N__44486,dangling_wire_248,N__46256,dangling_wire_249,N__20495,dangling_wire_250,N__40783,dangling_wire_251,N__45680}),
            .RCLKE(),
            .RCLK(N__51313),
            .RE(N__28848),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN_net),
            .WE(N__28353));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical (
            .RDATA({dangling_wire_252,buf_data1_23,dangling_wire_253,buf_data4_23,dangling_wire_254,buf_data3_23,dangling_wire_255,buf_data2_23,dangling_wire_256,buf_data1_22,dangling_wire_257,buf_data4_22,dangling_wire_258,buf_data3_22,dangling_wire_259,buf_data2_22}),
            .RADDR({dangling_wire_260,dangling_wire_261,N__42563,N__30524,N__30380,N__51494,N__28181,N__32477,N__29684,N__28466,N__29864}),
            .WADDR({dangling_wire_262,dangling_wire_263,N__35867,N__35975,N__36083,N__36191,N__36302,N__35063,N__35168,N__35273,N__35378}),
            .MASK({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279}),
            .WDATA({dangling_wire_280,N__22736,dangling_wire_281,N__45878,dangling_wire_282,N__25685,dangling_wire_283,N__48122,dangling_wire_284,N__21365,dangling_wire_285,N__29078,dangling_wire_286,N__43718,dangling_wire_287,N__48179}),
            .RCLKE(),
            .RCLK(N__51134),
            .RE(N__28774),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN_net),
            .WE(N__28364));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical (
            .RDATA({dangling_wire_288,buf_data1_3,dangling_wire_289,buf_data4_3,dangling_wire_290,buf_data3_3,dangling_wire_291,buf_data2_3,dangling_wire_292,buf_data1_2,dangling_wire_293,buf_data4_2,dangling_wire_294,buf_data3_2,dangling_wire_295,buf_data2_2}),
            .RADDR({dangling_wire_296,dangling_wire_297,N__42551,N__30512,N__30368,N__51482,N__28169,N__32465,N__29672,N__28454,N__29852}),
            .WADDR({dangling_wire_298,dangling_wire_299,N__35855,N__35963,N__36071,N__36179,N__36290,N__35051,N__35156,N__35261,N__35366}),
            .MASK({dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .WDATA({dangling_wire_316,N__18785,dangling_wire_317,N__20819,dangling_wire_318,N__32624,dangling_wire_319,N__17582,dangling_wire_320,N__44426,dangling_wire_321,N__17921,dangling_wire_322,N__18482,dangling_wire_323,N__46666}),
            .RCLKE(),
            .RCLK(N__51192),
            .RE(N__28807),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN_net),
            .WE(N__28359));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical (
            .RDATA({dangling_wire_324,buf_data1_11,dangling_wire_325,buf_data4_11,dangling_wire_326,buf_data3_11,dangling_wire_327,buf_data2_11,dangling_wire_328,buf_data1_10,dangling_wire_329,buf_data4_10,dangling_wire_330,buf_data3_10,dangling_wire_331,buf_data2_10}),
            .RADDR({dangling_wire_332,dangling_wire_333,N__42508,N__30472,N__30325,N__51433,N__28126,N__32419,N__29632,N__28411,N__29812}),
            .WADDR({dangling_wire_334,dangling_wire_335,N__35818,N__35926,N__36031,N__36139,N__36247,N__35011,N__35119,N__35224,N__35329}),
            .MASK({dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .WDATA({dangling_wire_352,N__24539,dangling_wire_353,N__26552,dangling_wire_354,N__43778,dangling_wire_355,N__42620,dangling_wire_356,N__52505,dangling_wire_357,N__19708,dangling_wire_358,N__44207,dangling_wire_359,N__38261}),
            .RCLKE(),
            .RCLK(N__51317),
            .RE(N__28849),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN_net),
            .WE(N__28354));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical (
            .RDATA({dangling_wire_360,buf_data1_21,dangling_wire_361,buf_data4_21,dangling_wire_362,buf_data3_21,dangling_wire_363,buf_data2_21,dangling_wire_364,buf_data1_20,dangling_wire_365,buf_data4_20,dangling_wire_366,buf_data3_20,dangling_wire_367,buf_data2_20}),
            .RADDR({dangling_wire_368,dangling_wire_369,N__42557,N__30518,N__30374,N__51488,N__28175,N__32471,N__29678,N__28460,N__29858}),
            .WADDR({dangling_wire_370,dangling_wire_371,N__35861,N__35969,N__36077,N__36185,N__36296,N__35057,N__35162,N__35267,N__35372}),
            .MASK({dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387}),
            .WDATA({dangling_wire_388,N__21167,dangling_wire_389,N__23173,dangling_wire_390,N__36845,dangling_wire_391,N__46331,dangling_wire_392,N__20189,dangling_wire_393,N__24653,dangling_wire_394,N__24073,dangling_wire_395,N__45707}),
            .RCLKE(),
            .RCLK(N__51158),
            .RE(N__28806),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN_net),
            .WE(N__28358));
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.WRITE_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.READ_MODE=1;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical (
            .RDATA({dangling_wire_396,buf_data1_9,dangling_wire_397,buf_data4_9,dangling_wire_398,buf_data3_9,dangling_wire_399,buf_data2_9,dangling_wire_400,buf_data1_8,dangling_wire_401,buf_data4_8,dangling_wire_402,buf_data3_8,dangling_wire_403,buf_data2_8}),
            .RADDR({dangling_wire_404,dangling_wire_405,N__42496,N__30460,N__30313,N__51421,N__28114,N__32407,N__29620,N__28399,N__29800}),
            .WADDR({dangling_wire_406,dangling_wire_407,N__35806,N__35914,N__36019,N__36127,N__36235,N__34999,N__35107,N__35212,N__35317}),
            .MASK({dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423}),
            .WDATA({dangling_wire_424,N__24602,dangling_wire_425,N__42670,dangling_wire_426,N__42095,dangling_wire_427,N__46202,dangling_wire_428,N__32147,dangling_wire_429,N__24350,dangling_wire_430,N__24511,dangling_wire_431,N__20420}),
            .RCLKE(),
            .RCLK(N__51319),
            .RE(N__28853),
            .WCLKE(),
            .WCLK(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN_net),
            .WE(N__28363));
    IO_PAD ipInertedIOPad_M_CS1_iopad (
            .OE(N__54255),
            .DIN(N__54254),
            .DOUT(N__54253),
            .PACKAGEPIN(M_CS1));
    defparam ipInertedIOPad_M_CS1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CS1_preio (
            .PADOEN(N__54255),
            .PADOUT(N__54254),
            .PADIN(N__54253),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18920),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_SYSCLK_iopad (
            .OE(N__54246),
            .DIN(N__54245),
            .DOUT(N__54244),
            .PACKAGEPIN(ICE_SYSCLK));
    defparam ipInertedIOPad_ICE_SYSCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SYSCLK_preio (
            .PADOEN(N__54246),
            .PADOUT(N__54245),
            .PADIN(N__54244),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SYSCLK),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MOSI1_iopad (
            .OE(N__54237),
            .DIN(N__54236),
            .DOUT(N__54235),
            .PACKAGEPIN(M_MOSI1));
    defparam ipInertedIOPad_M_MOSI1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_MOSI1_preio (
            .PADOEN(N__54237),
            .PADOUT(N__54236),
            .PADIN(N__54235),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_DRDY1_iopad (
            .OE(N__54228),
            .DIN(N__54227),
            .DOUT(N__54226),
            .PACKAGEPIN(M_DRDY1));
    defparam ipInertedIOPad_M_DRDY1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_DRDY1_preio (
            .PADOEN(N__54228),
            .PADOUT(N__54227),
            .PADIN(N__54226),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_DRDY1),
            .DIN1());
    IO_PAD ipInertedIOPad_M_CLK2_iopad (
            .OE(N__54219),
            .DIN(N__54218),
            .DOUT(N__54217),
            .PACKAGEPIN(M_CLK2));
    defparam ipInertedIOPad_M_CLK2_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CLK2_preio (
            .PADOEN(N__54219),
            .PADOUT(N__54218),
            .PADIN(N__54217),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16753),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_SCLK1_iopad (
            .OE(N__54210),
            .DIN(N__54209),
            .DOUT(N__54208),
            .PACKAGEPIN(M_SCLK1));
    defparam ipInertedIOPad_M_SCLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_SCLK1_preio (
            .PADOEN(N__54210),
            .PADOUT(N__54209),
            .PADIN(N__54208),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18890),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_FLT0_iopad (
            .OE(N__54201),
            .DIN(N__54200),
            .DOUT(N__54199),
            .PACKAGEPIN(M_FLT0));
    defparam ipInertedIOPad_M_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_FLT0_preio (
            .PADOEN(N__54201),
            .PADOUT(N__54200),
            .PADIN(N__54199),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__28568),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_CS3_iopad (
            .OE(N__54192),
            .DIN(N__54191),
            .DOUT(N__54190),
            .PACKAGEPIN(M_CS3));
    defparam ipInertedIOPad_M_CS3_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CS3_preio (
            .PADOEN(N__54192),
            .PADOUT(N__54191),
            .PADIN(N__54190),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20708),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_CHKCABLE_iopad (
            .OE(N__54183),
            .DIN(N__54182),
            .DOUT(N__54181),
            .PACKAGEPIN(ICE_CHKCABLE));
    defparam ipInertedIOPad_ICE_CHKCABLE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_CHKCABLE_preio (
            .PADOEN(N__54183),
            .PADOUT(N__54182),
            .PADIN(N__54181),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_CHKCABLE),
            .DIN1());
    IO_PAD ipInertedIOPad_M_OSR1_iopad (
            .OE(N__54174),
            .DIN(N__54173),
            .DOUT(N__54172),
            .PACKAGEPIN(M_OSR1));
    defparam ipInertedIOPad_M_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_OSR1_preio (
            .PADOEN(N__54174),
            .PADOUT(N__54173),
            .PADIN(N__54172),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29441),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_1_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_1_iopad (
            .OE(N__54165),
            .DIN(N__54164),
            .DOUT(N__54163),
            .PACKAGEPIN(ICE_GPMO_1));
    defparam ipInertedIOPad_ICE_GPMO_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_1_preio (
            .PADOEN(N__54165),
            .PADOUT(N__54164),
            .PADIN(N__54163),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_EIS_SYNCCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_EIS_SYNCCLK_iopad (
            .OE(N__54156),
            .DIN(N__54155),
            .DOUT(N__54154),
            .PACKAGEPIN(EIS_SYNCCLK));
    defparam ipInertedIOPad_EIS_SYNCCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_EIS_SYNCCLK_preio (
            .PADOEN(N__54156),
            .PADOUT(N__54155),
            .PADIN(N__54154),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_CLK4),
            .DIN1());
    IO_PAD ipInertedIOPad_M_SCLK3_iopad (
            .OE(N__54147),
            .DIN(N__54146),
            .DOUT(N__54145),
            .PACKAGEPIN(M_SCLK3));
    defparam ipInertedIOPad_M_SCLK3_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_SCLK3_preio (
            .PADOEN(N__54147),
            .PADOUT(N__54146),
            .PADIN(N__54145),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20678),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_OSR0_iopad (
            .OE(N__54138),
            .DIN(N__54137),
            .DOUT(N__54136),
            .PACKAGEPIN(M_OSR0));
    defparam ipInertedIOPad_M_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_OSR0_preio (
            .PADOEN(N__54138),
            .PADOUT(N__54137),
            .PADIN(N__54136),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__28085),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MISO4_iopad (
            .OE(N__54129),
            .DIN(N__54128),
            .DOUT(N__54127),
            .PACKAGEPIN(M_MISO4));
    defparam ipInertedIOPad_M_MISO4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_MISO4_preio (
            .PADOEN(N__54129),
            .PADOUT(N__54128),
            .PADIN(N__54127),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_MISO4),
            .DIN1());
    IO_PAD ipInertedIOPad_M_DRDY4_iopad (
            .OE(N__54120),
            .DIN(N__54119),
            .DOUT(N__54118),
            .PACKAGEPIN(M_DRDY4));
    defparam ipInertedIOPad_M_DRDY4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_DRDY4_preio (
            .PADOEN(N__54120),
            .PADOUT(N__54119),
            .PADIN(N__54118),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_DRDY4),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_MOSI_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_MOSI_iopad (
            .OE(N__54111),
            .DIN(N__54110),
            .DOUT(N__54109),
            .PACKAGEPIN(ICE_SPI_MOSI));
    defparam ipInertedIOPad_ICE_SPI_MOSI_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_MOSI_preio (
            .PADOEN(N__54111),
            .PADOUT(N__54110),
            .PADIN(N__54109),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_MOSI),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_0_iopad (
            .OE(N__54102),
            .DIN(N__54101),
            .DOUT(N__54100),
            .PACKAGEPIN(ICE_GPMO_0));
    defparam ipInertedIOPad_ICE_GPMO_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_0_preio (
            .PADOEN(N__54102),
            .PADOUT(N__54101),
            .PADIN(N__54100),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_0),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI1_iopad (
            .OE(N__54093),
            .DIN(N__54092),
            .DOUT(N__54091),
            .PACKAGEPIN(DDS_MOSI1));
    defparam ipInertedIOPad_DDS_MOSI1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI1_preio (
            .PADOEN(N__54093),
            .PADOUT(N__54092),
            .PADIN(N__54091),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21224),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_SCLK4_iopad (
            .OE(N__54084),
            .DIN(N__54083),
            .DOUT(N__54082),
            .PACKAGEPIN(M_SCLK4));
    defparam ipInertedIOPad_M_SCLK4_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_SCLK4_preio (
            .PADOEN(N__54084),
            .PADOUT(N__54083),
            .PADIN(N__54082),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21650),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MISO3_iopad (
            .OE(N__54075),
            .DIN(N__54074),
            .DOUT(N__54073),
            .PACKAGEPIN(M_MISO3));
    defparam ipInertedIOPad_M_MISO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_MISO3_preio (
            .PADOEN(N__54075),
            .PADOUT(N__54074),
            .PADIN(N__54073),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_MISO3),
            .DIN1());
    IO_PAD ipInertedIOPad_M_CS4_iopad (
            .OE(N__54066),
            .DIN(N__54065),
            .DOUT(N__54064),
            .PACKAGEPIN(M_CS4));
    defparam ipInertedIOPad_M_CS4_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CS4_preio (
            .PADOEN(N__54066),
            .PADOUT(N__54065),
            .PADIN(N__54064),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26594),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_SCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_SCLK_iopad (
            .OE(N__54057),
            .DIN(N__54056),
            .DOUT(N__54055),
            .PACKAGEPIN(ICE_SPI_SCLK));
    defparam ipInertedIOPad_ICE_SPI_SCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_SCLK_preio (
            .PADOEN(N__54057),
            .PADOUT(N__54056),
            .PADIN(N__54055),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_SCLK),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MOSI4_iopad (
            .OE(N__54048),
            .DIN(N__54047),
            .DOUT(N__54046),
            .PACKAGEPIN(M_MOSI4));
    defparam ipInertedIOPad_M_MOSI4_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_MOSI4_preio (
            .PADOEN(N__54048),
            .PADOUT(N__54047),
            .PADIN(N__54046),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MISO2_iopad (
            .OE(N__54039),
            .DIN(N__54038),
            .DOUT(N__54037),
            .PACKAGEPIN(M_MISO2));
    defparam ipInertedIOPad_M_MISO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_MISO2_preio (
            .PADOEN(N__54039),
            .PADOUT(N__54038),
            .PADIN(N__54037),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_MISO2),
            .DIN1());
    IO_PAD ipInertedIOPad_M_DRDY2_iopad (
            .OE(N__54030),
            .DIN(N__54029),
            .DOUT(N__54028),
            .PACKAGEPIN(M_DRDY2));
    defparam ipInertedIOPad_M_DRDY2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_DRDY2_preio (
            .PADOEN(N__54030),
            .PADOUT(N__54029),
            .PADIN(N__54028),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_DRDY2),
            .DIN1());
    IO_PAD ipInertedIOPad_M_CLK1_iopad (
            .OE(N__54021),
            .DIN(N__54020),
            .DOUT(N__54019),
            .PACKAGEPIN(M_CLK1));
    defparam ipInertedIOPad_M_CLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CLK1_preio (
            .PADOEN(N__54021),
            .PADOUT(N__54020),
            .PADIN(N__54019),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16745),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_SPI_MISO_iopad (
            .OE(N__54012),
            .DIN(N__54011),
            .DOUT(N__54010),
            .PACKAGEPIN(ICE_SPI_MISO));
    defparam ipInertedIOPad_ICE_SPI_MISO_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_SPI_MISO_preio (
            .PADOEN(N__54012),
            .PADOUT(N__54011),
            .PADIN(N__54010),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30290),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_2_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_2_iopad (
            .OE(N__54003),
            .DIN(N__54002),
            .DOUT(N__54001),
            .PACKAGEPIN(ICE_GPMO_2));
    defparam ipInertedIOPad_ICE_GPMO_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_2_preio (
            .PADOEN(N__54003),
            .PADOUT(N__54002),
            .PADIN(N__54001),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_2),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_GPMI_0_iopad (
            .OE(N__53994),
            .DIN(N__53993),
            .DOUT(N__53992),
            .PACKAGEPIN(ICE_GPMI_0));
    defparam ipInertedIOPad_ICE_GPMI_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_GPMI_0_preio (
            .PADOEN(N__53994),
            .PADOUT(N__53993),
            .PADIN(N__53992),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__46313),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TEST_LED_iopad (
            .OE(N__53985),
            .DIN(N__53984),
            .DOUT(N__53983),
            .PACKAGEPIN(TEST_LED));
    defparam ipInertedIOPad_TEST_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_TEST_LED_preio (
            .PADOEN(N__53985),
            .PADOUT(N__53984),
            .PADIN(N__53983),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16796),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_POW_iopad (
            .OE(N__53976),
            .DIN(N__53975),
            .DOUT(N__53974),
            .PACKAGEPIN(M_POW));
    defparam ipInertedIOPad_M_POW_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_POW_preio (
            .PADOEN(N__53976),
            .PADOUT(N__53975),
            .PADIN(N__53974),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26267),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MOSI3_iopad (
            .OE(N__53967),
            .DIN(N__53966),
            .DOUT(N__53965),
            .PACKAGEPIN(M_MOSI3));
    defparam ipInertedIOPad_M_MOSI3_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_MOSI3_preio (
            .PADOEN(N__53967),
            .PADOUT(N__53966),
            .PADIN(N__53965),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MISO1_iopad (
            .OE(N__53958),
            .DIN(N__53957),
            .DOUT(N__53956),
            .PACKAGEPIN(M_MISO1));
    defparam ipInertedIOPad_M_MISO1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_MISO1_preio (
            .PADOEN(N__53958),
            .PADOUT(N__53957),
            .PADIN(N__53956),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_MISO1),
            .DIN1());
    IO_PAD ipInertedIOPad_M_DRDY3_iopad (
            .OE(N__53949),
            .DIN(N__53948),
            .DOUT(N__53947),
            .PACKAGEPIN(M_DRDY3));
    defparam ipInertedIOPad_M_DRDY3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_M_DRDY3_preio (
            .PADOEN(N__53949),
            .PADOUT(N__53948),
            .PADIN(N__53947),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(M_DRDY3),
            .DIN1());
    IO_PAD ipInertedIOPad_M_DCSEL_iopad (
            .OE(N__53940),
            .DIN(N__53939),
            .DOUT(N__53938),
            .PACKAGEPIN(M_DCSEL));
    defparam ipInertedIOPad_M_DCSEL_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_DCSEL_preio (
            .PADOEN(N__53940),
            .PADOUT(N__53939),
            .PADIN(N__53938),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27932),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_START_iopad (
            .OE(N__53931),
            .DIN(N__53930),
            .DOUT(N__53929),
            .PACKAGEPIN(M_START));
    defparam ipInertedIOPad_M_START_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_START_preio (
            .PADOEN(N__53931),
            .PADOUT(N__53930),
            .PADIN(N__53929),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19766),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_MOSI2_iopad (
            .OE(N__53922),
            .DIN(N__53921),
            .DOUT(N__53920),
            .PACKAGEPIN(M_MOSI2));
    defparam ipInertedIOPad_M_MOSI2_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_MOSI2_preio (
            .PADOEN(N__53922),
            .PADOUT(N__53921),
            .PADIN(N__53920),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_CLK3_iopad (
            .OE(N__53913),
            .DIN(N__53912),
            .DOUT(N__53911),
            .PACKAGEPIN(M_CLK3));
    defparam ipInertedIOPad_M_CLK3_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CLK3_preio (
            .PADOEN(N__53913),
            .PADOUT(N__53912),
            .PADIN(N__53911),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16749),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS1_iopad (
            .OE(N__53904),
            .DIN(N__53903),
            .DOUT(N__53902),
            .PACKAGEPIN(DDS_CS1));
    defparam ipInertedIOPad_DDS_CS1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS1_preio (
            .PADOEN(N__53904),
            .PADOUT(N__53903),
            .PADIN(N__53902),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26900),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_FLT1_iopad (
            .OE(N__53895),
            .DIN(N__53894),
            .DOUT(N__53893),
            .PACKAGEPIN(M_FLT1));
    defparam ipInertedIOPad_M_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_FLT1_preio (
            .PADOEN(N__53895),
            .PADOUT(N__53894),
            .PADIN(N__53893),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29585),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DISP_COMM_iopad (
            .OE(N__53886),
            .DIN(N__53885),
            .DOUT(N__53884),
            .PACKAGEPIN(DISP_COMM));
    defparam ipInertedIOPad_DISP_COMM_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DISP_COMM_preio (
            .PADOEN(N__53886),
            .PADOUT(N__53885),
            .PADIN(N__53884),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16673),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK1_iopad (
            .OE(N__53877),
            .DIN(N__53876),
            .DOUT(N__53875),
            .PACKAGEPIN(DDS_MCLK1));
    defparam ipInertedIOPad_DDS_MCLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK1_preio (
            .PADOEN(N__53877),
            .PADOUT(N__53876),
            .PADIN(N__53875),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16889),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_CE0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_CE0_iopad (
            .OE(N__53868),
            .DIN(N__53867),
            .DOUT(N__53866),
            .PACKAGEPIN(ICE_SPI_CE0));
    defparam ipInertedIOPad_ICE_SPI_CE0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_CE0_preio (
            .PADOEN(N__53868),
            .PADOUT(N__53867),
            .PADIN(N__53866),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_CE0),
            .DIN1());
    IO_PAD ipInertedIOPad_M_SCLK2_iopad (
            .OE(N__53859),
            .DIN(N__53858),
            .DOUT(N__53857),
            .PACKAGEPIN(M_SCLK2));
    defparam ipInertedIOPad_M_SCLK2_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_SCLK2_preio (
            .PADOEN(N__53859),
            .PADOUT(N__53858),
            .PADIN(N__53857),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19361),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_CS2_iopad (
            .OE(N__53850),
            .DIN(N__53849),
            .DOUT(N__53848),
            .PACKAGEPIN(M_CS2));
    defparam ipInertedIOPad_M_CS2_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CS2_preio (
            .PADOEN(N__53850),
            .PADOUT(N__53849),
            .PADIN(N__53848),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17387),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_M_CLK4_iopad (
            .OE(N__53841),
            .DIN(N__53840),
            .DOUT(N__53839),
            .PACKAGEPIN(M_CLK4));
    defparam ipInertedIOPad_M_CLK4_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_M_CLK4_preio (
            .PADOEN(N__53841),
            .PADOUT(N__53840),
            .PADIN(N__53839),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16754),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK1_iopad (
            .OE(N__53832),
            .DIN(N__53831),
            .DOUT(N__53830),
            .PACKAGEPIN(DDS_SCK1));
    defparam ipInertedIOPad_DDS_SCK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK1_preio (
            .PADOEN(N__53832),
            .PADOUT(N__53831),
            .PADIN(N__53830),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21059),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__13727 (
            .O(N__53813),
            .I(N__53806));
    InMux I__13726 (
            .O(N__53812),
            .I(N__53803));
    InMux I__13725 (
            .O(N__53811),
            .I(N__53800));
    InMux I__13724 (
            .O(N__53810),
            .I(N__53795));
    InMux I__13723 (
            .O(N__53809),
            .I(N__53792));
    LocalMux I__13722 (
            .O(N__53806),
            .I(N__53785));
    LocalMux I__13721 (
            .O(N__53803),
            .I(N__53785));
    LocalMux I__13720 (
            .O(N__53800),
            .I(N__53785));
    InMux I__13719 (
            .O(N__53799),
            .I(N__53782));
    InMux I__13718 (
            .O(N__53798),
            .I(N__53779));
    LocalMux I__13717 (
            .O(N__53795),
            .I(N__53776));
    LocalMux I__13716 (
            .O(N__53792),
            .I(N__53771));
    Span4Mux_v I__13715 (
            .O(N__53785),
            .I(N__53766));
    LocalMux I__13714 (
            .O(N__53782),
            .I(N__53766));
    LocalMux I__13713 (
            .O(N__53779),
            .I(N__53761));
    Span4Mux_h I__13712 (
            .O(N__53776),
            .I(N__53761));
    InMux I__13711 (
            .O(N__53775),
            .I(N__53758));
    InMux I__13710 (
            .O(N__53774),
            .I(N__53755));
    Span4Mux_h I__13709 (
            .O(N__53771),
            .I(N__53740));
    Span4Mux_v I__13708 (
            .O(N__53766),
            .I(N__53740));
    Span4Mux_v I__13707 (
            .O(N__53761),
            .I(N__53740));
    LocalMux I__13706 (
            .O(N__53758),
            .I(N__53740));
    LocalMux I__13705 (
            .O(N__53755),
            .I(N__53740));
    InMux I__13704 (
            .O(N__53754),
            .I(N__53735));
    InMux I__13703 (
            .O(N__53753),
            .I(N__53735));
    InMux I__13702 (
            .O(N__53752),
            .I(N__53730));
    InMux I__13701 (
            .O(N__53751),
            .I(N__53727));
    Span4Mux_v I__13700 (
            .O(N__53740),
            .I(N__53722));
    LocalMux I__13699 (
            .O(N__53735),
            .I(N__53722));
    InMux I__13698 (
            .O(N__53734),
            .I(N__53717));
    InMux I__13697 (
            .O(N__53733),
            .I(N__53717));
    LocalMux I__13696 (
            .O(N__53730),
            .I(N__53713));
    LocalMux I__13695 (
            .O(N__53727),
            .I(N__53710));
    Span4Mux_v I__13694 (
            .O(N__53722),
            .I(N__53705));
    LocalMux I__13693 (
            .O(N__53717),
            .I(N__53705));
    InMux I__13692 (
            .O(N__53716),
            .I(N__53699));
    Span4Mux_h I__13691 (
            .O(N__53713),
            .I(N__53692));
    Span4Mux_h I__13690 (
            .O(N__53710),
            .I(N__53689));
    Span4Mux_v I__13689 (
            .O(N__53705),
            .I(N__53686));
    InMux I__13688 (
            .O(N__53704),
            .I(N__53678));
    InMux I__13687 (
            .O(N__53703),
            .I(N__53678));
    InMux I__13686 (
            .O(N__53702),
            .I(N__53678));
    LocalMux I__13685 (
            .O(N__53699),
            .I(N__53675));
    InMux I__13684 (
            .O(N__53698),
            .I(N__53672));
    InMux I__13683 (
            .O(N__53697),
            .I(N__53669));
    InMux I__13682 (
            .O(N__53696),
            .I(N__53664));
    InMux I__13681 (
            .O(N__53695),
            .I(N__53664));
    Span4Mux_h I__13680 (
            .O(N__53692),
            .I(N__53661));
    Span4Mux_v I__13679 (
            .O(N__53689),
            .I(N__53656));
    Span4Mux_h I__13678 (
            .O(N__53686),
            .I(N__53656));
    InMux I__13677 (
            .O(N__53685),
            .I(N__53653));
    LocalMux I__13676 (
            .O(N__53678),
            .I(N__53650));
    Span4Mux_h I__13675 (
            .O(N__53675),
            .I(N__53647));
    LocalMux I__13674 (
            .O(N__53672),
            .I(N__53642));
    LocalMux I__13673 (
            .O(N__53669),
            .I(N__53642));
    LocalMux I__13672 (
            .O(N__53664),
            .I(N__53639));
    Span4Mux_h I__13671 (
            .O(N__53661),
            .I(N__53636));
    Sp12to4 I__13670 (
            .O(N__53656),
            .I(N__53633));
    LocalMux I__13669 (
            .O(N__53653),
            .I(N__53626));
    Span4Mux_h I__13668 (
            .O(N__53650),
            .I(N__53626));
    Span4Mux_h I__13667 (
            .O(N__53647),
            .I(N__53626));
    Span4Mux_h I__13666 (
            .O(N__53642),
            .I(N__53619));
    Span4Mux_v I__13665 (
            .O(N__53639),
            .I(N__53619));
    Span4Mux_v I__13664 (
            .O(N__53636),
            .I(N__53619));
    Span12Mux_h I__13663 (
            .O(N__53633),
            .I(N__53616));
    Odrv4 I__13662 (
            .O(N__53626),
            .I(n15150));
    Odrv4 I__13661 (
            .O(N__53619),
            .I(n15150));
    Odrv12 I__13660 (
            .O(N__53616),
            .I(n15150));
    CascadeMux I__13659 (
            .O(N__53609),
            .I(N__53606));
    InMux I__13658 (
            .O(N__53606),
            .I(N__53602));
    InMux I__13657 (
            .O(N__53605),
            .I(N__53599));
    LocalMux I__13656 (
            .O(N__53602),
            .I(N__53596));
    LocalMux I__13655 (
            .O(N__53599),
            .I(N__53593));
    Span4Mux_h I__13654 (
            .O(N__53596),
            .I(N__53589));
    Span4Mux_h I__13653 (
            .O(N__53593),
            .I(N__53586));
    InMux I__13652 (
            .O(N__53592),
            .I(N__53583));
    Odrv4 I__13651 (
            .O(N__53589),
            .I(cmd_rdadctmp_22_adj_1054));
    Odrv4 I__13650 (
            .O(N__53586),
            .I(cmd_rdadctmp_22_adj_1054));
    LocalMux I__13649 (
            .O(N__53583),
            .I(cmd_rdadctmp_22_adj_1054));
    CascadeMux I__13648 (
            .O(N__53576),
            .I(N__53566));
    InMux I__13647 (
            .O(N__53575),
            .I(N__53561));
    InMux I__13646 (
            .O(N__53574),
            .I(N__53561));
    InMux I__13645 (
            .O(N__53573),
            .I(N__53552));
    InMux I__13644 (
            .O(N__53572),
            .I(N__53552));
    InMux I__13643 (
            .O(N__53571),
            .I(N__53552));
    InMux I__13642 (
            .O(N__53570),
            .I(N__53552));
    InMux I__13641 (
            .O(N__53569),
            .I(N__53549));
    InMux I__13640 (
            .O(N__53566),
            .I(N__53546));
    LocalMux I__13639 (
            .O(N__53561),
            .I(N__53543));
    LocalMux I__13638 (
            .O(N__53552),
            .I(N__53540));
    LocalMux I__13637 (
            .O(N__53549),
            .I(N__53528));
    LocalMux I__13636 (
            .O(N__53546),
            .I(N__53510));
    Span4Mux_v I__13635 (
            .O(N__53543),
            .I(N__53510));
    Span4Mux_h I__13634 (
            .O(N__53540),
            .I(N__53507));
    InMux I__13633 (
            .O(N__53539),
            .I(N__53494));
    InMux I__13632 (
            .O(N__53538),
            .I(N__53494));
    InMux I__13631 (
            .O(N__53537),
            .I(N__53494));
    InMux I__13630 (
            .O(N__53536),
            .I(N__53494));
    InMux I__13629 (
            .O(N__53535),
            .I(N__53494));
    InMux I__13628 (
            .O(N__53534),
            .I(N__53494));
    InMux I__13627 (
            .O(N__53533),
            .I(N__53489));
    InMux I__13626 (
            .O(N__53532),
            .I(N__53484));
    InMux I__13625 (
            .O(N__53531),
            .I(N__53484));
    Span4Mux_h I__13624 (
            .O(N__53528),
            .I(N__53478));
    InMux I__13623 (
            .O(N__53527),
            .I(N__53475));
    InMux I__13622 (
            .O(N__53526),
            .I(N__53471));
    InMux I__13621 (
            .O(N__53525),
            .I(N__53468));
    InMux I__13620 (
            .O(N__53524),
            .I(N__53457));
    InMux I__13619 (
            .O(N__53523),
            .I(N__53457));
    InMux I__13618 (
            .O(N__53522),
            .I(N__53457));
    InMux I__13617 (
            .O(N__53521),
            .I(N__53457));
    InMux I__13616 (
            .O(N__53520),
            .I(N__53457));
    InMux I__13615 (
            .O(N__53519),
            .I(N__53446));
    InMux I__13614 (
            .O(N__53518),
            .I(N__53446));
    InMux I__13613 (
            .O(N__53517),
            .I(N__53446));
    InMux I__13612 (
            .O(N__53516),
            .I(N__53446));
    InMux I__13611 (
            .O(N__53515),
            .I(N__53446));
    Span4Mux_v I__13610 (
            .O(N__53510),
            .I(N__53439));
    Span4Mux_v I__13609 (
            .O(N__53507),
            .I(N__53439));
    LocalMux I__13608 (
            .O(N__53494),
            .I(N__53439));
    InMux I__13607 (
            .O(N__53493),
            .I(N__53430));
    InMux I__13606 (
            .O(N__53492),
            .I(N__53427));
    LocalMux I__13605 (
            .O(N__53489),
            .I(N__53422));
    LocalMux I__13604 (
            .O(N__53484),
            .I(N__53422));
    InMux I__13603 (
            .O(N__53483),
            .I(N__53417));
    InMux I__13602 (
            .O(N__53482),
            .I(N__53417));
    InMux I__13601 (
            .O(N__53481),
            .I(N__53414));
    Span4Mux_v I__13600 (
            .O(N__53478),
            .I(N__53409));
    LocalMux I__13599 (
            .O(N__53475),
            .I(N__53409));
    InMux I__13598 (
            .O(N__53474),
            .I(N__53399));
    LocalMux I__13597 (
            .O(N__53471),
            .I(N__53394));
    LocalMux I__13596 (
            .O(N__53468),
            .I(N__53394));
    LocalMux I__13595 (
            .O(N__53457),
            .I(N__53385));
    LocalMux I__13594 (
            .O(N__53446),
            .I(N__53385));
    Span4Mux_h I__13593 (
            .O(N__53439),
            .I(N__53382));
    InMux I__13592 (
            .O(N__53438),
            .I(N__53379));
    InMux I__13591 (
            .O(N__53437),
            .I(N__53370));
    InMux I__13590 (
            .O(N__53436),
            .I(N__53370));
    InMux I__13589 (
            .O(N__53435),
            .I(N__53370));
    InMux I__13588 (
            .O(N__53434),
            .I(N__53370));
    InMux I__13587 (
            .O(N__53433),
            .I(N__53367));
    LocalMux I__13586 (
            .O(N__53430),
            .I(N__53362));
    LocalMux I__13585 (
            .O(N__53427),
            .I(N__53362));
    Span4Mux_h I__13584 (
            .O(N__53422),
            .I(N__53357));
    LocalMux I__13583 (
            .O(N__53417),
            .I(N__53357));
    LocalMux I__13582 (
            .O(N__53414),
            .I(N__53349));
    Span4Mux_h I__13581 (
            .O(N__53409),
            .I(N__53349));
    InMux I__13580 (
            .O(N__53408),
            .I(N__53336));
    InMux I__13579 (
            .O(N__53407),
            .I(N__53336));
    InMux I__13578 (
            .O(N__53406),
            .I(N__53336));
    InMux I__13577 (
            .O(N__53405),
            .I(N__53336));
    InMux I__13576 (
            .O(N__53404),
            .I(N__53336));
    InMux I__13575 (
            .O(N__53403),
            .I(N__53336));
    InMux I__13574 (
            .O(N__53402),
            .I(N__53332));
    LocalMux I__13573 (
            .O(N__53399),
            .I(N__53329));
    Span4Mux_h I__13572 (
            .O(N__53394),
            .I(N__53326));
    InMux I__13571 (
            .O(N__53393),
            .I(N__53316));
    InMux I__13570 (
            .O(N__53392),
            .I(N__53316));
    InMux I__13569 (
            .O(N__53391),
            .I(N__53316));
    InMux I__13568 (
            .O(N__53390),
            .I(N__53316));
    Span4Mux_v I__13567 (
            .O(N__53385),
            .I(N__53313));
    Span4Mux_h I__13566 (
            .O(N__53382),
            .I(N__53310));
    LocalMux I__13565 (
            .O(N__53379),
            .I(N__53307));
    LocalMux I__13564 (
            .O(N__53370),
            .I(N__53304));
    LocalMux I__13563 (
            .O(N__53367),
            .I(N__53301));
    Span4Mux_v I__13562 (
            .O(N__53362),
            .I(N__53298));
    Span4Mux_h I__13561 (
            .O(N__53357),
            .I(N__53295));
    InMux I__13560 (
            .O(N__53356),
            .I(N__53290));
    InMux I__13559 (
            .O(N__53355),
            .I(N__53285));
    InMux I__13558 (
            .O(N__53354),
            .I(N__53285));
    Span4Mux_h I__13557 (
            .O(N__53349),
            .I(N__53282));
    LocalMux I__13556 (
            .O(N__53336),
            .I(N__53279));
    InMux I__13555 (
            .O(N__53335),
            .I(N__53272));
    LocalMux I__13554 (
            .O(N__53332),
            .I(N__53269));
    Span4Mux_v I__13553 (
            .O(N__53329),
            .I(N__53264));
    Span4Mux_h I__13552 (
            .O(N__53326),
            .I(N__53264));
    InMux I__13551 (
            .O(N__53325),
            .I(N__53261));
    LocalMux I__13550 (
            .O(N__53316),
            .I(N__53258));
    Span4Mux_h I__13549 (
            .O(N__53313),
            .I(N__53253));
    Span4Mux_h I__13548 (
            .O(N__53310),
            .I(N__53253));
    Span4Mux_h I__13547 (
            .O(N__53307),
            .I(N__53248));
    Span4Mux_h I__13546 (
            .O(N__53304),
            .I(N__53248));
    Span4Mux_h I__13545 (
            .O(N__53301),
            .I(N__53243));
    Span4Mux_h I__13544 (
            .O(N__53298),
            .I(N__53243));
    Span4Mux_v I__13543 (
            .O(N__53295),
            .I(N__53240));
    InMux I__13542 (
            .O(N__53294),
            .I(N__53237));
    InMux I__13541 (
            .O(N__53293),
            .I(N__53234));
    LocalMux I__13540 (
            .O(N__53290),
            .I(N__53229));
    LocalMux I__13539 (
            .O(N__53285),
            .I(N__53229));
    Span4Mux_h I__13538 (
            .O(N__53282),
            .I(N__53224));
    Span4Mux_h I__13537 (
            .O(N__53279),
            .I(N__53224));
    InMux I__13536 (
            .O(N__53278),
            .I(N__53216));
    InMux I__13535 (
            .O(N__53277),
            .I(N__53213));
    InMux I__13534 (
            .O(N__53276),
            .I(N__53210));
    InMux I__13533 (
            .O(N__53275),
            .I(N__53207));
    LocalMux I__13532 (
            .O(N__53272),
            .I(N__53204));
    Span4Mux_h I__13531 (
            .O(N__53269),
            .I(N__53199));
    Span4Mux_h I__13530 (
            .O(N__53264),
            .I(N__53199));
    LocalMux I__13529 (
            .O(N__53261),
            .I(N__53192));
    Span12Mux_h I__13528 (
            .O(N__53258),
            .I(N__53192));
    Sp12to4 I__13527 (
            .O(N__53253),
            .I(N__53192));
    Span4Mux_h I__13526 (
            .O(N__53248),
            .I(N__53185));
    Span4Mux_h I__13525 (
            .O(N__53243),
            .I(N__53185));
    Span4Mux_h I__13524 (
            .O(N__53240),
            .I(N__53185));
    LocalMux I__13523 (
            .O(N__53237),
            .I(N__53176));
    LocalMux I__13522 (
            .O(N__53234),
            .I(N__53176));
    Span4Mux_h I__13521 (
            .O(N__53229),
            .I(N__53176));
    Span4Mux_h I__13520 (
            .O(N__53224),
            .I(N__53176));
    InMux I__13519 (
            .O(N__53223),
            .I(N__53165));
    InMux I__13518 (
            .O(N__53222),
            .I(N__53165));
    InMux I__13517 (
            .O(N__53221),
            .I(N__53165));
    InMux I__13516 (
            .O(N__53220),
            .I(N__53165));
    InMux I__13515 (
            .O(N__53219),
            .I(N__53165));
    LocalMux I__13514 (
            .O(N__53216),
            .I(adc_state_0_adj_1044));
    LocalMux I__13513 (
            .O(N__53213),
            .I(adc_state_0_adj_1044));
    LocalMux I__13512 (
            .O(N__53210),
            .I(adc_state_0_adj_1044));
    LocalMux I__13511 (
            .O(N__53207),
            .I(adc_state_0_adj_1044));
    Odrv12 I__13510 (
            .O(N__53204),
            .I(adc_state_0_adj_1044));
    Odrv4 I__13509 (
            .O(N__53199),
            .I(adc_state_0_adj_1044));
    Odrv12 I__13508 (
            .O(N__53192),
            .I(adc_state_0_adj_1044));
    Odrv4 I__13507 (
            .O(N__53185),
            .I(adc_state_0_adj_1044));
    Odrv4 I__13506 (
            .O(N__53176),
            .I(adc_state_0_adj_1044));
    LocalMux I__13505 (
            .O(N__53165),
            .I(adc_state_0_adj_1044));
    InMux I__13504 (
            .O(N__53144),
            .I(N__53140));
    InMux I__13503 (
            .O(N__53143),
            .I(N__53137));
    LocalMux I__13502 (
            .O(N__53140),
            .I(N__53134));
    LocalMux I__13501 (
            .O(N__53137),
            .I(buf_adcdata2_14));
    Odrv4 I__13500 (
            .O(N__53134),
            .I(buf_adcdata2_14));
    InMux I__13499 (
            .O(N__53129),
            .I(N__53118));
    InMux I__13498 (
            .O(N__53128),
            .I(N__53118));
    InMux I__13497 (
            .O(N__53127),
            .I(N__53107));
    InMux I__13496 (
            .O(N__53126),
            .I(N__53107));
    InMux I__13495 (
            .O(N__53125),
            .I(N__53107));
    InMux I__13494 (
            .O(N__53124),
            .I(N__53102));
    InMux I__13493 (
            .O(N__53123),
            .I(N__53102));
    LocalMux I__13492 (
            .O(N__53118),
            .I(N__53098));
    InMux I__13491 (
            .O(N__53117),
            .I(N__53095));
    InMux I__13490 (
            .O(N__53116),
            .I(N__53092));
    InMux I__13489 (
            .O(N__53115),
            .I(N__53089));
    InMux I__13488 (
            .O(N__53114),
            .I(N__53086));
    LocalMux I__13487 (
            .O(N__53107),
            .I(N__53079));
    LocalMux I__13486 (
            .O(N__53102),
            .I(N__53079));
    InMux I__13485 (
            .O(N__53101),
            .I(N__53072));
    Span4Mux_v I__13484 (
            .O(N__53098),
            .I(N__53065));
    LocalMux I__13483 (
            .O(N__53095),
            .I(N__53065));
    LocalMux I__13482 (
            .O(N__53092),
            .I(N__53065));
    LocalMux I__13481 (
            .O(N__53089),
            .I(N__53060));
    LocalMux I__13480 (
            .O(N__53086),
            .I(N__53057));
    InMux I__13479 (
            .O(N__53085),
            .I(N__53052));
    InMux I__13478 (
            .O(N__53084),
            .I(N__53052));
    Span4Mux_v I__13477 (
            .O(N__53079),
            .I(N__53046));
    InMux I__13476 (
            .O(N__53078),
            .I(N__53037));
    InMux I__13475 (
            .O(N__53077),
            .I(N__53037));
    InMux I__13474 (
            .O(N__53076),
            .I(N__53037));
    InMux I__13473 (
            .O(N__53075),
            .I(N__53037));
    LocalMux I__13472 (
            .O(N__53072),
            .I(N__53034));
    Span4Mux_v I__13471 (
            .O(N__53065),
            .I(N__53031));
    InMux I__13470 (
            .O(N__53064),
            .I(N__53028));
    InMux I__13469 (
            .O(N__53063),
            .I(N__53025));
    Span4Mux_v I__13468 (
            .O(N__53060),
            .I(N__53022));
    Span4Mux_h I__13467 (
            .O(N__53057),
            .I(N__53019));
    LocalMux I__13466 (
            .O(N__53052),
            .I(N__53016));
    InMux I__13465 (
            .O(N__53051),
            .I(N__53012));
    InMux I__13464 (
            .O(N__53050),
            .I(N__53009));
    InMux I__13463 (
            .O(N__53049),
            .I(N__53006));
    Span4Mux_h I__13462 (
            .O(N__53046),
            .I(N__53001));
    LocalMux I__13461 (
            .O(N__53037),
            .I(N__53001));
    Span4Mux_v I__13460 (
            .O(N__53034),
            .I(N__52998));
    Span4Mux_h I__13459 (
            .O(N__53031),
            .I(N__52995));
    LocalMux I__13458 (
            .O(N__53028),
            .I(N__52990));
    LocalMux I__13457 (
            .O(N__53025),
            .I(N__52990));
    Span4Mux_h I__13456 (
            .O(N__53022),
            .I(N__52987));
    Span4Mux_h I__13455 (
            .O(N__53019),
            .I(N__52984));
    Span4Mux_h I__13454 (
            .O(N__53016),
            .I(N__52981));
    InMux I__13453 (
            .O(N__53015),
            .I(N__52978));
    LocalMux I__13452 (
            .O(N__53012),
            .I(N__52969));
    LocalMux I__13451 (
            .O(N__53009),
            .I(N__52969));
    LocalMux I__13450 (
            .O(N__53006),
            .I(N__52969));
    Span4Mux_h I__13449 (
            .O(N__53001),
            .I(N__52969));
    Sp12to4 I__13448 (
            .O(N__52998),
            .I(N__52966));
    Sp12to4 I__13447 (
            .O(N__52995),
            .I(N__52963));
    Span4Mux_v I__13446 (
            .O(N__52990),
            .I(N__52956));
    Span4Mux_h I__13445 (
            .O(N__52987),
            .I(N__52956));
    Span4Mux_h I__13444 (
            .O(N__52984),
            .I(N__52956));
    Span4Mux_h I__13443 (
            .O(N__52981),
            .I(N__52953));
    LocalMux I__13442 (
            .O(N__52978),
            .I(N__52944));
    Sp12to4 I__13441 (
            .O(N__52969),
            .I(N__52944));
    Span12Mux_h I__13440 (
            .O(N__52966),
            .I(N__52944));
    Span12Mux_h I__13439 (
            .O(N__52963),
            .I(N__52944));
    Span4Mux_h I__13438 (
            .O(N__52956),
            .I(N__52941));
    Odrv4 I__13437 (
            .O(N__52953),
            .I(n15153));
    Odrv12 I__13436 (
            .O(N__52944),
            .I(n15153));
    Odrv4 I__13435 (
            .O(N__52941),
            .I(n15153));
    CascadeMux I__13434 (
            .O(N__52934),
            .I(N__52931));
    InMux I__13433 (
            .O(N__52931),
            .I(N__52928));
    LocalMux I__13432 (
            .O(N__52928),
            .I(N__52925));
    Span4Mux_h I__13431 (
            .O(N__52925),
            .I(N__52922));
    Span4Mux_h I__13430 (
            .O(N__52922),
            .I(N__52918));
    CascadeMux I__13429 (
            .O(N__52921),
            .I(N__52914));
    Span4Mux_h I__13428 (
            .O(N__52918),
            .I(N__52911));
    InMux I__13427 (
            .O(N__52917),
            .I(N__52908));
    InMux I__13426 (
            .O(N__52914),
            .I(N__52905));
    Odrv4 I__13425 (
            .O(N__52911),
            .I(cmd_rdadctmp_18));
    LocalMux I__13424 (
            .O(N__52908),
            .I(cmd_rdadctmp_18));
    LocalMux I__13423 (
            .O(N__52905),
            .I(cmd_rdadctmp_18));
    CascadeMux I__13422 (
            .O(N__52898),
            .I(N__52885));
    InMux I__13421 (
            .O(N__52897),
            .I(N__52871));
    InMux I__13420 (
            .O(N__52896),
            .I(N__52868));
    InMux I__13419 (
            .O(N__52895),
            .I(N__52863));
    InMux I__13418 (
            .O(N__52894),
            .I(N__52863));
    InMux I__13417 (
            .O(N__52893),
            .I(N__52860));
    InMux I__13416 (
            .O(N__52892),
            .I(N__52857));
    CascadeMux I__13415 (
            .O(N__52891),
            .I(N__52854));
    CascadeMux I__13414 (
            .O(N__52890),
            .I(N__52841));
    CascadeMux I__13413 (
            .O(N__52889),
            .I(N__52838));
    InMux I__13412 (
            .O(N__52888),
            .I(N__52814));
    InMux I__13411 (
            .O(N__52885),
            .I(N__52814));
    InMux I__13410 (
            .O(N__52884),
            .I(N__52814));
    InMux I__13409 (
            .O(N__52883),
            .I(N__52814));
    InMux I__13408 (
            .O(N__52882),
            .I(N__52814));
    InMux I__13407 (
            .O(N__52881),
            .I(N__52814));
    InMux I__13406 (
            .O(N__52880),
            .I(N__52814));
    InMux I__13405 (
            .O(N__52879),
            .I(N__52814));
    CascadeMux I__13404 (
            .O(N__52878),
            .I(N__52810));
    InMux I__13403 (
            .O(N__52877),
            .I(N__52806));
    InMux I__13402 (
            .O(N__52876),
            .I(N__52799));
    InMux I__13401 (
            .O(N__52875),
            .I(N__52799));
    InMux I__13400 (
            .O(N__52874),
            .I(N__52799));
    LocalMux I__13399 (
            .O(N__52871),
            .I(N__52790));
    LocalMux I__13398 (
            .O(N__52868),
            .I(N__52785));
    LocalMux I__13397 (
            .O(N__52863),
            .I(N__52785));
    LocalMux I__13396 (
            .O(N__52860),
            .I(N__52782));
    LocalMux I__13395 (
            .O(N__52857),
            .I(N__52779));
    InMux I__13394 (
            .O(N__52854),
            .I(N__52775));
    InMux I__13393 (
            .O(N__52853),
            .I(N__52763));
    InMux I__13392 (
            .O(N__52852),
            .I(N__52763));
    InMux I__13391 (
            .O(N__52851),
            .I(N__52763));
    InMux I__13390 (
            .O(N__52850),
            .I(N__52763));
    InMux I__13389 (
            .O(N__52849),
            .I(N__52763));
    InMux I__13388 (
            .O(N__52848),
            .I(N__52760));
    InMux I__13387 (
            .O(N__52847),
            .I(N__52757));
    InMux I__13386 (
            .O(N__52846),
            .I(N__52754));
    InMux I__13385 (
            .O(N__52845),
            .I(N__52751));
    InMux I__13384 (
            .O(N__52844),
            .I(N__52748));
    InMux I__13383 (
            .O(N__52841),
            .I(N__52745));
    InMux I__13382 (
            .O(N__52838),
            .I(N__52742));
    InMux I__13381 (
            .O(N__52837),
            .I(N__52739));
    InMux I__13380 (
            .O(N__52836),
            .I(N__52736));
    InMux I__13379 (
            .O(N__52835),
            .I(N__52725));
    InMux I__13378 (
            .O(N__52834),
            .I(N__52725));
    InMux I__13377 (
            .O(N__52833),
            .I(N__52725));
    InMux I__13376 (
            .O(N__52832),
            .I(N__52725));
    InMux I__13375 (
            .O(N__52831),
            .I(N__52725));
    LocalMux I__13374 (
            .O(N__52814),
            .I(N__52722));
    InMux I__13373 (
            .O(N__52813),
            .I(N__52719));
    InMux I__13372 (
            .O(N__52810),
            .I(N__52714));
    InMux I__13371 (
            .O(N__52809),
            .I(N__52714));
    LocalMux I__13370 (
            .O(N__52806),
            .I(N__52711));
    LocalMux I__13369 (
            .O(N__52799),
            .I(N__52708));
    InMux I__13368 (
            .O(N__52798),
            .I(N__52699));
    InMux I__13367 (
            .O(N__52797),
            .I(N__52699));
    InMux I__13366 (
            .O(N__52796),
            .I(N__52699));
    InMux I__13365 (
            .O(N__52795),
            .I(N__52699));
    InMux I__13364 (
            .O(N__52794),
            .I(N__52696));
    InMux I__13363 (
            .O(N__52793),
            .I(N__52693));
    Span4Mux_v I__13362 (
            .O(N__52790),
            .I(N__52690));
    Span4Mux_v I__13361 (
            .O(N__52785),
            .I(N__52683));
    Span4Mux_v I__13360 (
            .O(N__52782),
            .I(N__52683));
    Span4Mux_v I__13359 (
            .O(N__52779),
            .I(N__52683));
    CascadeMux I__13358 (
            .O(N__52778),
            .I(N__52680));
    LocalMux I__13357 (
            .O(N__52775),
            .I(N__52667));
    InMux I__13356 (
            .O(N__52774),
            .I(N__52664));
    LocalMux I__13355 (
            .O(N__52763),
            .I(N__52659));
    LocalMux I__13354 (
            .O(N__52760),
            .I(N__52659));
    LocalMux I__13353 (
            .O(N__52757),
            .I(N__52656));
    LocalMux I__13352 (
            .O(N__52754),
            .I(N__52653));
    LocalMux I__13351 (
            .O(N__52751),
            .I(N__52650));
    LocalMux I__13350 (
            .O(N__52748),
            .I(N__52645));
    LocalMux I__13349 (
            .O(N__52745),
            .I(N__52645));
    LocalMux I__13348 (
            .O(N__52742),
            .I(N__52636));
    LocalMux I__13347 (
            .O(N__52739),
            .I(N__52636));
    LocalMux I__13346 (
            .O(N__52736),
            .I(N__52636));
    LocalMux I__13345 (
            .O(N__52725),
            .I(N__52636));
    Span4Mux_h I__13344 (
            .O(N__52722),
            .I(N__52631));
    LocalMux I__13343 (
            .O(N__52719),
            .I(N__52631));
    LocalMux I__13342 (
            .O(N__52714),
            .I(N__52628));
    Span4Mux_v I__13341 (
            .O(N__52711),
            .I(N__52621));
    Span4Mux_v I__13340 (
            .O(N__52708),
            .I(N__52621));
    LocalMux I__13339 (
            .O(N__52699),
            .I(N__52621));
    LocalMux I__13338 (
            .O(N__52696),
            .I(N__52607));
    LocalMux I__13337 (
            .O(N__52693),
            .I(N__52607));
    Sp12to4 I__13336 (
            .O(N__52690),
            .I(N__52607));
    Sp12to4 I__13335 (
            .O(N__52683),
            .I(N__52607));
    InMux I__13334 (
            .O(N__52680),
            .I(N__52598));
    InMux I__13333 (
            .O(N__52679),
            .I(N__52598));
    InMux I__13332 (
            .O(N__52678),
            .I(N__52595));
    InMux I__13331 (
            .O(N__52677),
            .I(N__52578));
    InMux I__13330 (
            .O(N__52676),
            .I(N__52578));
    InMux I__13329 (
            .O(N__52675),
            .I(N__52578));
    InMux I__13328 (
            .O(N__52674),
            .I(N__52578));
    InMux I__13327 (
            .O(N__52673),
            .I(N__52578));
    InMux I__13326 (
            .O(N__52672),
            .I(N__52578));
    InMux I__13325 (
            .O(N__52671),
            .I(N__52578));
    InMux I__13324 (
            .O(N__52670),
            .I(N__52578));
    Span4Mux_h I__13323 (
            .O(N__52667),
            .I(N__52571));
    LocalMux I__13322 (
            .O(N__52664),
            .I(N__52571));
    Span4Mux_v I__13321 (
            .O(N__52659),
            .I(N__52571));
    Span4Mux_v I__13320 (
            .O(N__52656),
            .I(N__52564));
    Span4Mux_v I__13319 (
            .O(N__52653),
            .I(N__52564));
    Span4Mux_v I__13318 (
            .O(N__52650),
            .I(N__52564));
    Span4Mux_h I__13317 (
            .O(N__52645),
            .I(N__52559));
    Span4Mux_h I__13316 (
            .O(N__52636),
            .I(N__52559));
    Span4Mux_v I__13315 (
            .O(N__52631),
            .I(N__52552));
    Span4Mux_v I__13314 (
            .O(N__52628),
            .I(N__52552));
    Span4Mux_v I__13313 (
            .O(N__52621),
            .I(N__52552));
    InMux I__13312 (
            .O(N__52620),
            .I(N__52545));
    InMux I__13311 (
            .O(N__52619),
            .I(N__52545));
    InMux I__13310 (
            .O(N__52618),
            .I(N__52545));
    InMux I__13309 (
            .O(N__52617),
            .I(N__52540));
    InMux I__13308 (
            .O(N__52616),
            .I(N__52540));
    Span12Mux_h I__13307 (
            .O(N__52607),
            .I(N__52537));
    InMux I__13306 (
            .O(N__52606),
            .I(N__52528));
    InMux I__13305 (
            .O(N__52605),
            .I(N__52528));
    InMux I__13304 (
            .O(N__52604),
            .I(N__52528));
    InMux I__13303 (
            .O(N__52603),
            .I(N__52528));
    LocalMux I__13302 (
            .O(N__52598),
            .I(adc_state_0));
    LocalMux I__13301 (
            .O(N__52595),
            .I(adc_state_0));
    LocalMux I__13300 (
            .O(N__52578),
            .I(adc_state_0));
    Odrv4 I__13299 (
            .O(N__52571),
            .I(adc_state_0));
    Odrv4 I__13298 (
            .O(N__52564),
            .I(adc_state_0));
    Odrv4 I__13297 (
            .O(N__52559),
            .I(adc_state_0));
    Odrv4 I__13296 (
            .O(N__52552),
            .I(adc_state_0));
    LocalMux I__13295 (
            .O(N__52545),
            .I(adc_state_0));
    LocalMux I__13294 (
            .O(N__52540),
            .I(adc_state_0));
    Odrv12 I__13293 (
            .O(N__52537),
            .I(adc_state_0));
    LocalMux I__13292 (
            .O(N__52528),
            .I(adc_state_0));
    InMux I__13291 (
            .O(N__52505),
            .I(N__52501));
    InMux I__13290 (
            .O(N__52504),
            .I(N__52498));
    LocalMux I__13289 (
            .O(N__52501),
            .I(N__52495));
    LocalMux I__13288 (
            .O(N__52498),
            .I(buf_adcdata1_10));
    Odrv4 I__13287 (
            .O(N__52495),
            .I(buf_adcdata1_10));
    InMux I__13286 (
            .O(N__52490),
            .I(N__52486));
    CascadeMux I__13285 (
            .O(N__52489),
            .I(N__52483));
    LocalMux I__13284 (
            .O(N__52486),
            .I(N__52480));
    InMux I__13283 (
            .O(N__52483),
            .I(N__52477));
    Span12Mux_s11_v I__13282 (
            .O(N__52480),
            .I(N__52474));
    LocalMux I__13281 (
            .O(N__52477),
            .I(n8_adj_1225));
    Odrv12 I__13280 (
            .O(N__52474),
            .I(n8_adj_1225));
    InMux I__13279 (
            .O(N__52469),
            .I(N__52463));
    InMux I__13278 (
            .O(N__52468),
            .I(N__52439));
    InMux I__13277 (
            .O(N__52467),
            .I(N__52436));
    InMux I__13276 (
            .O(N__52466),
            .I(N__52427));
    LocalMux I__13275 (
            .O(N__52463),
            .I(N__52420));
    CascadeMux I__13274 (
            .O(N__52462),
            .I(N__52415));
    CascadeMux I__13273 (
            .O(N__52461),
            .I(N__52411));
    CascadeMux I__13272 (
            .O(N__52460),
            .I(N__52407));
    CascadeMux I__13271 (
            .O(N__52459),
            .I(N__52403));
    CascadeMux I__13270 (
            .O(N__52458),
            .I(N__52399));
    CascadeMux I__13269 (
            .O(N__52457),
            .I(N__52395));
    CascadeMux I__13268 (
            .O(N__52456),
            .I(N__52391));
    InMux I__13267 (
            .O(N__52455),
            .I(N__52387));
    CascadeMux I__13266 (
            .O(N__52454),
            .I(N__52381));
    InMux I__13265 (
            .O(N__52453),
            .I(N__52377));
    InMux I__13264 (
            .O(N__52452),
            .I(N__52369));
    InMux I__13263 (
            .O(N__52451),
            .I(N__52369));
    InMux I__13262 (
            .O(N__52450),
            .I(N__52369));
    InMux I__13261 (
            .O(N__52449),
            .I(N__52364));
    InMux I__13260 (
            .O(N__52448),
            .I(N__52364));
    CascadeMux I__13259 (
            .O(N__52447),
            .I(N__52361));
    CascadeMux I__13258 (
            .O(N__52446),
            .I(N__52357));
    InMux I__13257 (
            .O(N__52445),
            .I(N__52351));
    InMux I__13256 (
            .O(N__52444),
            .I(N__52351));
    InMux I__13255 (
            .O(N__52443),
            .I(N__52346));
    InMux I__13254 (
            .O(N__52442),
            .I(N__52342));
    LocalMux I__13253 (
            .O(N__52439),
            .I(N__52337));
    LocalMux I__13252 (
            .O(N__52436),
            .I(N__52337));
    InMux I__13251 (
            .O(N__52435),
            .I(N__52332));
    InMux I__13250 (
            .O(N__52434),
            .I(N__52332));
    InMux I__13249 (
            .O(N__52433),
            .I(N__52327));
    InMux I__13248 (
            .O(N__52432),
            .I(N__52327));
    InMux I__13247 (
            .O(N__52431),
            .I(N__52322));
    InMux I__13246 (
            .O(N__52430),
            .I(N__52322));
    LocalMux I__13245 (
            .O(N__52427),
            .I(N__52319));
    InMux I__13244 (
            .O(N__52426),
            .I(N__52314));
    InMux I__13243 (
            .O(N__52425),
            .I(N__52314));
    SRMux I__13242 (
            .O(N__52424),
            .I(N__52306));
    CascadeMux I__13241 (
            .O(N__52423),
            .I(N__52303));
    Span4Mux_h I__13240 (
            .O(N__52420),
            .I(N__52297));
    InMux I__13239 (
            .O(N__52419),
            .I(N__52280));
    InMux I__13238 (
            .O(N__52418),
            .I(N__52280));
    InMux I__13237 (
            .O(N__52415),
            .I(N__52280));
    InMux I__13236 (
            .O(N__52414),
            .I(N__52280));
    InMux I__13235 (
            .O(N__52411),
            .I(N__52280));
    InMux I__13234 (
            .O(N__52410),
            .I(N__52280));
    InMux I__13233 (
            .O(N__52407),
            .I(N__52280));
    InMux I__13232 (
            .O(N__52406),
            .I(N__52280));
    InMux I__13231 (
            .O(N__52403),
            .I(N__52265));
    InMux I__13230 (
            .O(N__52402),
            .I(N__52265));
    InMux I__13229 (
            .O(N__52399),
            .I(N__52265));
    InMux I__13228 (
            .O(N__52398),
            .I(N__52265));
    InMux I__13227 (
            .O(N__52395),
            .I(N__52265));
    InMux I__13226 (
            .O(N__52394),
            .I(N__52265));
    InMux I__13225 (
            .O(N__52391),
            .I(N__52265));
    CascadeMux I__13224 (
            .O(N__52390),
            .I(N__52262));
    LocalMux I__13223 (
            .O(N__52387),
            .I(N__52259));
    InMux I__13222 (
            .O(N__52386),
            .I(N__52254));
    InMux I__13221 (
            .O(N__52385),
            .I(N__52254));
    InMux I__13220 (
            .O(N__52384),
            .I(N__52247));
    InMux I__13219 (
            .O(N__52381),
            .I(N__52247));
    InMux I__13218 (
            .O(N__52380),
            .I(N__52247));
    LocalMux I__13217 (
            .O(N__52377),
            .I(N__52244));
    InMux I__13216 (
            .O(N__52376),
            .I(N__52241));
    LocalMux I__13215 (
            .O(N__52369),
            .I(N__52233));
    LocalMux I__13214 (
            .O(N__52364),
            .I(N__52233));
    InMux I__13213 (
            .O(N__52361),
            .I(N__52230));
    InMux I__13212 (
            .O(N__52360),
            .I(N__52225));
    InMux I__13211 (
            .O(N__52357),
            .I(N__52225));
    CascadeMux I__13210 (
            .O(N__52356),
            .I(N__52222));
    LocalMux I__13209 (
            .O(N__52351),
            .I(N__52214));
    InMux I__13208 (
            .O(N__52350),
            .I(N__52211));
    InMux I__13207 (
            .O(N__52349),
            .I(N__52208));
    LocalMux I__13206 (
            .O(N__52346),
            .I(N__52205));
    InMux I__13205 (
            .O(N__52345),
            .I(N__52202));
    LocalMux I__13204 (
            .O(N__52342),
            .I(N__52187));
    Span4Mux_v I__13203 (
            .O(N__52337),
            .I(N__52187));
    LocalMux I__13202 (
            .O(N__52332),
            .I(N__52187));
    LocalMux I__13201 (
            .O(N__52327),
            .I(N__52187));
    LocalMux I__13200 (
            .O(N__52322),
            .I(N__52187));
    Span4Mux_h I__13199 (
            .O(N__52319),
            .I(N__52187));
    LocalMux I__13198 (
            .O(N__52314),
            .I(N__52187));
    InMux I__13197 (
            .O(N__52313),
            .I(N__52172));
    InMux I__13196 (
            .O(N__52312),
            .I(N__52172));
    InMux I__13195 (
            .O(N__52311),
            .I(N__52172));
    InMux I__13194 (
            .O(N__52310),
            .I(N__52172));
    InMux I__13193 (
            .O(N__52309),
            .I(N__52172));
    LocalMux I__13192 (
            .O(N__52306),
            .I(N__52169));
    InMux I__13191 (
            .O(N__52303),
            .I(N__52166));
    InMux I__13190 (
            .O(N__52302),
            .I(N__52162));
    InMux I__13189 (
            .O(N__52301),
            .I(N__52159));
    InMux I__13188 (
            .O(N__52300),
            .I(N__52156));
    Span4Mux_v I__13187 (
            .O(N__52297),
            .I(N__52149));
    LocalMux I__13186 (
            .O(N__52280),
            .I(N__52149));
    LocalMux I__13185 (
            .O(N__52265),
            .I(N__52149));
    InMux I__13184 (
            .O(N__52262),
            .I(N__52146));
    Span4Mux_v I__13183 (
            .O(N__52259),
            .I(N__52143));
    LocalMux I__13182 (
            .O(N__52254),
            .I(N__52140));
    LocalMux I__13181 (
            .O(N__52247),
            .I(N__52133));
    Span4Mux_h I__13180 (
            .O(N__52244),
            .I(N__52133));
    LocalMux I__13179 (
            .O(N__52241),
            .I(N__52133));
    InMux I__13178 (
            .O(N__52240),
            .I(N__52126));
    InMux I__13177 (
            .O(N__52239),
            .I(N__52126));
    InMux I__13176 (
            .O(N__52238),
            .I(N__52126));
    Span4Mux_h I__13175 (
            .O(N__52233),
            .I(N__52119));
    LocalMux I__13174 (
            .O(N__52230),
            .I(N__52119));
    LocalMux I__13173 (
            .O(N__52225),
            .I(N__52119));
    InMux I__13172 (
            .O(N__52222),
            .I(N__52110));
    InMux I__13171 (
            .O(N__52221),
            .I(N__52110));
    InMux I__13170 (
            .O(N__52220),
            .I(N__52110));
    InMux I__13169 (
            .O(N__52219),
            .I(N__52110));
    InMux I__13168 (
            .O(N__52218),
            .I(N__52105));
    InMux I__13167 (
            .O(N__52217),
            .I(N__52105));
    Span4Mux_h I__13166 (
            .O(N__52214),
            .I(N__52102));
    LocalMux I__13165 (
            .O(N__52211),
            .I(N__52091));
    LocalMux I__13164 (
            .O(N__52208),
            .I(N__52091));
    Span4Mux_h I__13163 (
            .O(N__52205),
            .I(N__52091));
    LocalMux I__13162 (
            .O(N__52202),
            .I(N__52091));
    Span4Mux_v I__13161 (
            .O(N__52187),
            .I(N__52091));
    InMux I__13160 (
            .O(N__52186),
            .I(N__52086));
    InMux I__13159 (
            .O(N__52185),
            .I(N__52086));
    InMux I__13158 (
            .O(N__52184),
            .I(N__52083));
    InMux I__13157 (
            .O(N__52183),
            .I(N__52078));
    LocalMux I__13156 (
            .O(N__52172),
            .I(N__52075));
    Span4Mux_v I__13155 (
            .O(N__52169),
            .I(N__52070));
    LocalMux I__13154 (
            .O(N__52166),
            .I(N__52067));
    CascadeMux I__13153 (
            .O(N__52165),
            .I(N__52063));
    LocalMux I__13152 (
            .O(N__52162),
            .I(N__52058));
    LocalMux I__13151 (
            .O(N__52159),
            .I(N__52051));
    LocalMux I__13150 (
            .O(N__52156),
            .I(N__52051));
    Span4Mux_v I__13149 (
            .O(N__52149),
            .I(N__52051));
    LocalMux I__13148 (
            .O(N__52146),
            .I(N__52046));
    Span4Mux_v I__13147 (
            .O(N__52143),
            .I(N__52046));
    Span4Mux_h I__13146 (
            .O(N__52140),
            .I(N__52039));
    Span4Mux_v I__13145 (
            .O(N__52133),
            .I(N__52039));
    LocalMux I__13144 (
            .O(N__52126),
            .I(N__52039));
    Span4Mux_h I__13143 (
            .O(N__52119),
            .I(N__52034));
    LocalMux I__13142 (
            .O(N__52110),
            .I(N__52034));
    LocalMux I__13141 (
            .O(N__52105),
            .I(N__52025));
    Span4Mux_h I__13140 (
            .O(N__52102),
            .I(N__52025));
    Span4Mux_v I__13139 (
            .O(N__52091),
            .I(N__52025));
    LocalMux I__13138 (
            .O(N__52086),
            .I(N__52022));
    LocalMux I__13137 (
            .O(N__52083),
            .I(N__52019));
    InMux I__13136 (
            .O(N__52082),
            .I(N__52016));
    InMux I__13135 (
            .O(N__52081),
            .I(N__52013));
    LocalMux I__13134 (
            .O(N__52078),
            .I(N__52010));
    Span12Mux_v I__13133 (
            .O(N__52075),
            .I(N__52007));
    InMux I__13132 (
            .O(N__52074),
            .I(N__52004));
    InMux I__13131 (
            .O(N__52073),
            .I(N__52001));
    Span4Mux_h I__13130 (
            .O(N__52070),
            .I(N__51996));
    Span4Mux_v I__13129 (
            .O(N__52067),
            .I(N__51996));
    InMux I__13128 (
            .O(N__52066),
            .I(N__51991));
    InMux I__13127 (
            .O(N__52063),
            .I(N__51991));
    InMux I__13126 (
            .O(N__52062),
            .I(N__51986));
    InMux I__13125 (
            .O(N__52061),
            .I(N__51986));
    Span4Mux_v I__13124 (
            .O(N__52058),
            .I(N__51977));
    Span4Mux_v I__13123 (
            .O(N__52051),
            .I(N__51977));
    Span4Mux_v I__13122 (
            .O(N__52046),
            .I(N__51977));
    Span4Mux_h I__13121 (
            .O(N__52039),
            .I(N__51977));
    Span4Mux_h I__13120 (
            .O(N__52034),
            .I(N__51974));
    InMux I__13119 (
            .O(N__52033),
            .I(N__51969));
    InMux I__13118 (
            .O(N__52032),
            .I(N__51969));
    Span4Mux_h I__13117 (
            .O(N__52025),
            .I(N__51964));
    Span4Mux_h I__13116 (
            .O(N__52022),
            .I(N__51964));
    Span12Mux_h I__13115 (
            .O(N__52019),
            .I(N__51953));
    LocalMux I__13114 (
            .O(N__52016),
            .I(N__51953));
    LocalMux I__13113 (
            .O(N__52013),
            .I(N__51953));
    Span12Mux_s10_v I__13112 (
            .O(N__52010),
            .I(N__51953));
    Span12Mux_h I__13111 (
            .O(N__52007),
            .I(N__51953));
    LocalMux I__13110 (
            .O(N__52004),
            .I(comm_state_3));
    LocalMux I__13109 (
            .O(N__52001),
            .I(comm_state_3));
    Odrv4 I__13108 (
            .O(N__51996),
            .I(comm_state_3));
    LocalMux I__13107 (
            .O(N__51991),
            .I(comm_state_3));
    LocalMux I__13106 (
            .O(N__51986),
            .I(comm_state_3));
    Odrv4 I__13105 (
            .O(N__51977),
            .I(comm_state_3));
    Odrv4 I__13104 (
            .O(N__51974),
            .I(comm_state_3));
    LocalMux I__13103 (
            .O(N__51969),
            .I(comm_state_3));
    Odrv4 I__13102 (
            .O(N__51964),
            .I(comm_state_3));
    Odrv12 I__13101 (
            .O(N__51953),
            .I(comm_state_3));
    CascadeMux I__13100 (
            .O(N__51932),
            .I(N__51924));
    CascadeMux I__13099 (
            .O(N__51931),
            .I(N__51919));
    CascadeMux I__13098 (
            .O(N__51930),
            .I(N__51910));
    CascadeMux I__13097 (
            .O(N__51929),
            .I(N__51906));
    CascadeMux I__13096 (
            .O(N__51928),
            .I(N__51903));
    InMux I__13095 (
            .O(N__51927),
            .I(N__51900));
    InMux I__13094 (
            .O(N__51924),
            .I(N__51890));
    InMux I__13093 (
            .O(N__51923),
            .I(N__51887));
    InMux I__13092 (
            .O(N__51922),
            .I(N__51884));
    InMux I__13091 (
            .O(N__51919),
            .I(N__51881));
    CascadeMux I__13090 (
            .O(N__51918),
            .I(N__51876));
    CascadeMux I__13089 (
            .O(N__51917),
            .I(N__51873));
    CascadeMux I__13088 (
            .O(N__51916),
            .I(N__51870));
    InMux I__13087 (
            .O(N__51915),
            .I(N__51863));
    CascadeMux I__13086 (
            .O(N__51914),
            .I(N__51860));
    CascadeMux I__13085 (
            .O(N__51913),
            .I(N__51857));
    InMux I__13084 (
            .O(N__51910),
            .I(N__51854));
    CascadeMux I__13083 (
            .O(N__51909),
            .I(N__51848));
    InMux I__13082 (
            .O(N__51906),
            .I(N__51845));
    InMux I__13081 (
            .O(N__51903),
            .I(N__51838));
    LocalMux I__13080 (
            .O(N__51900),
            .I(N__51835));
    InMux I__13079 (
            .O(N__51899),
            .I(N__51830));
    InMux I__13078 (
            .O(N__51898),
            .I(N__51830));
    CascadeMux I__13077 (
            .O(N__51897),
            .I(N__51826));
    InMux I__13076 (
            .O(N__51896),
            .I(N__51822));
    InMux I__13075 (
            .O(N__51895),
            .I(N__51817));
    InMux I__13074 (
            .O(N__51894),
            .I(N__51817));
    InMux I__13073 (
            .O(N__51893),
            .I(N__51814));
    LocalMux I__13072 (
            .O(N__51890),
            .I(N__51811));
    LocalMux I__13071 (
            .O(N__51887),
            .I(N__51808));
    LocalMux I__13070 (
            .O(N__51884),
            .I(N__51805));
    LocalMux I__13069 (
            .O(N__51881),
            .I(N__51802));
    InMux I__13068 (
            .O(N__51880),
            .I(N__51797));
    InMux I__13067 (
            .O(N__51879),
            .I(N__51797));
    InMux I__13066 (
            .O(N__51876),
            .I(N__51794));
    InMux I__13065 (
            .O(N__51873),
            .I(N__51787));
    InMux I__13064 (
            .O(N__51870),
            .I(N__51787));
    InMux I__13063 (
            .O(N__51869),
            .I(N__51787));
    InMux I__13062 (
            .O(N__51868),
            .I(N__51784));
    InMux I__13061 (
            .O(N__51867),
            .I(N__51779));
    InMux I__13060 (
            .O(N__51866),
            .I(N__51779));
    LocalMux I__13059 (
            .O(N__51863),
            .I(N__51776));
    InMux I__13058 (
            .O(N__51860),
            .I(N__51771));
    InMux I__13057 (
            .O(N__51857),
            .I(N__51771));
    LocalMux I__13056 (
            .O(N__51854),
            .I(N__51763));
    InMux I__13055 (
            .O(N__51853),
            .I(N__51758));
    InMux I__13054 (
            .O(N__51852),
            .I(N__51758));
    InMux I__13053 (
            .O(N__51851),
            .I(N__51753));
    InMux I__13052 (
            .O(N__51848),
            .I(N__51753));
    LocalMux I__13051 (
            .O(N__51845),
            .I(N__51750));
    CascadeMux I__13050 (
            .O(N__51844),
            .I(N__51746));
    CascadeMux I__13049 (
            .O(N__51843),
            .I(N__51743));
    CascadeMux I__13048 (
            .O(N__51842),
            .I(N__51740));
    InMux I__13047 (
            .O(N__51841),
            .I(N__51734));
    LocalMux I__13046 (
            .O(N__51838),
            .I(N__51731));
    Span4Mux_h I__13045 (
            .O(N__51835),
            .I(N__51726));
    LocalMux I__13044 (
            .O(N__51830),
            .I(N__51726));
    CascadeMux I__13043 (
            .O(N__51829),
            .I(N__51722));
    InMux I__13042 (
            .O(N__51826),
            .I(N__51719));
    CascadeMux I__13041 (
            .O(N__51825),
            .I(N__51716));
    LocalMux I__13040 (
            .O(N__51822),
            .I(N__51711));
    LocalMux I__13039 (
            .O(N__51817),
            .I(N__51711));
    LocalMux I__13038 (
            .O(N__51814),
            .I(N__51708));
    Span4Mux_v I__13037 (
            .O(N__51811),
            .I(N__51705));
    Span4Mux_v I__13036 (
            .O(N__51808),
            .I(N__51700));
    Span4Mux_v I__13035 (
            .O(N__51805),
            .I(N__51700));
    Span4Mux_v I__13034 (
            .O(N__51802),
            .I(N__51683));
    LocalMux I__13033 (
            .O(N__51797),
            .I(N__51683));
    LocalMux I__13032 (
            .O(N__51794),
            .I(N__51683));
    LocalMux I__13031 (
            .O(N__51787),
            .I(N__51683));
    LocalMux I__13030 (
            .O(N__51784),
            .I(N__51683));
    LocalMux I__13029 (
            .O(N__51779),
            .I(N__51683));
    Span4Mux_v I__13028 (
            .O(N__51776),
            .I(N__51683));
    LocalMux I__13027 (
            .O(N__51771),
            .I(N__51683));
    CascadeMux I__13026 (
            .O(N__51770),
            .I(N__51680));
    CascadeMux I__13025 (
            .O(N__51769),
            .I(N__51676));
    CascadeMux I__13024 (
            .O(N__51768),
            .I(N__51672));
    CascadeMux I__13023 (
            .O(N__51767),
            .I(N__51669));
    CascadeMux I__13022 (
            .O(N__51766),
            .I(N__51665));
    Span4Mux_h I__13021 (
            .O(N__51763),
            .I(N__51658));
    LocalMux I__13020 (
            .O(N__51758),
            .I(N__51658));
    LocalMux I__13019 (
            .O(N__51753),
            .I(N__51655));
    Span4Mux_v I__13018 (
            .O(N__51750),
            .I(N__51652));
    InMux I__13017 (
            .O(N__51749),
            .I(N__51643));
    InMux I__13016 (
            .O(N__51746),
            .I(N__51643));
    InMux I__13015 (
            .O(N__51743),
            .I(N__51643));
    InMux I__13014 (
            .O(N__51740),
            .I(N__51643));
    CascadeMux I__13013 (
            .O(N__51739),
            .I(N__51640));
    CascadeMux I__13012 (
            .O(N__51738),
            .I(N__51637));
    CascadeMux I__13011 (
            .O(N__51737),
            .I(N__51633));
    LocalMux I__13010 (
            .O(N__51734),
            .I(N__51630));
    Span4Mux_h I__13009 (
            .O(N__51731),
            .I(N__51625));
    Span4Mux_h I__13008 (
            .O(N__51726),
            .I(N__51625));
    InMux I__13007 (
            .O(N__51725),
            .I(N__51620));
    InMux I__13006 (
            .O(N__51722),
            .I(N__51620));
    LocalMux I__13005 (
            .O(N__51719),
            .I(N__51617));
    InMux I__13004 (
            .O(N__51716),
            .I(N__51614));
    Span4Mux_v I__13003 (
            .O(N__51711),
            .I(N__51607));
    Span4Mux_v I__13002 (
            .O(N__51708),
            .I(N__51607));
    Span4Mux_v I__13001 (
            .O(N__51705),
            .I(N__51607));
    Span4Mux_v I__13000 (
            .O(N__51700),
            .I(N__51602));
    Span4Mux_v I__12999 (
            .O(N__51683),
            .I(N__51602));
    InMux I__12998 (
            .O(N__51680),
            .I(N__51599));
    InMux I__12997 (
            .O(N__51679),
            .I(N__51594));
    InMux I__12996 (
            .O(N__51676),
            .I(N__51594));
    InMux I__12995 (
            .O(N__51675),
            .I(N__51583));
    InMux I__12994 (
            .O(N__51672),
            .I(N__51583));
    InMux I__12993 (
            .O(N__51669),
            .I(N__51583));
    InMux I__12992 (
            .O(N__51668),
            .I(N__51583));
    InMux I__12991 (
            .O(N__51665),
            .I(N__51583));
    InMux I__12990 (
            .O(N__51664),
            .I(N__51578));
    InMux I__12989 (
            .O(N__51663),
            .I(N__51578));
    Span4Mux_h I__12988 (
            .O(N__51658),
            .I(N__51569));
    Span4Mux_v I__12987 (
            .O(N__51655),
            .I(N__51569));
    Span4Mux_h I__12986 (
            .O(N__51652),
            .I(N__51569));
    LocalMux I__12985 (
            .O(N__51643),
            .I(N__51569));
    InMux I__12984 (
            .O(N__51640),
            .I(N__51566));
    InMux I__12983 (
            .O(N__51637),
            .I(N__51561));
    InMux I__12982 (
            .O(N__51636),
            .I(N__51561));
    InMux I__12981 (
            .O(N__51633),
            .I(N__51558));
    Span12Mux_v I__12980 (
            .O(N__51630),
            .I(N__51555));
    Span4Mux_v I__12979 (
            .O(N__51625),
            .I(N__51550));
    LocalMux I__12978 (
            .O(N__51620),
            .I(N__51550));
    Span12Mux_v I__12977 (
            .O(N__51617),
            .I(N__51541));
    LocalMux I__12976 (
            .O(N__51614),
            .I(N__51541));
    Sp12to4 I__12975 (
            .O(N__51607),
            .I(N__51541));
    Sp12to4 I__12974 (
            .O(N__51602),
            .I(N__51541));
    LocalMux I__12973 (
            .O(N__51599),
            .I(N__51530));
    LocalMux I__12972 (
            .O(N__51594),
            .I(N__51530));
    LocalMux I__12971 (
            .O(N__51583),
            .I(N__51530));
    LocalMux I__12970 (
            .O(N__51578),
            .I(N__51530));
    Span4Mux_v I__12969 (
            .O(N__51569),
            .I(N__51530));
    LocalMux I__12968 (
            .O(N__51566),
            .I(n6791));
    LocalMux I__12967 (
            .O(N__51561),
            .I(n6791));
    LocalMux I__12966 (
            .O(N__51558),
            .I(n6791));
    Odrv12 I__12965 (
            .O(N__51555),
            .I(n6791));
    Odrv4 I__12964 (
            .O(N__51550),
            .I(n6791));
    Odrv12 I__12963 (
            .O(N__51541),
            .I(n6791));
    Odrv4 I__12962 (
            .O(N__51530),
            .I(n6791));
    InMux I__12961 (
            .O(N__51515),
            .I(N__51512));
    LocalMux I__12960 (
            .O(N__51512),
            .I(N__51509));
    Span4Mux_h I__12959 (
            .O(N__51509),
            .I(N__51505));
    InMux I__12958 (
            .O(N__51508),
            .I(N__51502));
    Span4Mux_h I__12957 (
            .O(N__51505),
            .I(N__51499));
    LocalMux I__12956 (
            .O(N__51502),
            .I(n7_adj_1224));
    Odrv4 I__12955 (
            .O(N__51499),
            .I(n7_adj_1224));
    CascadeMux I__12954 (
            .O(N__51494),
            .I(N__51491));
    CascadeBuf I__12953 (
            .O(N__51491),
            .I(N__51488));
    CascadeMux I__12952 (
            .O(N__51488),
            .I(N__51485));
    CascadeBuf I__12951 (
            .O(N__51485),
            .I(N__51482));
    CascadeMux I__12950 (
            .O(N__51482),
            .I(N__51479));
    CascadeBuf I__12949 (
            .O(N__51479),
            .I(N__51476));
    CascadeMux I__12948 (
            .O(N__51476),
            .I(N__51473));
    CascadeBuf I__12947 (
            .O(N__51473),
            .I(N__51470));
    CascadeMux I__12946 (
            .O(N__51470),
            .I(N__51467));
    CascadeBuf I__12945 (
            .O(N__51467),
            .I(N__51464));
    CascadeMux I__12944 (
            .O(N__51464),
            .I(N__51461));
    CascadeBuf I__12943 (
            .O(N__51461),
            .I(N__51457));
    CascadeMux I__12942 (
            .O(N__51460),
            .I(N__51454));
    CascadeMux I__12941 (
            .O(N__51457),
            .I(N__51451));
    CascadeBuf I__12940 (
            .O(N__51454),
            .I(N__51448));
    CascadeBuf I__12939 (
            .O(N__51451),
            .I(N__51445));
    CascadeMux I__12938 (
            .O(N__51448),
            .I(N__51442));
    CascadeMux I__12937 (
            .O(N__51445),
            .I(N__51439));
    InMux I__12936 (
            .O(N__51442),
            .I(N__51436));
    CascadeBuf I__12935 (
            .O(N__51439),
            .I(N__51433));
    LocalMux I__12934 (
            .O(N__51436),
            .I(N__51430));
    CascadeMux I__12933 (
            .O(N__51433),
            .I(N__51427));
    Span12Mux_s11_h I__12932 (
            .O(N__51430),
            .I(N__51424));
    CascadeBuf I__12931 (
            .O(N__51427),
            .I(N__51421));
    Span12Mux_h I__12930 (
            .O(N__51424),
            .I(N__51418));
    CascadeMux I__12929 (
            .O(N__51421),
            .I(N__51415));
    Span12Mux_v I__12928 (
            .O(N__51418),
            .I(N__51412));
    InMux I__12927 (
            .O(N__51415),
            .I(N__51409));
    Odrv12 I__12926 (
            .O(N__51412),
            .I(data_index_9_N_258_5));
    LocalMux I__12925 (
            .O(N__51409),
            .I(data_index_9_N_258_5));
    InMux I__12924 (
            .O(N__51404),
            .I(N__51401));
    LocalMux I__12923 (
            .O(N__51401),
            .I(N__51398));
    Span4Mux_v I__12922 (
            .O(N__51398),
            .I(N__51394));
    InMux I__12921 (
            .O(N__51397),
            .I(N__51391));
    Span4Mux_h I__12920 (
            .O(N__51394),
            .I(N__51385));
    LocalMux I__12919 (
            .O(N__51391),
            .I(N__51385));
    InMux I__12918 (
            .O(N__51390),
            .I(N__51382));
    Span4Mux_v I__12917 (
            .O(N__51385),
            .I(N__51379));
    LocalMux I__12916 (
            .O(N__51382),
            .I(N__51376));
    Span4Mux_h I__12915 (
            .O(N__51379),
            .I(N__51371));
    Span4Mux_h I__12914 (
            .O(N__51376),
            .I(N__51368));
    InMux I__12913 (
            .O(N__51375),
            .I(N__51365));
    InMux I__12912 (
            .O(N__51374),
            .I(N__51362));
    Sp12to4 I__12911 (
            .O(N__51371),
            .I(N__51359));
    Span4Mux_h I__12910 (
            .O(N__51368),
            .I(N__51354));
    LocalMux I__12909 (
            .O(N__51365),
            .I(N__51354));
    LocalMux I__12908 (
            .O(N__51362),
            .I(N__51351));
    Span12Mux_s4_h I__12907 (
            .O(N__51359),
            .I(N__51346));
    Sp12to4 I__12906 (
            .O(N__51354),
            .I(N__51346));
    Span12Mux_v I__12905 (
            .O(N__51351),
            .I(N__51343));
    Span12Mux_v I__12904 (
            .O(N__51346),
            .I(N__51340));
    Odrv12 I__12903 (
            .O(N__51343),
            .I(ICE_SPI_SCLK));
    Odrv12 I__12902 (
            .O(N__51340),
            .I(ICE_SPI_SCLK));
    InMux I__12901 (
            .O(N__51335),
            .I(N__51332));
    LocalMux I__12900 (
            .O(N__51332),
            .I(N__51329));
    Span4Mux_v I__12899 (
            .O(N__51329),
            .I(N__51326));
    Span4Mux_h I__12898 (
            .O(N__51326),
            .I(N__51323));
    Odrv4 I__12897 (
            .O(N__51323),
            .I(\comm_spi.n10437 ));
    ClkMux I__12896 (
            .O(N__51320),
            .I(N__50675));
    ClkMux I__12895 (
            .O(N__51319),
            .I(N__50675));
    ClkMux I__12894 (
            .O(N__51318),
            .I(N__50675));
    ClkMux I__12893 (
            .O(N__51317),
            .I(N__50675));
    ClkMux I__12892 (
            .O(N__51316),
            .I(N__50675));
    ClkMux I__12891 (
            .O(N__51315),
            .I(N__50675));
    ClkMux I__12890 (
            .O(N__51314),
            .I(N__50675));
    ClkMux I__12889 (
            .O(N__51313),
            .I(N__50675));
    ClkMux I__12888 (
            .O(N__51312),
            .I(N__50675));
    ClkMux I__12887 (
            .O(N__51311),
            .I(N__50675));
    ClkMux I__12886 (
            .O(N__51310),
            .I(N__50675));
    ClkMux I__12885 (
            .O(N__51309),
            .I(N__50675));
    ClkMux I__12884 (
            .O(N__51308),
            .I(N__50675));
    ClkMux I__12883 (
            .O(N__51307),
            .I(N__50675));
    ClkMux I__12882 (
            .O(N__51306),
            .I(N__50675));
    ClkMux I__12881 (
            .O(N__51305),
            .I(N__50675));
    ClkMux I__12880 (
            .O(N__51304),
            .I(N__50675));
    ClkMux I__12879 (
            .O(N__51303),
            .I(N__50675));
    ClkMux I__12878 (
            .O(N__51302),
            .I(N__50675));
    ClkMux I__12877 (
            .O(N__51301),
            .I(N__50675));
    ClkMux I__12876 (
            .O(N__51300),
            .I(N__50675));
    ClkMux I__12875 (
            .O(N__51299),
            .I(N__50675));
    ClkMux I__12874 (
            .O(N__51298),
            .I(N__50675));
    ClkMux I__12873 (
            .O(N__51297),
            .I(N__50675));
    ClkMux I__12872 (
            .O(N__51296),
            .I(N__50675));
    ClkMux I__12871 (
            .O(N__51295),
            .I(N__50675));
    ClkMux I__12870 (
            .O(N__51294),
            .I(N__50675));
    ClkMux I__12869 (
            .O(N__51293),
            .I(N__50675));
    ClkMux I__12868 (
            .O(N__51292),
            .I(N__50675));
    ClkMux I__12867 (
            .O(N__51291),
            .I(N__50675));
    ClkMux I__12866 (
            .O(N__51290),
            .I(N__50675));
    ClkMux I__12865 (
            .O(N__51289),
            .I(N__50675));
    ClkMux I__12864 (
            .O(N__51288),
            .I(N__50675));
    ClkMux I__12863 (
            .O(N__51287),
            .I(N__50675));
    ClkMux I__12862 (
            .O(N__51286),
            .I(N__50675));
    ClkMux I__12861 (
            .O(N__51285),
            .I(N__50675));
    ClkMux I__12860 (
            .O(N__51284),
            .I(N__50675));
    ClkMux I__12859 (
            .O(N__51283),
            .I(N__50675));
    ClkMux I__12858 (
            .O(N__51282),
            .I(N__50675));
    ClkMux I__12857 (
            .O(N__51281),
            .I(N__50675));
    ClkMux I__12856 (
            .O(N__51280),
            .I(N__50675));
    ClkMux I__12855 (
            .O(N__51279),
            .I(N__50675));
    ClkMux I__12854 (
            .O(N__51278),
            .I(N__50675));
    ClkMux I__12853 (
            .O(N__51277),
            .I(N__50675));
    ClkMux I__12852 (
            .O(N__51276),
            .I(N__50675));
    ClkMux I__12851 (
            .O(N__51275),
            .I(N__50675));
    ClkMux I__12850 (
            .O(N__51274),
            .I(N__50675));
    ClkMux I__12849 (
            .O(N__51273),
            .I(N__50675));
    ClkMux I__12848 (
            .O(N__51272),
            .I(N__50675));
    ClkMux I__12847 (
            .O(N__51271),
            .I(N__50675));
    ClkMux I__12846 (
            .O(N__51270),
            .I(N__50675));
    ClkMux I__12845 (
            .O(N__51269),
            .I(N__50675));
    ClkMux I__12844 (
            .O(N__51268),
            .I(N__50675));
    ClkMux I__12843 (
            .O(N__51267),
            .I(N__50675));
    ClkMux I__12842 (
            .O(N__51266),
            .I(N__50675));
    ClkMux I__12841 (
            .O(N__51265),
            .I(N__50675));
    ClkMux I__12840 (
            .O(N__51264),
            .I(N__50675));
    ClkMux I__12839 (
            .O(N__51263),
            .I(N__50675));
    ClkMux I__12838 (
            .O(N__51262),
            .I(N__50675));
    ClkMux I__12837 (
            .O(N__51261),
            .I(N__50675));
    ClkMux I__12836 (
            .O(N__51260),
            .I(N__50675));
    ClkMux I__12835 (
            .O(N__51259),
            .I(N__50675));
    ClkMux I__12834 (
            .O(N__51258),
            .I(N__50675));
    ClkMux I__12833 (
            .O(N__51257),
            .I(N__50675));
    ClkMux I__12832 (
            .O(N__51256),
            .I(N__50675));
    ClkMux I__12831 (
            .O(N__51255),
            .I(N__50675));
    ClkMux I__12830 (
            .O(N__51254),
            .I(N__50675));
    ClkMux I__12829 (
            .O(N__51253),
            .I(N__50675));
    ClkMux I__12828 (
            .O(N__51252),
            .I(N__50675));
    ClkMux I__12827 (
            .O(N__51251),
            .I(N__50675));
    ClkMux I__12826 (
            .O(N__51250),
            .I(N__50675));
    ClkMux I__12825 (
            .O(N__51249),
            .I(N__50675));
    ClkMux I__12824 (
            .O(N__51248),
            .I(N__50675));
    ClkMux I__12823 (
            .O(N__51247),
            .I(N__50675));
    ClkMux I__12822 (
            .O(N__51246),
            .I(N__50675));
    ClkMux I__12821 (
            .O(N__51245),
            .I(N__50675));
    ClkMux I__12820 (
            .O(N__51244),
            .I(N__50675));
    ClkMux I__12819 (
            .O(N__51243),
            .I(N__50675));
    ClkMux I__12818 (
            .O(N__51242),
            .I(N__50675));
    ClkMux I__12817 (
            .O(N__51241),
            .I(N__50675));
    ClkMux I__12816 (
            .O(N__51240),
            .I(N__50675));
    ClkMux I__12815 (
            .O(N__51239),
            .I(N__50675));
    ClkMux I__12814 (
            .O(N__51238),
            .I(N__50675));
    ClkMux I__12813 (
            .O(N__51237),
            .I(N__50675));
    ClkMux I__12812 (
            .O(N__51236),
            .I(N__50675));
    ClkMux I__12811 (
            .O(N__51235),
            .I(N__50675));
    ClkMux I__12810 (
            .O(N__51234),
            .I(N__50675));
    ClkMux I__12809 (
            .O(N__51233),
            .I(N__50675));
    ClkMux I__12808 (
            .O(N__51232),
            .I(N__50675));
    ClkMux I__12807 (
            .O(N__51231),
            .I(N__50675));
    ClkMux I__12806 (
            .O(N__51230),
            .I(N__50675));
    ClkMux I__12805 (
            .O(N__51229),
            .I(N__50675));
    ClkMux I__12804 (
            .O(N__51228),
            .I(N__50675));
    ClkMux I__12803 (
            .O(N__51227),
            .I(N__50675));
    ClkMux I__12802 (
            .O(N__51226),
            .I(N__50675));
    ClkMux I__12801 (
            .O(N__51225),
            .I(N__50675));
    ClkMux I__12800 (
            .O(N__51224),
            .I(N__50675));
    ClkMux I__12799 (
            .O(N__51223),
            .I(N__50675));
    ClkMux I__12798 (
            .O(N__51222),
            .I(N__50675));
    ClkMux I__12797 (
            .O(N__51221),
            .I(N__50675));
    ClkMux I__12796 (
            .O(N__51220),
            .I(N__50675));
    ClkMux I__12795 (
            .O(N__51219),
            .I(N__50675));
    ClkMux I__12794 (
            .O(N__51218),
            .I(N__50675));
    ClkMux I__12793 (
            .O(N__51217),
            .I(N__50675));
    ClkMux I__12792 (
            .O(N__51216),
            .I(N__50675));
    ClkMux I__12791 (
            .O(N__51215),
            .I(N__50675));
    ClkMux I__12790 (
            .O(N__51214),
            .I(N__50675));
    ClkMux I__12789 (
            .O(N__51213),
            .I(N__50675));
    ClkMux I__12788 (
            .O(N__51212),
            .I(N__50675));
    ClkMux I__12787 (
            .O(N__51211),
            .I(N__50675));
    ClkMux I__12786 (
            .O(N__51210),
            .I(N__50675));
    ClkMux I__12785 (
            .O(N__51209),
            .I(N__50675));
    ClkMux I__12784 (
            .O(N__51208),
            .I(N__50675));
    ClkMux I__12783 (
            .O(N__51207),
            .I(N__50675));
    ClkMux I__12782 (
            .O(N__51206),
            .I(N__50675));
    ClkMux I__12781 (
            .O(N__51205),
            .I(N__50675));
    ClkMux I__12780 (
            .O(N__51204),
            .I(N__50675));
    ClkMux I__12779 (
            .O(N__51203),
            .I(N__50675));
    ClkMux I__12778 (
            .O(N__51202),
            .I(N__50675));
    ClkMux I__12777 (
            .O(N__51201),
            .I(N__50675));
    ClkMux I__12776 (
            .O(N__51200),
            .I(N__50675));
    ClkMux I__12775 (
            .O(N__51199),
            .I(N__50675));
    ClkMux I__12774 (
            .O(N__51198),
            .I(N__50675));
    ClkMux I__12773 (
            .O(N__51197),
            .I(N__50675));
    ClkMux I__12772 (
            .O(N__51196),
            .I(N__50675));
    ClkMux I__12771 (
            .O(N__51195),
            .I(N__50675));
    ClkMux I__12770 (
            .O(N__51194),
            .I(N__50675));
    ClkMux I__12769 (
            .O(N__51193),
            .I(N__50675));
    ClkMux I__12768 (
            .O(N__51192),
            .I(N__50675));
    ClkMux I__12767 (
            .O(N__51191),
            .I(N__50675));
    ClkMux I__12766 (
            .O(N__51190),
            .I(N__50675));
    ClkMux I__12765 (
            .O(N__51189),
            .I(N__50675));
    ClkMux I__12764 (
            .O(N__51188),
            .I(N__50675));
    ClkMux I__12763 (
            .O(N__51187),
            .I(N__50675));
    ClkMux I__12762 (
            .O(N__51186),
            .I(N__50675));
    ClkMux I__12761 (
            .O(N__51185),
            .I(N__50675));
    ClkMux I__12760 (
            .O(N__51184),
            .I(N__50675));
    ClkMux I__12759 (
            .O(N__51183),
            .I(N__50675));
    ClkMux I__12758 (
            .O(N__51182),
            .I(N__50675));
    ClkMux I__12757 (
            .O(N__51181),
            .I(N__50675));
    ClkMux I__12756 (
            .O(N__51180),
            .I(N__50675));
    ClkMux I__12755 (
            .O(N__51179),
            .I(N__50675));
    ClkMux I__12754 (
            .O(N__51178),
            .I(N__50675));
    ClkMux I__12753 (
            .O(N__51177),
            .I(N__50675));
    ClkMux I__12752 (
            .O(N__51176),
            .I(N__50675));
    ClkMux I__12751 (
            .O(N__51175),
            .I(N__50675));
    ClkMux I__12750 (
            .O(N__51174),
            .I(N__50675));
    ClkMux I__12749 (
            .O(N__51173),
            .I(N__50675));
    ClkMux I__12748 (
            .O(N__51172),
            .I(N__50675));
    ClkMux I__12747 (
            .O(N__51171),
            .I(N__50675));
    ClkMux I__12746 (
            .O(N__51170),
            .I(N__50675));
    ClkMux I__12745 (
            .O(N__51169),
            .I(N__50675));
    ClkMux I__12744 (
            .O(N__51168),
            .I(N__50675));
    ClkMux I__12743 (
            .O(N__51167),
            .I(N__50675));
    ClkMux I__12742 (
            .O(N__51166),
            .I(N__50675));
    ClkMux I__12741 (
            .O(N__51165),
            .I(N__50675));
    ClkMux I__12740 (
            .O(N__51164),
            .I(N__50675));
    ClkMux I__12739 (
            .O(N__51163),
            .I(N__50675));
    ClkMux I__12738 (
            .O(N__51162),
            .I(N__50675));
    ClkMux I__12737 (
            .O(N__51161),
            .I(N__50675));
    ClkMux I__12736 (
            .O(N__51160),
            .I(N__50675));
    ClkMux I__12735 (
            .O(N__51159),
            .I(N__50675));
    ClkMux I__12734 (
            .O(N__51158),
            .I(N__50675));
    ClkMux I__12733 (
            .O(N__51157),
            .I(N__50675));
    ClkMux I__12732 (
            .O(N__51156),
            .I(N__50675));
    ClkMux I__12731 (
            .O(N__51155),
            .I(N__50675));
    ClkMux I__12730 (
            .O(N__51154),
            .I(N__50675));
    ClkMux I__12729 (
            .O(N__51153),
            .I(N__50675));
    ClkMux I__12728 (
            .O(N__51152),
            .I(N__50675));
    ClkMux I__12727 (
            .O(N__51151),
            .I(N__50675));
    ClkMux I__12726 (
            .O(N__51150),
            .I(N__50675));
    ClkMux I__12725 (
            .O(N__51149),
            .I(N__50675));
    ClkMux I__12724 (
            .O(N__51148),
            .I(N__50675));
    ClkMux I__12723 (
            .O(N__51147),
            .I(N__50675));
    ClkMux I__12722 (
            .O(N__51146),
            .I(N__50675));
    ClkMux I__12721 (
            .O(N__51145),
            .I(N__50675));
    ClkMux I__12720 (
            .O(N__51144),
            .I(N__50675));
    ClkMux I__12719 (
            .O(N__51143),
            .I(N__50675));
    ClkMux I__12718 (
            .O(N__51142),
            .I(N__50675));
    ClkMux I__12717 (
            .O(N__51141),
            .I(N__50675));
    ClkMux I__12716 (
            .O(N__51140),
            .I(N__50675));
    ClkMux I__12715 (
            .O(N__51139),
            .I(N__50675));
    ClkMux I__12714 (
            .O(N__51138),
            .I(N__50675));
    ClkMux I__12713 (
            .O(N__51137),
            .I(N__50675));
    ClkMux I__12712 (
            .O(N__51136),
            .I(N__50675));
    ClkMux I__12711 (
            .O(N__51135),
            .I(N__50675));
    ClkMux I__12710 (
            .O(N__51134),
            .I(N__50675));
    ClkMux I__12709 (
            .O(N__51133),
            .I(N__50675));
    ClkMux I__12708 (
            .O(N__51132),
            .I(N__50675));
    ClkMux I__12707 (
            .O(N__51131),
            .I(N__50675));
    ClkMux I__12706 (
            .O(N__51130),
            .I(N__50675));
    ClkMux I__12705 (
            .O(N__51129),
            .I(N__50675));
    ClkMux I__12704 (
            .O(N__51128),
            .I(N__50675));
    ClkMux I__12703 (
            .O(N__51127),
            .I(N__50675));
    ClkMux I__12702 (
            .O(N__51126),
            .I(N__50675));
    ClkMux I__12701 (
            .O(N__51125),
            .I(N__50675));
    ClkMux I__12700 (
            .O(N__51124),
            .I(N__50675));
    ClkMux I__12699 (
            .O(N__51123),
            .I(N__50675));
    ClkMux I__12698 (
            .O(N__51122),
            .I(N__50675));
    ClkMux I__12697 (
            .O(N__51121),
            .I(N__50675));
    ClkMux I__12696 (
            .O(N__51120),
            .I(N__50675));
    ClkMux I__12695 (
            .O(N__51119),
            .I(N__50675));
    ClkMux I__12694 (
            .O(N__51118),
            .I(N__50675));
    ClkMux I__12693 (
            .O(N__51117),
            .I(N__50675));
    ClkMux I__12692 (
            .O(N__51116),
            .I(N__50675));
    ClkMux I__12691 (
            .O(N__51115),
            .I(N__50675));
    ClkMux I__12690 (
            .O(N__51114),
            .I(N__50675));
    ClkMux I__12689 (
            .O(N__51113),
            .I(N__50675));
    ClkMux I__12688 (
            .O(N__51112),
            .I(N__50675));
    ClkMux I__12687 (
            .O(N__51111),
            .I(N__50675));
    ClkMux I__12686 (
            .O(N__51110),
            .I(N__50675));
    ClkMux I__12685 (
            .O(N__51109),
            .I(N__50675));
    ClkMux I__12684 (
            .O(N__51108),
            .I(N__50675));
    ClkMux I__12683 (
            .O(N__51107),
            .I(N__50675));
    ClkMux I__12682 (
            .O(N__51106),
            .I(N__50675));
    GlobalMux I__12681 (
            .O(N__50675),
            .I(clk_32MHz));
    SRMux I__12680 (
            .O(N__50672),
            .I(N__50669));
    LocalMux I__12679 (
            .O(N__50669),
            .I(N__50666));
    Span4Mux_h I__12678 (
            .O(N__50666),
            .I(N__50663));
    Odrv4 I__12677 (
            .O(N__50663),
            .I(\comm_spi.iclk_N_801 ));
    CEMux I__12676 (
            .O(N__50660),
            .I(N__50657));
    LocalMux I__12675 (
            .O(N__50657),
            .I(N__50653));
    CEMux I__12674 (
            .O(N__50656),
            .I(N__50650));
    Span4Mux_v I__12673 (
            .O(N__50653),
            .I(N__50647));
    LocalMux I__12672 (
            .O(N__50650),
            .I(N__50644));
    Span4Mux_h I__12671 (
            .O(N__50647),
            .I(N__50641));
    Span4Mux_h I__12670 (
            .O(N__50644),
            .I(N__50638));
    Odrv4 I__12669 (
            .O(N__50641),
            .I(n8576));
    Odrv4 I__12668 (
            .O(N__50638),
            .I(n8576));
    CEMux I__12667 (
            .O(N__50633),
            .I(N__50630));
    LocalMux I__12666 (
            .O(N__50630),
            .I(N__50627));
    Span4Mux_h I__12665 (
            .O(N__50627),
            .I(N__50624));
    Odrv4 I__12664 (
            .O(N__50624),
            .I(n8117));
    InMux I__12663 (
            .O(N__50621),
            .I(N__50618));
    LocalMux I__12662 (
            .O(N__50618),
            .I(N__50615));
    Span4Mux_h I__12661 (
            .O(N__50615),
            .I(N__50612));
    Odrv4 I__12660 (
            .O(N__50612),
            .I(n6_adj_1175));
    InMux I__12659 (
            .O(N__50609),
            .I(N__50606));
    LocalMux I__12658 (
            .O(N__50606),
            .I(N__50590));
    InMux I__12657 (
            .O(N__50605),
            .I(N__50583));
    InMux I__12656 (
            .O(N__50604),
            .I(N__50583));
    InMux I__12655 (
            .O(N__50603),
            .I(N__50583));
    InMux I__12654 (
            .O(N__50602),
            .I(N__50575));
    InMux I__12653 (
            .O(N__50601),
            .I(N__50575));
    InMux I__12652 (
            .O(N__50600),
            .I(N__50570));
    InMux I__12651 (
            .O(N__50599),
            .I(N__50570));
    InMux I__12650 (
            .O(N__50598),
            .I(N__50565));
    InMux I__12649 (
            .O(N__50597),
            .I(N__50565));
    InMux I__12648 (
            .O(N__50596),
            .I(N__50562));
    InMux I__12647 (
            .O(N__50595),
            .I(N__50555));
    InMux I__12646 (
            .O(N__50594),
            .I(N__50547));
    InMux I__12645 (
            .O(N__50593),
            .I(N__50544));
    Span4Mux_v I__12644 (
            .O(N__50590),
            .I(N__50541));
    LocalMux I__12643 (
            .O(N__50583),
            .I(N__50538));
    InMux I__12642 (
            .O(N__50582),
            .I(N__50533));
    InMux I__12641 (
            .O(N__50581),
            .I(N__50528));
    InMux I__12640 (
            .O(N__50580),
            .I(N__50528));
    LocalMux I__12639 (
            .O(N__50575),
            .I(N__50525));
    LocalMux I__12638 (
            .O(N__50570),
            .I(N__50520));
    LocalMux I__12637 (
            .O(N__50565),
            .I(N__50520));
    LocalMux I__12636 (
            .O(N__50562),
            .I(N__50517));
    InMux I__12635 (
            .O(N__50561),
            .I(N__50514));
    InMux I__12634 (
            .O(N__50560),
            .I(N__50493));
    InMux I__12633 (
            .O(N__50559),
            .I(N__50493));
    InMux I__12632 (
            .O(N__50558),
            .I(N__50490));
    LocalMux I__12631 (
            .O(N__50555),
            .I(N__50487));
    InMux I__12630 (
            .O(N__50554),
            .I(N__50478));
    InMux I__12629 (
            .O(N__50553),
            .I(N__50478));
    InMux I__12628 (
            .O(N__50552),
            .I(N__50478));
    InMux I__12627 (
            .O(N__50551),
            .I(N__50478));
    CascadeMux I__12626 (
            .O(N__50550),
            .I(N__50473));
    LocalMux I__12625 (
            .O(N__50547),
            .I(N__50468));
    LocalMux I__12624 (
            .O(N__50544),
            .I(N__50468));
    Span4Mux_h I__12623 (
            .O(N__50541),
            .I(N__50465));
    Span12Mux_v I__12622 (
            .O(N__50538),
            .I(N__50462));
    InMux I__12621 (
            .O(N__50537),
            .I(N__50459));
    InMux I__12620 (
            .O(N__50536),
            .I(N__50456));
    LocalMux I__12619 (
            .O(N__50533),
            .I(N__50447));
    LocalMux I__12618 (
            .O(N__50528),
            .I(N__50447));
    Span4Mux_v I__12617 (
            .O(N__50525),
            .I(N__50447));
    Span4Mux_v I__12616 (
            .O(N__50520),
            .I(N__50447));
    Span4Mux_h I__12615 (
            .O(N__50517),
            .I(N__50442));
    LocalMux I__12614 (
            .O(N__50514),
            .I(N__50442));
    InMux I__12613 (
            .O(N__50513),
            .I(N__50439));
    InMux I__12612 (
            .O(N__50512),
            .I(N__50428));
    InMux I__12611 (
            .O(N__50511),
            .I(N__50428));
    InMux I__12610 (
            .O(N__50510),
            .I(N__50428));
    InMux I__12609 (
            .O(N__50509),
            .I(N__50428));
    InMux I__12608 (
            .O(N__50508),
            .I(N__50428));
    InMux I__12607 (
            .O(N__50507),
            .I(N__50421));
    InMux I__12606 (
            .O(N__50506),
            .I(N__50421));
    InMux I__12605 (
            .O(N__50505),
            .I(N__50421));
    InMux I__12604 (
            .O(N__50504),
            .I(N__50416));
    InMux I__12603 (
            .O(N__50503),
            .I(N__50416));
    InMux I__12602 (
            .O(N__50502),
            .I(N__50413));
    InMux I__12601 (
            .O(N__50501),
            .I(N__50408));
    InMux I__12600 (
            .O(N__50500),
            .I(N__50408));
    InMux I__12599 (
            .O(N__50499),
            .I(N__50403));
    InMux I__12598 (
            .O(N__50498),
            .I(N__50403));
    LocalMux I__12597 (
            .O(N__50493),
            .I(N__50394));
    LocalMux I__12596 (
            .O(N__50490),
            .I(N__50394));
    Span4Mux_v I__12595 (
            .O(N__50487),
            .I(N__50394));
    LocalMux I__12594 (
            .O(N__50478),
            .I(N__50394));
    InMux I__12593 (
            .O(N__50477),
            .I(N__50387));
    InMux I__12592 (
            .O(N__50476),
            .I(N__50387));
    InMux I__12591 (
            .O(N__50473),
            .I(N__50387));
    Span4Mux_v I__12590 (
            .O(N__50468),
            .I(N__50384));
    Sp12to4 I__12589 (
            .O(N__50465),
            .I(N__50377));
    Span12Mux_h I__12588 (
            .O(N__50462),
            .I(N__50377));
    LocalMux I__12587 (
            .O(N__50459),
            .I(N__50377));
    LocalMux I__12586 (
            .O(N__50456),
            .I(N__50370));
    Span4Mux_h I__12585 (
            .O(N__50447),
            .I(N__50370));
    Span4Mux_v I__12584 (
            .O(N__50442),
            .I(N__50370));
    LocalMux I__12583 (
            .O(N__50439),
            .I(comm_state_0));
    LocalMux I__12582 (
            .O(N__50428),
            .I(comm_state_0));
    LocalMux I__12581 (
            .O(N__50421),
            .I(comm_state_0));
    LocalMux I__12580 (
            .O(N__50416),
            .I(comm_state_0));
    LocalMux I__12579 (
            .O(N__50413),
            .I(comm_state_0));
    LocalMux I__12578 (
            .O(N__50408),
            .I(comm_state_0));
    LocalMux I__12577 (
            .O(N__50403),
            .I(comm_state_0));
    Odrv4 I__12576 (
            .O(N__50394),
            .I(comm_state_0));
    LocalMux I__12575 (
            .O(N__50387),
            .I(comm_state_0));
    Odrv4 I__12574 (
            .O(N__50384),
            .I(comm_state_0));
    Odrv12 I__12573 (
            .O(N__50377),
            .I(comm_state_0));
    Odrv4 I__12572 (
            .O(N__50370),
            .I(comm_state_0));
    InMux I__12571 (
            .O(N__50345),
            .I(N__50334));
    InMux I__12570 (
            .O(N__50344),
            .I(N__50331));
    InMux I__12569 (
            .O(N__50343),
            .I(N__50297));
    InMux I__12568 (
            .O(N__50342),
            .I(N__50294));
    InMux I__12567 (
            .O(N__50341),
            .I(N__50247));
    InMux I__12566 (
            .O(N__50340),
            .I(N__50247));
    InMux I__12565 (
            .O(N__50339),
            .I(N__50240));
    InMux I__12564 (
            .O(N__50338),
            .I(N__50240));
    InMux I__12563 (
            .O(N__50337),
            .I(N__50240));
    LocalMux I__12562 (
            .O(N__50334),
            .I(N__50235));
    LocalMux I__12561 (
            .O(N__50331),
            .I(N__50235));
    InMux I__12560 (
            .O(N__50330),
            .I(N__50230));
    InMux I__12559 (
            .O(N__50329),
            .I(N__50230));
    InMux I__12558 (
            .O(N__50328),
            .I(N__50221));
    InMux I__12557 (
            .O(N__50327),
            .I(N__50221));
    InMux I__12556 (
            .O(N__50326),
            .I(N__50221));
    InMux I__12555 (
            .O(N__50325),
            .I(N__50221));
    CascadeMux I__12554 (
            .O(N__50324),
            .I(N__50216));
    InMux I__12553 (
            .O(N__50323),
            .I(N__50212));
    CascadeMux I__12552 (
            .O(N__50322),
            .I(N__50207));
    InMux I__12551 (
            .O(N__50321),
            .I(N__50204));
    InMux I__12550 (
            .O(N__50320),
            .I(N__50183));
    InMux I__12549 (
            .O(N__50319),
            .I(N__50183));
    InMux I__12548 (
            .O(N__50318),
            .I(N__50183));
    InMux I__12547 (
            .O(N__50317),
            .I(N__50183));
    InMux I__12546 (
            .O(N__50316),
            .I(N__50183));
    InMux I__12545 (
            .O(N__50315),
            .I(N__50183));
    InMux I__12544 (
            .O(N__50314),
            .I(N__50183));
    InMux I__12543 (
            .O(N__50313),
            .I(N__50183));
    InMux I__12542 (
            .O(N__50312),
            .I(N__50178));
    InMux I__12541 (
            .O(N__50311),
            .I(N__50178));
    InMux I__12540 (
            .O(N__50310),
            .I(N__50167));
    InMux I__12539 (
            .O(N__50309),
            .I(N__50167));
    InMux I__12538 (
            .O(N__50308),
            .I(N__50167));
    InMux I__12537 (
            .O(N__50307),
            .I(N__50167));
    InMux I__12536 (
            .O(N__50306),
            .I(N__50167));
    InMux I__12535 (
            .O(N__50305),
            .I(N__50164));
    InMux I__12534 (
            .O(N__50304),
            .I(N__50153));
    InMux I__12533 (
            .O(N__50303),
            .I(N__50153));
    InMux I__12532 (
            .O(N__50302),
            .I(N__50153));
    InMux I__12531 (
            .O(N__50301),
            .I(N__50153));
    InMux I__12530 (
            .O(N__50300),
            .I(N__50153));
    LocalMux I__12529 (
            .O(N__50297),
            .I(N__50144));
    LocalMux I__12528 (
            .O(N__50294),
            .I(N__50144));
    CascadeMux I__12527 (
            .O(N__50293),
            .I(N__50138));
    CascadeMux I__12526 (
            .O(N__50292),
            .I(N__50135));
    InMux I__12525 (
            .O(N__50291),
            .I(N__50132));
    CascadeMux I__12524 (
            .O(N__50290),
            .I(N__50128));
    InMux I__12523 (
            .O(N__50289),
            .I(N__50124));
    InMux I__12522 (
            .O(N__50288),
            .I(N__50115));
    InMux I__12521 (
            .O(N__50287),
            .I(N__50115));
    InMux I__12520 (
            .O(N__50286),
            .I(N__50099));
    InMux I__12519 (
            .O(N__50285),
            .I(N__50099));
    InMux I__12518 (
            .O(N__50284),
            .I(N__50099));
    InMux I__12517 (
            .O(N__50283),
            .I(N__50094));
    InMux I__12516 (
            .O(N__50282),
            .I(N__50094));
    InMux I__12515 (
            .O(N__50281),
            .I(N__50085));
    InMux I__12514 (
            .O(N__50280),
            .I(N__50078));
    InMux I__12513 (
            .O(N__50279),
            .I(N__50078));
    InMux I__12512 (
            .O(N__50278),
            .I(N__50078));
    InMux I__12511 (
            .O(N__50277),
            .I(N__50069));
    InMux I__12510 (
            .O(N__50276),
            .I(N__50069));
    InMux I__12509 (
            .O(N__50275),
            .I(N__50069));
    InMux I__12508 (
            .O(N__50274),
            .I(N__50069));
    InMux I__12507 (
            .O(N__50273),
            .I(N__50060));
    InMux I__12506 (
            .O(N__50272),
            .I(N__50060));
    InMux I__12505 (
            .O(N__50271),
            .I(N__50060));
    InMux I__12504 (
            .O(N__50270),
            .I(N__50060));
    InMux I__12503 (
            .O(N__50269),
            .I(N__50057));
    InMux I__12502 (
            .O(N__50268),
            .I(N__50054));
    InMux I__12501 (
            .O(N__50267),
            .I(N__50051));
    InMux I__12500 (
            .O(N__50266),
            .I(N__50048));
    InMux I__12499 (
            .O(N__50265),
            .I(N__50031));
    InMux I__12498 (
            .O(N__50264),
            .I(N__50031));
    InMux I__12497 (
            .O(N__50263),
            .I(N__50031));
    InMux I__12496 (
            .O(N__50262),
            .I(N__50031));
    InMux I__12495 (
            .O(N__50261),
            .I(N__50031));
    InMux I__12494 (
            .O(N__50260),
            .I(N__50031));
    InMux I__12493 (
            .O(N__50259),
            .I(N__50031));
    InMux I__12492 (
            .O(N__50258),
            .I(N__50031));
    InMux I__12491 (
            .O(N__50257),
            .I(N__50018));
    InMux I__12490 (
            .O(N__50256),
            .I(N__50018));
    InMux I__12489 (
            .O(N__50255),
            .I(N__50018));
    InMux I__12488 (
            .O(N__50254),
            .I(N__50018));
    InMux I__12487 (
            .O(N__50253),
            .I(N__50018));
    InMux I__12486 (
            .O(N__50252),
            .I(N__50018));
    LocalMux I__12485 (
            .O(N__50247),
            .I(N__50015));
    LocalMux I__12484 (
            .O(N__50240),
            .I(N__50012));
    Span4Mux_h I__12483 (
            .O(N__50235),
            .I(N__50005));
    LocalMux I__12482 (
            .O(N__50230),
            .I(N__50005));
    LocalMux I__12481 (
            .O(N__50221),
            .I(N__50005));
    CascadeMux I__12480 (
            .O(N__50220),
            .I(N__50001));
    CascadeMux I__12479 (
            .O(N__50219),
            .I(N__49997));
    InMux I__12478 (
            .O(N__50216),
            .I(N__49993));
    InMux I__12477 (
            .O(N__50215),
            .I(N__49990));
    LocalMux I__12476 (
            .O(N__50212),
            .I(N__49987));
    InMux I__12475 (
            .O(N__50211),
            .I(N__49980));
    InMux I__12474 (
            .O(N__50210),
            .I(N__49980));
    InMux I__12473 (
            .O(N__50207),
            .I(N__49980));
    LocalMux I__12472 (
            .O(N__50204),
            .I(N__49977));
    InMux I__12471 (
            .O(N__50203),
            .I(N__49972));
    InMux I__12470 (
            .O(N__50202),
            .I(N__49972));
    InMux I__12469 (
            .O(N__50201),
            .I(N__49967));
    InMux I__12468 (
            .O(N__50200),
            .I(N__49967));
    LocalMux I__12467 (
            .O(N__50183),
            .I(N__49962));
    LocalMux I__12466 (
            .O(N__50178),
            .I(N__49957));
    LocalMux I__12465 (
            .O(N__50167),
            .I(N__49957));
    LocalMux I__12464 (
            .O(N__50164),
            .I(N__49952));
    LocalMux I__12463 (
            .O(N__50153),
            .I(N__49952));
    InMux I__12462 (
            .O(N__50152),
            .I(N__49943));
    InMux I__12461 (
            .O(N__50151),
            .I(N__49943));
    InMux I__12460 (
            .O(N__50150),
            .I(N__49943));
    InMux I__12459 (
            .O(N__50149),
            .I(N__49943));
    Span4Mux_h I__12458 (
            .O(N__50144),
            .I(N__49940));
    CascadeMux I__12457 (
            .O(N__50143),
            .I(N__49935));
    InMux I__12456 (
            .O(N__50142),
            .I(N__49932));
    InMux I__12455 (
            .O(N__50141),
            .I(N__49929));
    InMux I__12454 (
            .O(N__50138),
            .I(N__49924));
    InMux I__12453 (
            .O(N__50135),
            .I(N__49924));
    LocalMux I__12452 (
            .O(N__50132),
            .I(N__49921));
    InMux I__12451 (
            .O(N__50131),
            .I(N__49914));
    InMux I__12450 (
            .O(N__50128),
            .I(N__49914));
    InMux I__12449 (
            .O(N__50127),
            .I(N__49914));
    LocalMux I__12448 (
            .O(N__50124),
            .I(N__49911));
    InMux I__12447 (
            .O(N__50123),
            .I(N__49902));
    InMux I__12446 (
            .O(N__50122),
            .I(N__49902));
    InMux I__12445 (
            .O(N__50121),
            .I(N__49902));
    InMux I__12444 (
            .O(N__50120),
            .I(N__49902));
    LocalMux I__12443 (
            .O(N__50115),
            .I(N__49899));
    InMux I__12442 (
            .O(N__50114),
            .I(N__49882));
    InMux I__12441 (
            .O(N__50113),
            .I(N__49882));
    InMux I__12440 (
            .O(N__50112),
            .I(N__49882));
    CascadeMux I__12439 (
            .O(N__50111),
            .I(N__49876));
    InMux I__12438 (
            .O(N__50110),
            .I(N__49871));
    InMux I__12437 (
            .O(N__50109),
            .I(N__49865));
    InMux I__12436 (
            .O(N__50108),
            .I(N__49862));
    InMux I__12435 (
            .O(N__50107),
            .I(N__49859));
    InMux I__12434 (
            .O(N__50106),
            .I(N__49856));
    LocalMux I__12433 (
            .O(N__50099),
            .I(N__49851));
    LocalMux I__12432 (
            .O(N__50094),
            .I(N__49851));
    InMux I__12431 (
            .O(N__50093),
            .I(N__49848));
    InMux I__12430 (
            .O(N__50092),
            .I(N__49845));
    InMux I__12429 (
            .O(N__50091),
            .I(N__49836));
    InMux I__12428 (
            .O(N__50090),
            .I(N__49836));
    InMux I__12427 (
            .O(N__50089),
            .I(N__49836));
    InMux I__12426 (
            .O(N__50088),
            .I(N__49836));
    LocalMux I__12425 (
            .O(N__50085),
            .I(N__49831));
    LocalMux I__12424 (
            .O(N__50078),
            .I(N__49831));
    LocalMux I__12423 (
            .O(N__50069),
            .I(N__49820));
    LocalMux I__12422 (
            .O(N__50060),
            .I(N__49820));
    LocalMux I__12421 (
            .O(N__50057),
            .I(N__49820));
    LocalMux I__12420 (
            .O(N__50054),
            .I(N__49820));
    LocalMux I__12419 (
            .O(N__50051),
            .I(N__49820));
    LocalMux I__12418 (
            .O(N__50048),
            .I(N__49806));
    LocalMux I__12417 (
            .O(N__50031),
            .I(N__49806));
    LocalMux I__12416 (
            .O(N__50018),
            .I(N__49806));
    Span4Mux_h I__12415 (
            .O(N__50015),
            .I(N__49806));
    Span4Mux_h I__12414 (
            .O(N__50012),
            .I(N__49806));
    Span4Mux_v I__12413 (
            .O(N__50005),
            .I(N__49806));
    InMux I__12412 (
            .O(N__50004),
            .I(N__49795));
    InMux I__12411 (
            .O(N__50001),
            .I(N__49795));
    InMux I__12410 (
            .O(N__50000),
            .I(N__49795));
    InMux I__12409 (
            .O(N__49997),
            .I(N__49795));
    InMux I__12408 (
            .O(N__49996),
            .I(N__49795));
    LocalMux I__12407 (
            .O(N__49993),
            .I(N__49792));
    LocalMux I__12406 (
            .O(N__49990),
            .I(N__49779));
    Span4Mux_h I__12405 (
            .O(N__49987),
            .I(N__49779));
    LocalMux I__12404 (
            .O(N__49980),
            .I(N__49779));
    Span4Mux_h I__12403 (
            .O(N__49977),
            .I(N__49779));
    LocalMux I__12402 (
            .O(N__49972),
            .I(N__49779));
    LocalMux I__12401 (
            .O(N__49967),
            .I(N__49779));
    InMux I__12400 (
            .O(N__49966),
            .I(N__49776));
    InMux I__12399 (
            .O(N__49965),
            .I(N__49770));
    Span4Mux_v I__12398 (
            .O(N__49962),
            .I(N__49763));
    Span4Mux_v I__12397 (
            .O(N__49957),
            .I(N__49763));
    Span4Mux_v I__12396 (
            .O(N__49952),
            .I(N__49763));
    LocalMux I__12395 (
            .O(N__49943),
            .I(N__49758));
    Span4Mux_h I__12394 (
            .O(N__49940),
            .I(N__49758));
    InMux I__12393 (
            .O(N__49939),
            .I(N__49753));
    InMux I__12392 (
            .O(N__49938),
            .I(N__49753));
    InMux I__12391 (
            .O(N__49935),
            .I(N__49750));
    LocalMux I__12390 (
            .O(N__49932),
            .I(N__49747));
    LocalMux I__12389 (
            .O(N__49929),
            .I(N__49742));
    LocalMux I__12388 (
            .O(N__49924),
            .I(N__49742));
    Span4Mux_h I__12387 (
            .O(N__49921),
            .I(N__49736));
    LocalMux I__12386 (
            .O(N__49914),
            .I(N__49736));
    Span4Mux_v I__12385 (
            .O(N__49911),
            .I(N__49726));
    LocalMux I__12384 (
            .O(N__49902),
            .I(N__49726));
    Span4Mux_h I__12383 (
            .O(N__49899),
            .I(N__49726));
    InMux I__12382 (
            .O(N__49898),
            .I(N__49721));
    InMux I__12381 (
            .O(N__49897),
            .I(N__49721));
    InMux I__12380 (
            .O(N__49896),
            .I(N__49716));
    InMux I__12379 (
            .O(N__49895),
            .I(N__49716));
    InMux I__12378 (
            .O(N__49894),
            .I(N__49703));
    InMux I__12377 (
            .O(N__49893),
            .I(N__49703));
    InMux I__12376 (
            .O(N__49892),
            .I(N__49703));
    InMux I__12375 (
            .O(N__49891),
            .I(N__49703));
    InMux I__12374 (
            .O(N__49890),
            .I(N__49703));
    InMux I__12373 (
            .O(N__49889),
            .I(N__49703));
    LocalMux I__12372 (
            .O(N__49882),
            .I(N__49700));
    InMux I__12371 (
            .O(N__49881),
            .I(N__49695));
    InMux I__12370 (
            .O(N__49880),
            .I(N__49695));
    InMux I__12369 (
            .O(N__49879),
            .I(N__49688));
    InMux I__12368 (
            .O(N__49876),
            .I(N__49688));
    InMux I__12367 (
            .O(N__49875),
            .I(N__49688));
    InMux I__12366 (
            .O(N__49874),
            .I(N__49685));
    LocalMux I__12365 (
            .O(N__49871),
            .I(N__49682));
    InMux I__12364 (
            .O(N__49870),
            .I(N__49675));
    InMux I__12363 (
            .O(N__49869),
            .I(N__49675));
    InMux I__12362 (
            .O(N__49868),
            .I(N__49675));
    LocalMux I__12361 (
            .O(N__49865),
            .I(N__49660));
    LocalMux I__12360 (
            .O(N__49862),
            .I(N__49660));
    LocalMux I__12359 (
            .O(N__49859),
            .I(N__49660));
    LocalMux I__12358 (
            .O(N__49856),
            .I(N__49660));
    Sp12to4 I__12357 (
            .O(N__49851),
            .I(N__49660));
    LocalMux I__12356 (
            .O(N__49848),
            .I(N__49660));
    LocalMux I__12355 (
            .O(N__49845),
            .I(N__49660));
    LocalMux I__12354 (
            .O(N__49836),
            .I(N__49653));
    Span4Mux_v I__12353 (
            .O(N__49831),
            .I(N__49653));
    Span4Mux_v I__12352 (
            .O(N__49820),
            .I(N__49653));
    InMux I__12351 (
            .O(N__49819),
            .I(N__49650));
    Span4Mux_h I__12350 (
            .O(N__49806),
            .I(N__49645));
    LocalMux I__12349 (
            .O(N__49795),
            .I(N__49645));
    Span4Mux_h I__12348 (
            .O(N__49792),
            .I(N__49638));
    Span4Mux_v I__12347 (
            .O(N__49779),
            .I(N__49638));
    LocalMux I__12346 (
            .O(N__49776),
            .I(N__49638));
    InMux I__12345 (
            .O(N__49775),
            .I(N__49631));
    InMux I__12344 (
            .O(N__49774),
            .I(N__49631));
    InMux I__12343 (
            .O(N__49773),
            .I(N__49631));
    LocalMux I__12342 (
            .O(N__49770),
            .I(N__49628));
    Span4Mux_h I__12341 (
            .O(N__49763),
            .I(N__49615));
    Span4Mux_v I__12340 (
            .O(N__49758),
            .I(N__49615));
    LocalMux I__12339 (
            .O(N__49753),
            .I(N__49615));
    LocalMux I__12338 (
            .O(N__49750),
            .I(N__49615));
    Span4Mux_v I__12337 (
            .O(N__49747),
            .I(N__49615));
    Span4Mux_h I__12336 (
            .O(N__49742),
            .I(N__49615));
    InMux I__12335 (
            .O(N__49741),
            .I(N__49612));
    Span4Mux_h I__12334 (
            .O(N__49736),
            .I(N__49609));
    InMux I__12333 (
            .O(N__49735),
            .I(N__49602));
    InMux I__12332 (
            .O(N__49734),
            .I(N__49602));
    InMux I__12331 (
            .O(N__49733),
            .I(N__49602));
    Span4Mux_v I__12330 (
            .O(N__49726),
            .I(N__49599));
    LocalMux I__12329 (
            .O(N__49721),
            .I(N__49576));
    LocalMux I__12328 (
            .O(N__49716),
            .I(N__49576));
    LocalMux I__12327 (
            .O(N__49703),
            .I(N__49576));
    Span12Mux_v I__12326 (
            .O(N__49700),
            .I(N__49576));
    LocalMux I__12325 (
            .O(N__49695),
            .I(N__49576));
    LocalMux I__12324 (
            .O(N__49688),
            .I(N__49576));
    LocalMux I__12323 (
            .O(N__49685),
            .I(N__49576));
    Span12Mux_v I__12322 (
            .O(N__49682),
            .I(N__49576));
    LocalMux I__12321 (
            .O(N__49675),
            .I(N__49576));
    Span12Mux_v I__12320 (
            .O(N__49660),
            .I(N__49576));
    Sp12to4 I__12319 (
            .O(N__49653),
            .I(N__49576));
    LocalMux I__12318 (
            .O(N__49650),
            .I(N__49569));
    Span4Mux_h I__12317 (
            .O(N__49645),
            .I(N__49569));
    Span4Mux_h I__12316 (
            .O(N__49638),
            .I(N__49569));
    LocalMux I__12315 (
            .O(N__49631),
            .I(comm_state_1));
    Odrv4 I__12314 (
            .O(N__49628),
            .I(comm_state_1));
    Odrv4 I__12313 (
            .O(N__49615),
            .I(comm_state_1));
    LocalMux I__12312 (
            .O(N__49612),
            .I(comm_state_1));
    Odrv4 I__12311 (
            .O(N__49609),
            .I(comm_state_1));
    LocalMux I__12310 (
            .O(N__49602),
            .I(comm_state_1));
    Odrv4 I__12309 (
            .O(N__49599),
            .I(comm_state_1));
    Odrv12 I__12308 (
            .O(N__49576),
            .I(comm_state_1));
    Odrv4 I__12307 (
            .O(N__49569),
            .I(comm_state_1));
    InMux I__12306 (
            .O(N__49550),
            .I(N__49532));
    InMux I__12305 (
            .O(N__49549),
            .I(N__49528));
    InMux I__12304 (
            .O(N__49548),
            .I(N__49521));
    InMux I__12303 (
            .O(N__49547),
            .I(N__49521));
    InMux I__12302 (
            .O(N__49546),
            .I(N__49521));
    InMux I__12301 (
            .O(N__49545),
            .I(N__49514));
    InMux I__12300 (
            .O(N__49544),
            .I(N__49514));
    InMux I__12299 (
            .O(N__49543),
            .I(N__49514));
    InMux I__12298 (
            .O(N__49542),
            .I(N__49509));
    InMux I__12297 (
            .O(N__49541),
            .I(N__49509));
    InMux I__12296 (
            .O(N__49540),
            .I(N__49499));
    InMux I__12295 (
            .O(N__49539),
            .I(N__49499));
    CascadeMux I__12294 (
            .O(N__49538),
            .I(N__49496));
    InMux I__12293 (
            .O(N__49537),
            .I(N__49493));
    InMux I__12292 (
            .O(N__49536),
            .I(N__49488));
    InMux I__12291 (
            .O(N__49535),
            .I(N__49488));
    LocalMux I__12290 (
            .O(N__49532),
            .I(N__49485));
    InMux I__12289 (
            .O(N__49531),
            .I(N__49482));
    LocalMux I__12288 (
            .O(N__49528),
            .I(N__49474));
    LocalMux I__12287 (
            .O(N__49521),
            .I(N__49474));
    LocalMux I__12286 (
            .O(N__49514),
            .I(N__49464));
    LocalMux I__12285 (
            .O(N__49509),
            .I(N__49464));
    InMux I__12284 (
            .O(N__49508),
            .I(N__49453));
    InMux I__12283 (
            .O(N__49507),
            .I(N__49453));
    InMux I__12282 (
            .O(N__49506),
            .I(N__49453));
    InMux I__12281 (
            .O(N__49505),
            .I(N__49453));
    InMux I__12280 (
            .O(N__49504),
            .I(N__49453));
    LocalMux I__12279 (
            .O(N__49499),
            .I(N__49450));
    InMux I__12278 (
            .O(N__49496),
            .I(N__49447));
    LocalMux I__12277 (
            .O(N__49493),
            .I(N__49442));
    LocalMux I__12276 (
            .O(N__49488),
            .I(N__49439));
    Span4Mux_v I__12275 (
            .O(N__49485),
            .I(N__49427));
    LocalMux I__12274 (
            .O(N__49482),
            .I(N__49427));
    InMux I__12273 (
            .O(N__49481),
            .I(N__49422));
    InMux I__12272 (
            .O(N__49480),
            .I(N__49422));
    InMux I__12271 (
            .O(N__49479),
            .I(N__49419));
    Span4Mux_v I__12270 (
            .O(N__49474),
            .I(N__49416));
    InMux I__12269 (
            .O(N__49473),
            .I(N__49407));
    InMux I__12268 (
            .O(N__49472),
            .I(N__49407));
    InMux I__12267 (
            .O(N__49471),
            .I(N__49407));
    InMux I__12266 (
            .O(N__49470),
            .I(N__49407));
    InMux I__12265 (
            .O(N__49469),
            .I(N__49399));
    Span4Mux_v I__12264 (
            .O(N__49464),
            .I(N__49394));
    LocalMux I__12263 (
            .O(N__49453),
            .I(N__49394));
    Span4Mux_v I__12262 (
            .O(N__49450),
            .I(N__49389));
    LocalMux I__12261 (
            .O(N__49447),
            .I(N__49389));
    InMux I__12260 (
            .O(N__49446),
            .I(N__49386));
    InMux I__12259 (
            .O(N__49445),
            .I(N__49383));
    Span12Mux_v I__12258 (
            .O(N__49442),
            .I(N__49378));
    Span12Mux_s10_h I__12257 (
            .O(N__49439),
            .I(N__49378));
    InMux I__12256 (
            .O(N__49438),
            .I(N__49375));
    InMux I__12255 (
            .O(N__49437),
            .I(N__49372));
    InMux I__12254 (
            .O(N__49436),
            .I(N__49369));
    InMux I__12253 (
            .O(N__49435),
            .I(N__49360));
    InMux I__12252 (
            .O(N__49434),
            .I(N__49360));
    InMux I__12251 (
            .O(N__49433),
            .I(N__49360));
    InMux I__12250 (
            .O(N__49432),
            .I(N__49360));
    Span4Mux_h I__12249 (
            .O(N__49427),
            .I(N__49357));
    LocalMux I__12248 (
            .O(N__49422),
            .I(N__49348));
    LocalMux I__12247 (
            .O(N__49419),
            .I(N__49348));
    Sp12to4 I__12246 (
            .O(N__49416),
            .I(N__49348));
    LocalMux I__12245 (
            .O(N__49407),
            .I(N__49348));
    InMux I__12244 (
            .O(N__49406),
            .I(N__49343));
    InMux I__12243 (
            .O(N__49405),
            .I(N__49343));
    InMux I__12242 (
            .O(N__49404),
            .I(N__49338));
    InMux I__12241 (
            .O(N__49403),
            .I(N__49338));
    InMux I__12240 (
            .O(N__49402),
            .I(N__49335));
    LocalMux I__12239 (
            .O(N__49399),
            .I(N__49328));
    Span4Mux_h I__12238 (
            .O(N__49394),
            .I(N__49328));
    Span4Mux_h I__12237 (
            .O(N__49389),
            .I(N__49328));
    LocalMux I__12236 (
            .O(N__49386),
            .I(N__49321));
    LocalMux I__12235 (
            .O(N__49383),
            .I(N__49321));
    Span12Mux_h I__12234 (
            .O(N__49378),
            .I(N__49321));
    LocalMux I__12233 (
            .O(N__49375),
            .I(comm_state_2));
    LocalMux I__12232 (
            .O(N__49372),
            .I(comm_state_2));
    LocalMux I__12231 (
            .O(N__49369),
            .I(comm_state_2));
    LocalMux I__12230 (
            .O(N__49360),
            .I(comm_state_2));
    Odrv4 I__12229 (
            .O(N__49357),
            .I(comm_state_2));
    Odrv12 I__12228 (
            .O(N__49348),
            .I(comm_state_2));
    LocalMux I__12227 (
            .O(N__49343),
            .I(comm_state_2));
    LocalMux I__12226 (
            .O(N__49338),
            .I(comm_state_2));
    LocalMux I__12225 (
            .O(N__49335),
            .I(comm_state_2));
    Odrv4 I__12224 (
            .O(N__49328),
            .I(comm_state_2));
    Odrv12 I__12223 (
            .O(N__49321),
            .I(comm_state_2));
    CEMux I__12222 (
            .O(N__49298),
            .I(N__49295));
    LocalMux I__12221 (
            .O(N__49295),
            .I(N__49292));
    Span4Mux_v I__12220 (
            .O(N__49292),
            .I(N__49289));
    Odrv4 I__12219 (
            .O(N__49289),
            .I(n8129));
    CascadeMux I__12218 (
            .O(N__49286),
            .I(N__49282));
    InMux I__12217 (
            .O(N__49285),
            .I(N__49278));
    InMux I__12216 (
            .O(N__49282),
            .I(N__49273));
    InMux I__12215 (
            .O(N__49281),
            .I(N__49273));
    LocalMux I__12214 (
            .O(N__49278),
            .I(cmd_rdadctmp_19_adj_1093));
    LocalMux I__12213 (
            .O(N__49273),
            .I(cmd_rdadctmp_19_adj_1093));
    InMux I__12212 (
            .O(N__49268),
            .I(N__49257));
    InMux I__12211 (
            .O(N__49267),
            .I(N__49257));
    CascadeMux I__12210 (
            .O(N__49266),
            .I(N__49253));
    InMux I__12209 (
            .O(N__49265),
            .I(N__49244));
    InMux I__12208 (
            .O(N__49264),
            .I(N__49244));
    InMux I__12207 (
            .O(N__49263),
            .I(N__49244));
    InMux I__12206 (
            .O(N__49262),
            .I(N__49244));
    LocalMux I__12205 (
            .O(N__49257),
            .I(N__49234));
    CascadeMux I__12204 (
            .O(N__49256),
            .I(N__49228));
    InMux I__12203 (
            .O(N__49253),
            .I(N__49222));
    LocalMux I__12202 (
            .O(N__49244),
            .I(N__49217));
    InMux I__12201 (
            .O(N__49243),
            .I(N__49214));
    InMux I__12200 (
            .O(N__49242),
            .I(N__49209));
    CascadeMux I__12199 (
            .O(N__49241),
            .I(N__49206));
    InMux I__12198 (
            .O(N__49240),
            .I(N__49186));
    InMux I__12197 (
            .O(N__49239),
            .I(N__49183));
    InMux I__12196 (
            .O(N__49238),
            .I(N__49178));
    InMux I__12195 (
            .O(N__49237),
            .I(N__49178));
    Span4Mux_h I__12194 (
            .O(N__49234),
            .I(N__49175));
    InMux I__12193 (
            .O(N__49233),
            .I(N__49170));
    InMux I__12192 (
            .O(N__49232),
            .I(N__49170));
    InMux I__12191 (
            .O(N__49231),
            .I(N__49167));
    InMux I__12190 (
            .O(N__49228),
            .I(N__49158));
    InMux I__12189 (
            .O(N__49227),
            .I(N__49158));
    InMux I__12188 (
            .O(N__49226),
            .I(N__49158));
    InMux I__12187 (
            .O(N__49225),
            .I(N__49158));
    LocalMux I__12186 (
            .O(N__49222),
            .I(N__49155));
    InMux I__12185 (
            .O(N__49221),
            .I(N__49150));
    InMux I__12184 (
            .O(N__49220),
            .I(N__49150));
    Span4Mux_h I__12183 (
            .O(N__49217),
            .I(N__49145));
    LocalMux I__12182 (
            .O(N__49214),
            .I(N__49145));
    InMux I__12181 (
            .O(N__49213),
            .I(N__49142));
    InMux I__12180 (
            .O(N__49212),
            .I(N__49139));
    LocalMux I__12179 (
            .O(N__49209),
            .I(N__49136));
    InMux I__12178 (
            .O(N__49206),
            .I(N__49131));
    InMux I__12177 (
            .O(N__49205),
            .I(N__49131));
    CascadeMux I__12176 (
            .O(N__49204),
            .I(N__49125));
    CascadeMux I__12175 (
            .O(N__49203),
            .I(N__49115));
    CascadeMux I__12174 (
            .O(N__49202),
            .I(N__49112));
    InMux I__12173 (
            .O(N__49201),
            .I(N__49102));
    InMux I__12172 (
            .O(N__49200),
            .I(N__49102));
    InMux I__12171 (
            .O(N__49199),
            .I(N__49095));
    InMux I__12170 (
            .O(N__49198),
            .I(N__49095));
    InMux I__12169 (
            .O(N__49197),
            .I(N__49095));
    InMux I__12168 (
            .O(N__49196),
            .I(N__49090));
    InMux I__12167 (
            .O(N__49195),
            .I(N__49090));
    InMux I__12166 (
            .O(N__49194),
            .I(N__49079));
    InMux I__12165 (
            .O(N__49193),
            .I(N__49079));
    InMux I__12164 (
            .O(N__49192),
            .I(N__49079));
    InMux I__12163 (
            .O(N__49191),
            .I(N__49079));
    InMux I__12162 (
            .O(N__49190),
            .I(N__49079));
    InMux I__12161 (
            .O(N__49189),
            .I(N__49074));
    LocalMux I__12160 (
            .O(N__49186),
            .I(N__49071));
    LocalMux I__12159 (
            .O(N__49183),
            .I(N__49066));
    LocalMux I__12158 (
            .O(N__49178),
            .I(N__49066));
    Span4Mux_h I__12157 (
            .O(N__49175),
            .I(N__49061));
    LocalMux I__12156 (
            .O(N__49170),
            .I(N__49061));
    LocalMux I__12155 (
            .O(N__49167),
            .I(N__49056));
    LocalMux I__12154 (
            .O(N__49158),
            .I(N__49056));
    Span4Mux_v I__12153 (
            .O(N__49155),
            .I(N__49049));
    LocalMux I__12152 (
            .O(N__49150),
            .I(N__49049));
    Span4Mux_v I__12151 (
            .O(N__49145),
            .I(N__49049));
    LocalMux I__12150 (
            .O(N__49142),
            .I(N__49046));
    LocalMux I__12149 (
            .O(N__49139),
            .I(N__49043));
    Span4Mux_v I__12148 (
            .O(N__49136),
            .I(N__49040));
    LocalMux I__12147 (
            .O(N__49131),
            .I(N__49037));
    InMux I__12146 (
            .O(N__49130),
            .I(N__49030));
    InMux I__12145 (
            .O(N__49129),
            .I(N__49030));
    InMux I__12144 (
            .O(N__49128),
            .I(N__49030));
    InMux I__12143 (
            .O(N__49125),
            .I(N__49024));
    InMux I__12142 (
            .O(N__49124),
            .I(N__49024));
    InMux I__12141 (
            .O(N__49123),
            .I(N__49021));
    InMux I__12140 (
            .O(N__49122),
            .I(N__49013));
    InMux I__12139 (
            .O(N__49121),
            .I(N__49013));
    InMux I__12138 (
            .O(N__49120),
            .I(N__49013));
    CascadeMux I__12137 (
            .O(N__49119),
            .I(N__49008));
    InMux I__12136 (
            .O(N__49118),
            .I(N__49004));
    InMux I__12135 (
            .O(N__49115),
            .I(N__48993));
    InMux I__12134 (
            .O(N__49112),
            .I(N__48993));
    InMux I__12133 (
            .O(N__49111),
            .I(N__48993));
    InMux I__12132 (
            .O(N__49110),
            .I(N__48993));
    InMux I__12131 (
            .O(N__49109),
            .I(N__48993));
    InMux I__12130 (
            .O(N__49108),
            .I(N__48988));
    InMux I__12129 (
            .O(N__49107),
            .I(N__48988));
    LocalMux I__12128 (
            .O(N__49102),
            .I(N__48979));
    LocalMux I__12127 (
            .O(N__49095),
            .I(N__48979));
    LocalMux I__12126 (
            .O(N__49090),
            .I(N__48979));
    LocalMux I__12125 (
            .O(N__49079),
            .I(N__48979));
    InMux I__12124 (
            .O(N__49078),
            .I(N__48972));
    InMux I__12123 (
            .O(N__49077),
            .I(N__48972));
    LocalMux I__12122 (
            .O(N__49074),
            .I(N__48961));
    Span4Mux_v I__12121 (
            .O(N__49071),
            .I(N__48961));
    Span4Mux_v I__12120 (
            .O(N__49066),
            .I(N__48961));
    Span4Mux_v I__12119 (
            .O(N__49061),
            .I(N__48961));
    Span4Mux_v I__12118 (
            .O(N__49056),
            .I(N__48961));
    Span4Mux_h I__12117 (
            .O(N__49049),
            .I(N__48958));
    Span4Mux_v I__12116 (
            .O(N__49046),
            .I(N__48955));
    Span4Mux_v I__12115 (
            .O(N__49043),
            .I(N__48950));
    Span4Mux_v I__12114 (
            .O(N__49040),
            .I(N__48950));
    Span4Mux_v I__12113 (
            .O(N__49037),
            .I(N__48947));
    LocalMux I__12112 (
            .O(N__49030),
            .I(N__48944));
    InMux I__12111 (
            .O(N__49029),
            .I(N__48939));
    LocalMux I__12110 (
            .O(N__49024),
            .I(N__48936));
    LocalMux I__12109 (
            .O(N__49021),
            .I(N__48933));
    InMux I__12108 (
            .O(N__49020),
            .I(N__48930));
    LocalMux I__12107 (
            .O(N__49013),
            .I(N__48927));
    InMux I__12106 (
            .O(N__49012),
            .I(N__48924));
    InMux I__12105 (
            .O(N__49011),
            .I(N__48919));
    InMux I__12104 (
            .O(N__49008),
            .I(N__48919));
    InMux I__12103 (
            .O(N__49007),
            .I(N__48916));
    LocalMux I__12102 (
            .O(N__49004),
            .I(N__48913));
    LocalMux I__12101 (
            .O(N__48993),
            .I(N__48910));
    LocalMux I__12100 (
            .O(N__48988),
            .I(N__48905));
    Span4Mux_v I__12099 (
            .O(N__48979),
            .I(N__48905));
    InMux I__12098 (
            .O(N__48978),
            .I(N__48900));
    InMux I__12097 (
            .O(N__48977),
            .I(N__48900));
    LocalMux I__12096 (
            .O(N__48972),
            .I(N__48889));
    Sp12to4 I__12095 (
            .O(N__48961),
            .I(N__48889));
    Sp12to4 I__12094 (
            .O(N__48958),
            .I(N__48889));
    Sp12to4 I__12093 (
            .O(N__48955),
            .I(N__48889));
    Sp12to4 I__12092 (
            .O(N__48950),
            .I(N__48889));
    Span4Mux_h I__12091 (
            .O(N__48947),
            .I(N__48884));
    Span4Mux_h I__12090 (
            .O(N__48944),
            .I(N__48884));
    InMux I__12089 (
            .O(N__48943),
            .I(N__48879));
    InMux I__12088 (
            .O(N__48942),
            .I(N__48879));
    LocalMux I__12087 (
            .O(N__48939),
            .I(N__48868));
    Span4Mux_h I__12086 (
            .O(N__48936),
            .I(N__48868));
    Span4Mux_v I__12085 (
            .O(N__48933),
            .I(N__48868));
    LocalMux I__12084 (
            .O(N__48930),
            .I(N__48868));
    Span4Mux_h I__12083 (
            .O(N__48927),
            .I(N__48868));
    LocalMux I__12082 (
            .O(N__48924),
            .I(adc_state_0_adj_1080));
    LocalMux I__12081 (
            .O(N__48919),
            .I(adc_state_0_adj_1080));
    LocalMux I__12080 (
            .O(N__48916),
            .I(adc_state_0_adj_1080));
    Odrv4 I__12079 (
            .O(N__48913),
            .I(adc_state_0_adj_1080));
    Odrv4 I__12078 (
            .O(N__48910),
            .I(adc_state_0_adj_1080));
    Odrv4 I__12077 (
            .O(N__48905),
            .I(adc_state_0_adj_1080));
    LocalMux I__12076 (
            .O(N__48900),
            .I(adc_state_0_adj_1080));
    Odrv12 I__12075 (
            .O(N__48889),
            .I(adc_state_0_adj_1080));
    Odrv4 I__12074 (
            .O(N__48884),
            .I(adc_state_0_adj_1080));
    LocalMux I__12073 (
            .O(N__48879),
            .I(adc_state_0_adj_1080));
    Odrv4 I__12072 (
            .O(N__48868),
            .I(adc_state_0_adj_1080));
    CascadeMux I__12071 (
            .O(N__48845),
            .I(N__48842));
    InMux I__12070 (
            .O(N__48842),
            .I(N__48836));
    InMux I__12069 (
            .O(N__48841),
            .I(N__48833));
    InMux I__12068 (
            .O(N__48840),
            .I(N__48825));
    InMux I__12067 (
            .O(N__48839),
            .I(N__48825));
    LocalMux I__12066 (
            .O(N__48836),
            .I(N__48819));
    LocalMux I__12065 (
            .O(N__48833),
            .I(N__48819));
    InMux I__12064 (
            .O(N__48832),
            .I(N__48811));
    CascadeMux I__12063 (
            .O(N__48831),
            .I(N__48806));
    InMux I__12062 (
            .O(N__48830),
            .I(N__48800));
    LocalMux I__12061 (
            .O(N__48825),
            .I(N__48797));
    InMux I__12060 (
            .O(N__48824),
            .I(N__48794));
    Span4Mux_v I__12059 (
            .O(N__48819),
            .I(N__48791));
    InMux I__12058 (
            .O(N__48818),
            .I(N__48786));
    InMux I__12057 (
            .O(N__48817),
            .I(N__48786));
    InMux I__12056 (
            .O(N__48816),
            .I(N__48781));
    InMux I__12055 (
            .O(N__48815),
            .I(N__48778));
    InMux I__12054 (
            .O(N__48814),
            .I(N__48773));
    LocalMux I__12053 (
            .O(N__48811),
            .I(N__48770));
    InMux I__12052 (
            .O(N__48810),
            .I(N__48767));
    InMux I__12051 (
            .O(N__48809),
            .I(N__48764));
    InMux I__12050 (
            .O(N__48806),
            .I(N__48758));
    InMux I__12049 (
            .O(N__48805),
            .I(N__48758));
    InMux I__12048 (
            .O(N__48804),
            .I(N__48752));
    InMux I__12047 (
            .O(N__48803),
            .I(N__48749));
    LocalMux I__12046 (
            .O(N__48800),
            .I(N__48746));
    Span4Mux_h I__12045 (
            .O(N__48797),
            .I(N__48741));
    LocalMux I__12044 (
            .O(N__48794),
            .I(N__48741));
    Span4Mux_h I__12043 (
            .O(N__48791),
            .I(N__48736));
    LocalMux I__12042 (
            .O(N__48786),
            .I(N__48736));
    InMux I__12041 (
            .O(N__48785),
            .I(N__48728));
    InMux I__12040 (
            .O(N__48784),
            .I(N__48728));
    LocalMux I__12039 (
            .O(N__48781),
            .I(N__48723));
    LocalMux I__12038 (
            .O(N__48778),
            .I(N__48723));
    InMux I__12037 (
            .O(N__48777),
            .I(N__48718));
    InMux I__12036 (
            .O(N__48776),
            .I(N__48718));
    LocalMux I__12035 (
            .O(N__48773),
            .I(N__48715));
    Span4Mux_v I__12034 (
            .O(N__48770),
            .I(N__48712));
    LocalMux I__12033 (
            .O(N__48767),
            .I(N__48707));
    LocalMux I__12032 (
            .O(N__48764),
            .I(N__48707));
    InMux I__12031 (
            .O(N__48763),
            .I(N__48704));
    LocalMux I__12030 (
            .O(N__48758),
            .I(N__48701));
    InMux I__12029 (
            .O(N__48757),
            .I(N__48698));
    InMux I__12028 (
            .O(N__48756),
            .I(N__48693));
    InMux I__12027 (
            .O(N__48755),
            .I(N__48693));
    LocalMux I__12026 (
            .O(N__48752),
            .I(N__48686));
    LocalMux I__12025 (
            .O(N__48749),
            .I(N__48686));
    Span4Mux_h I__12024 (
            .O(N__48746),
            .I(N__48686));
    Span4Mux_h I__12023 (
            .O(N__48741),
            .I(N__48681));
    Span4Mux_h I__12022 (
            .O(N__48736),
            .I(N__48681));
    InMux I__12021 (
            .O(N__48735),
            .I(N__48671));
    InMux I__12020 (
            .O(N__48734),
            .I(N__48671));
    InMux I__12019 (
            .O(N__48733),
            .I(N__48671));
    LocalMux I__12018 (
            .O(N__48728),
            .I(N__48668));
    Span4Mux_v I__12017 (
            .O(N__48723),
            .I(N__48661));
    LocalMux I__12016 (
            .O(N__48718),
            .I(N__48661));
    Span4Mux_h I__12015 (
            .O(N__48715),
            .I(N__48661));
    Sp12to4 I__12014 (
            .O(N__48712),
            .I(N__48658));
    Span4Mux_v I__12013 (
            .O(N__48707),
            .I(N__48655));
    LocalMux I__12012 (
            .O(N__48704),
            .I(N__48652));
    Span4Mux_h I__12011 (
            .O(N__48701),
            .I(N__48649));
    LocalMux I__12010 (
            .O(N__48698),
            .I(N__48640));
    LocalMux I__12009 (
            .O(N__48693),
            .I(N__48640));
    Span4Mux_h I__12008 (
            .O(N__48686),
            .I(N__48640));
    Span4Mux_v I__12007 (
            .O(N__48681),
            .I(N__48640));
    InMux I__12006 (
            .O(N__48680),
            .I(N__48637));
    InMux I__12005 (
            .O(N__48679),
            .I(N__48632));
    InMux I__12004 (
            .O(N__48678),
            .I(N__48632));
    LocalMux I__12003 (
            .O(N__48671),
            .I(N__48627));
    Span4Mux_h I__12002 (
            .O(N__48668),
            .I(N__48627));
    Span4Mux_v I__12001 (
            .O(N__48661),
            .I(N__48624));
    Span12Mux_s9_v I__12000 (
            .O(N__48658),
            .I(N__48619));
    Sp12to4 I__11999 (
            .O(N__48655),
            .I(N__48619));
    Span4Mux_v I__11998 (
            .O(N__48652),
            .I(N__48612));
    Span4Mux_v I__11997 (
            .O(N__48649),
            .I(N__48612));
    Span4Mux_h I__11996 (
            .O(N__48640),
            .I(N__48612));
    LocalMux I__11995 (
            .O(N__48637),
            .I(n8332));
    LocalMux I__11994 (
            .O(N__48632),
            .I(n8332));
    Odrv4 I__11993 (
            .O(N__48627),
            .I(n8332));
    Odrv4 I__11992 (
            .O(N__48624),
            .I(n8332));
    Odrv12 I__11991 (
            .O(N__48619),
            .I(n8332));
    Odrv4 I__11990 (
            .O(N__48612),
            .I(n8332));
    CascadeMux I__11989 (
            .O(N__48599),
            .I(N__48595));
    InMux I__11988 (
            .O(N__48598),
            .I(N__48590));
    InMux I__11987 (
            .O(N__48595),
            .I(N__48590));
    LocalMux I__11986 (
            .O(N__48590),
            .I(N__48586));
    CascadeMux I__11985 (
            .O(N__48589),
            .I(N__48583));
    Span12Mux_h I__11984 (
            .O(N__48586),
            .I(N__48580));
    InMux I__11983 (
            .O(N__48583),
            .I(N__48577));
    Odrv12 I__11982 (
            .O(N__48580),
            .I(cmd_rdadctmp_20_adj_1092));
    LocalMux I__11981 (
            .O(N__48577),
            .I(cmd_rdadctmp_20_adj_1092));
    InMux I__11980 (
            .O(N__48572),
            .I(N__48569));
    LocalMux I__11979 (
            .O(N__48569),
            .I(N__48566));
    Odrv12 I__11978 (
            .O(N__48566),
            .I(n15640));
    CascadeMux I__11977 (
            .O(N__48563),
            .I(N__48560));
    InMux I__11976 (
            .O(N__48560),
            .I(N__48557));
    LocalMux I__11975 (
            .O(N__48557),
            .I(N__48554));
    Span12Mux_v I__11974 (
            .O(N__48554),
            .I(N__48551));
    Odrv12 I__11973 (
            .O(N__48551),
            .I(n10_adj_1172));
    CEMux I__11972 (
            .O(N__48548),
            .I(N__48539));
    CascadeMux I__11971 (
            .O(N__48547),
            .I(N__48533));
    CascadeMux I__11970 (
            .O(N__48546),
            .I(N__48530));
    InMux I__11969 (
            .O(N__48545),
            .I(N__48510));
    InMux I__11968 (
            .O(N__48544),
            .I(N__48510));
    InMux I__11967 (
            .O(N__48543),
            .I(N__48510));
    InMux I__11966 (
            .O(N__48542),
            .I(N__48507));
    LocalMux I__11965 (
            .O(N__48539),
            .I(N__48500));
    SRMux I__11964 (
            .O(N__48538),
            .I(N__48497));
    InMux I__11963 (
            .O(N__48537),
            .I(N__48494));
    InMux I__11962 (
            .O(N__48536),
            .I(N__48477));
    InMux I__11961 (
            .O(N__48533),
            .I(N__48477));
    InMux I__11960 (
            .O(N__48530),
            .I(N__48477));
    InMux I__11959 (
            .O(N__48529),
            .I(N__48477));
    InMux I__11958 (
            .O(N__48528),
            .I(N__48477));
    InMux I__11957 (
            .O(N__48527),
            .I(N__48477));
    InMux I__11956 (
            .O(N__48526),
            .I(N__48477));
    InMux I__11955 (
            .O(N__48525),
            .I(N__48477));
    InMux I__11954 (
            .O(N__48524),
            .I(N__48460));
    InMux I__11953 (
            .O(N__48523),
            .I(N__48460));
    InMux I__11952 (
            .O(N__48522),
            .I(N__48460));
    InMux I__11951 (
            .O(N__48521),
            .I(N__48460));
    InMux I__11950 (
            .O(N__48520),
            .I(N__48460));
    InMux I__11949 (
            .O(N__48519),
            .I(N__48460));
    InMux I__11948 (
            .O(N__48518),
            .I(N__48460));
    InMux I__11947 (
            .O(N__48517),
            .I(N__48460));
    LocalMux I__11946 (
            .O(N__48510),
            .I(N__48457));
    LocalMux I__11945 (
            .O(N__48507),
            .I(N__48454));
    InMux I__11944 (
            .O(N__48506),
            .I(N__48445));
    InMux I__11943 (
            .O(N__48505),
            .I(N__48445));
    InMux I__11942 (
            .O(N__48504),
            .I(N__48445));
    InMux I__11941 (
            .O(N__48503),
            .I(N__48445));
    Span4Mux_v I__11940 (
            .O(N__48500),
            .I(N__48442));
    LocalMux I__11939 (
            .O(N__48497),
            .I(N__48439));
    LocalMux I__11938 (
            .O(N__48494),
            .I(N__48436));
    LocalMux I__11937 (
            .O(N__48477),
            .I(N__48431));
    LocalMux I__11936 (
            .O(N__48460),
            .I(N__48431));
    Span4Mux_h I__11935 (
            .O(N__48457),
            .I(N__48424));
    Span4Mux_h I__11934 (
            .O(N__48454),
            .I(N__48424));
    LocalMux I__11933 (
            .O(N__48445),
            .I(N__48424));
    Span4Mux_h I__11932 (
            .O(N__48442),
            .I(N__48421));
    Span4Mux_v I__11931 (
            .O(N__48439),
            .I(N__48413));
    Span4Mux_h I__11930 (
            .O(N__48436),
            .I(N__48413));
    Span4Mux_h I__11929 (
            .O(N__48431),
            .I(N__48413));
    Span4Mux_h I__11928 (
            .O(N__48424),
            .I(N__48410));
    Span4Mux_v I__11927 (
            .O(N__48421),
            .I(N__48407));
    InMux I__11926 (
            .O(N__48420),
            .I(N__48404));
    Span4Mux_v I__11925 (
            .O(N__48413),
            .I(N__48401));
    Span4Mux_v I__11924 (
            .O(N__48410),
            .I(N__48398));
    Odrv4 I__11923 (
            .O(N__48407),
            .I(dds_state_1));
    LocalMux I__11922 (
            .O(N__48404),
            .I(dds_state_1));
    Odrv4 I__11921 (
            .O(N__48401),
            .I(dds_state_1));
    Odrv4 I__11920 (
            .O(N__48398),
            .I(dds_state_1));
    CascadeMux I__11919 (
            .O(N__48389),
            .I(N__48384));
    InMux I__11918 (
            .O(N__48388),
            .I(N__48377));
    InMux I__11917 (
            .O(N__48387),
            .I(N__48374));
    InMux I__11916 (
            .O(N__48384),
            .I(N__48367));
    InMux I__11915 (
            .O(N__48383),
            .I(N__48367));
    InMux I__11914 (
            .O(N__48382),
            .I(N__48367));
    InMux I__11913 (
            .O(N__48381),
            .I(N__48364));
    InMux I__11912 (
            .O(N__48380),
            .I(N__48360));
    LocalMux I__11911 (
            .O(N__48377),
            .I(N__48357));
    LocalMux I__11910 (
            .O(N__48374),
            .I(N__48352));
    LocalMux I__11909 (
            .O(N__48367),
            .I(N__48352));
    LocalMux I__11908 (
            .O(N__48364),
            .I(N__48349));
    InMux I__11907 (
            .O(N__48363),
            .I(N__48346));
    LocalMux I__11906 (
            .O(N__48360),
            .I(N__48343));
    Span4Mux_v I__11905 (
            .O(N__48357),
            .I(N__48340));
    Span4Mux_v I__11904 (
            .O(N__48352),
            .I(N__48335));
    Span4Mux_h I__11903 (
            .O(N__48349),
            .I(N__48335));
    LocalMux I__11902 (
            .O(N__48346),
            .I(N__48331));
    Span4Mux_h I__11901 (
            .O(N__48343),
            .I(N__48328));
    Span4Mux_h I__11900 (
            .O(N__48340),
            .I(N__48325));
    Span4Mux_h I__11899 (
            .O(N__48335),
            .I(N__48322));
    InMux I__11898 (
            .O(N__48334),
            .I(N__48319));
    Span12Mux_h I__11897 (
            .O(N__48331),
            .I(N__48316));
    Span4Mux_v I__11896 (
            .O(N__48328),
            .I(N__48311));
    Span4Mux_h I__11895 (
            .O(N__48325),
            .I(N__48311));
    Span4Mux_h I__11894 (
            .O(N__48322),
            .I(N__48308));
    LocalMux I__11893 (
            .O(N__48319),
            .I(dds_state_0));
    Odrv12 I__11892 (
            .O(N__48316),
            .I(dds_state_0));
    Odrv4 I__11891 (
            .O(N__48311),
            .I(dds_state_0));
    Odrv4 I__11890 (
            .O(N__48308),
            .I(dds_state_0));
    CEMux I__11889 (
            .O(N__48299),
            .I(N__48295));
    CEMux I__11888 (
            .O(N__48298),
            .I(N__48292));
    LocalMux I__11887 (
            .O(N__48295),
            .I(N__48289));
    LocalMux I__11886 (
            .O(N__48292),
            .I(N__48286));
    Span4Mux_h I__11885 (
            .O(N__48289),
            .I(N__48283));
    Span4Mux_h I__11884 (
            .O(N__48286),
            .I(N__48280));
    Sp12to4 I__11883 (
            .O(N__48283),
            .I(N__48277));
    Odrv4 I__11882 (
            .O(N__48280),
            .I(\CLOCK_DDS.n9 ));
    Odrv12 I__11881 (
            .O(N__48277),
            .I(\CLOCK_DDS.n9 ));
    CascadeMux I__11880 (
            .O(N__48272),
            .I(N__48269));
    InMux I__11879 (
            .O(N__48269),
            .I(N__48266));
    LocalMux I__11878 (
            .O(N__48266),
            .I(N__48263));
    Span4Mux_v I__11877 (
            .O(N__48263),
            .I(N__48260));
    Span4Mux_h I__11876 (
            .O(N__48260),
            .I(N__48256));
    InMux I__11875 (
            .O(N__48259),
            .I(N__48253));
    Span4Mux_h I__11874 (
            .O(N__48256),
            .I(N__48249));
    LocalMux I__11873 (
            .O(N__48253),
            .I(N__48246));
    CascadeMux I__11872 (
            .O(N__48252),
            .I(N__48243));
    Span4Mux_h I__11871 (
            .O(N__48249),
            .I(N__48240));
    Span4Mux_h I__11870 (
            .O(N__48246),
            .I(N__48237));
    InMux I__11869 (
            .O(N__48243),
            .I(N__48234));
    Odrv4 I__11868 (
            .O(N__48240),
            .I(cmd_rdadctmp_24));
    Odrv4 I__11867 (
            .O(N__48237),
            .I(cmd_rdadctmp_24));
    LocalMux I__11866 (
            .O(N__48234),
            .I(cmd_rdadctmp_24));
    InMux I__11865 (
            .O(N__48227),
            .I(N__48223));
    InMux I__11864 (
            .O(N__48226),
            .I(N__48220));
    LocalMux I__11863 (
            .O(N__48223),
            .I(N__48217));
    LocalMux I__11862 (
            .O(N__48220),
            .I(buf_adcdata1_16));
    Odrv4 I__11861 (
            .O(N__48217),
            .I(buf_adcdata1_16));
    InMux I__11860 (
            .O(N__48212),
            .I(N__48209));
    LocalMux I__11859 (
            .O(N__48209),
            .I(N__48206));
    Span4Mux_v I__11858 (
            .O(N__48206),
            .I(N__48203));
    Span4Mux_h I__11857 (
            .O(N__48203),
            .I(N__48198));
    CascadeMux I__11856 (
            .O(N__48202),
            .I(N__48195));
    InMux I__11855 (
            .O(N__48201),
            .I(N__48192));
    Span4Mux_h I__11854 (
            .O(N__48198),
            .I(N__48189));
    InMux I__11853 (
            .O(N__48195),
            .I(N__48186));
    LocalMux I__11852 (
            .O(N__48192),
            .I(cmd_rdadctmp_30_adj_1046));
    Odrv4 I__11851 (
            .O(N__48189),
            .I(cmd_rdadctmp_30_adj_1046));
    LocalMux I__11850 (
            .O(N__48186),
            .I(cmd_rdadctmp_30_adj_1046));
    InMux I__11849 (
            .O(N__48179),
            .I(N__48176));
    LocalMux I__11848 (
            .O(N__48176),
            .I(N__48173));
    Span4Mux_v I__11847 (
            .O(N__48173),
            .I(N__48169));
    InMux I__11846 (
            .O(N__48172),
            .I(N__48166));
    Span4Mux_v I__11845 (
            .O(N__48169),
            .I(N__48163));
    LocalMux I__11844 (
            .O(N__48166),
            .I(buf_adcdata2_22));
    Odrv4 I__11843 (
            .O(N__48163),
            .I(buf_adcdata2_22));
    CascadeMux I__11842 (
            .O(N__48158),
            .I(N__48155));
    InMux I__11841 (
            .O(N__48155),
            .I(N__48152));
    LocalMux I__11840 (
            .O(N__48152),
            .I(N__48149));
    Span4Mux_h I__11839 (
            .O(N__48149),
            .I(N__48146));
    Span4Mux_h I__11838 (
            .O(N__48146),
            .I(N__48143));
    Span4Mux_v I__11837 (
            .O(N__48143),
            .I(N__48140));
    Span4Mux_h I__11836 (
            .O(N__48140),
            .I(N__48136));
    CascadeMux I__11835 (
            .O(N__48139),
            .I(N__48133));
    Span4Mux_h I__11834 (
            .O(N__48136),
            .I(N__48130));
    InMux I__11833 (
            .O(N__48133),
            .I(N__48127));
    Odrv4 I__11832 (
            .O(N__48130),
            .I(cmd_rdadctmp_31_adj_1045));
    LocalMux I__11831 (
            .O(N__48127),
            .I(cmd_rdadctmp_31_adj_1045));
    InMux I__11830 (
            .O(N__48122),
            .I(N__48119));
    LocalMux I__11829 (
            .O(N__48119),
            .I(N__48115));
    InMux I__11828 (
            .O(N__48118),
            .I(N__48112));
    Span4Mux_v I__11827 (
            .O(N__48115),
            .I(N__48109));
    LocalMux I__11826 (
            .O(N__48112),
            .I(buf_adcdata2_23));
    Odrv4 I__11825 (
            .O(N__48109),
            .I(buf_adcdata2_23));
    InMux I__11824 (
            .O(N__48104),
            .I(N__48101));
    LocalMux I__11823 (
            .O(N__48101),
            .I(N__48098));
    Span4Mux_v I__11822 (
            .O(N__48098),
            .I(N__48095));
    Odrv4 I__11821 (
            .O(N__48095),
            .I(buf_data2_16));
    CascadeMux I__11820 (
            .O(N__48092),
            .I(N__48088));
    InMux I__11819 (
            .O(N__48091),
            .I(N__48080));
    InMux I__11818 (
            .O(N__48088),
            .I(N__48075));
    InMux I__11817 (
            .O(N__48087),
            .I(N__48075));
    CascadeMux I__11816 (
            .O(N__48086),
            .I(N__48064));
    CascadeMux I__11815 (
            .O(N__48085),
            .I(N__48061));
    InMux I__11814 (
            .O(N__48084),
            .I(N__48057));
    InMux I__11813 (
            .O(N__48083),
            .I(N__48054));
    LocalMux I__11812 (
            .O(N__48080),
            .I(N__48049));
    LocalMux I__11811 (
            .O(N__48075),
            .I(N__48049));
    InMux I__11810 (
            .O(N__48074),
            .I(N__48043));
    InMux I__11809 (
            .O(N__48073),
            .I(N__48030));
    InMux I__11808 (
            .O(N__48072),
            .I(N__48030));
    InMux I__11807 (
            .O(N__48071),
            .I(N__48023));
    InMux I__11806 (
            .O(N__48070),
            .I(N__48023));
    InMux I__11805 (
            .O(N__48069),
            .I(N__48023));
    InMux I__11804 (
            .O(N__48068),
            .I(N__48020));
    InMux I__11803 (
            .O(N__48067),
            .I(N__48015));
    InMux I__11802 (
            .O(N__48064),
            .I(N__48015));
    InMux I__11801 (
            .O(N__48061),
            .I(N__48007));
    InMux I__11800 (
            .O(N__48060),
            .I(N__48007));
    LocalMux I__11799 (
            .O(N__48057),
            .I(N__48001));
    LocalMux I__11798 (
            .O(N__48054),
            .I(N__47996));
    Span4Mux_h I__11797 (
            .O(N__48049),
            .I(N__47996));
    InMux I__11796 (
            .O(N__48048),
            .I(N__47993));
    CascadeMux I__11795 (
            .O(N__48047),
            .I(N__47990));
    CascadeMux I__11794 (
            .O(N__48046),
            .I(N__47986));
    LocalMux I__11793 (
            .O(N__48043),
            .I(N__47980));
    InMux I__11792 (
            .O(N__48042),
            .I(N__47977));
    InMux I__11791 (
            .O(N__48041),
            .I(N__47974));
    InMux I__11790 (
            .O(N__48040),
            .I(N__47971));
    InMux I__11789 (
            .O(N__48039),
            .I(N__47966));
    InMux I__11788 (
            .O(N__48038),
            .I(N__47966));
    InMux I__11787 (
            .O(N__48037),
            .I(N__47963));
    InMux I__11786 (
            .O(N__48036),
            .I(N__47958));
    InMux I__11785 (
            .O(N__48035),
            .I(N__47958));
    LocalMux I__11784 (
            .O(N__48030),
            .I(N__47955));
    LocalMux I__11783 (
            .O(N__48023),
            .I(N__47948));
    LocalMux I__11782 (
            .O(N__48020),
            .I(N__47948));
    LocalMux I__11781 (
            .O(N__48015),
            .I(N__47948));
    InMux I__11780 (
            .O(N__48014),
            .I(N__47945));
    InMux I__11779 (
            .O(N__48013),
            .I(N__47941));
    InMux I__11778 (
            .O(N__48012),
            .I(N__47938));
    LocalMux I__11777 (
            .O(N__48007),
            .I(N__47935));
    InMux I__11776 (
            .O(N__48006),
            .I(N__47930));
    InMux I__11775 (
            .O(N__48005),
            .I(N__47930));
    InMux I__11774 (
            .O(N__48004),
            .I(N__47925));
    Span4Mux_v I__11773 (
            .O(N__48001),
            .I(N__47902));
    Span4Mux_h I__11772 (
            .O(N__47996),
            .I(N__47902));
    LocalMux I__11771 (
            .O(N__47993),
            .I(N__47902));
    InMux I__11770 (
            .O(N__47990),
            .I(N__47895));
    InMux I__11769 (
            .O(N__47989),
            .I(N__47895));
    InMux I__11768 (
            .O(N__47986),
            .I(N__47895));
    InMux I__11767 (
            .O(N__47985),
            .I(N__47888));
    InMux I__11766 (
            .O(N__47984),
            .I(N__47888));
    InMux I__11765 (
            .O(N__47983),
            .I(N__47888));
    Span4Mux_h I__11764 (
            .O(N__47980),
            .I(N__47877));
    LocalMux I__11763 (
            .O(N__47977),
            .I(N__47877));
    LocalMux I__11762 (
            .O(N__47974),
            .I(N__47877));
    LocalMux I__11761 (
            .O(N__47971),
            .I(N__47877));
    LocalMux I__11760 (
            .O(N__47966),
            .I(N__47877));
    LocalMux I__11759 (
            .O(N__47963),
            .I(N__47866));
    LocalMux I__11758 (
            .O(N__47958),
            .I(N__47866));
    Span4Mux_v I__11757 (
            .O(N__47955),
            .I(N__47866));
    Span4Mux_v I__11756 (
            .O(N__47948),
            .I(N__47866));
    LocalMux I__11755 (
            .O(N__47945),
            .I(N__47866));
    InMux I__11754 (
            .O(N__47944),
            .I(N__47861));
    LocalMux I__11753 (
            .O(N__47941),
            .I(N__47856));
    LocalMux I__11752 (
            .O(N__47938),
            .I(N__47849));
    Span4Mux_v I__11751 (
            .O(N__47935),
            .I(N__47844));
    LocalMux I__11750 (
            .O(N__47930),
            .I(N__47844));
    InMux I__11749 (
            .O(N__47929),
            .I(N__47841));
    InMux I__11748 (
            .O(N__47928),
            .I(N__47838));
    LocalMux I__11747 (
            .O(N__47925),
            .I(N__47835));
    InMux I__11746 (
            .O(N__47924),
            .I(N__47828));
    InMux I__11745 (
            .O(N__47923),
            .I(N__47828));
    InMux I__11744 (
            .O(N__47922),
            .I(N__47828));
    InMux I__11743 (
            .O(N__47921),
            .I(N__47825));
    InMux I__11742 (
            .O(N__47920),
            .I(N__47817));
    InMux I__11741 (
            .O(N__47919),
            .I(N__47817));
    CascadeMux I__11740 (
            .O(N__47918),
            .I(N__47812));
    InMux I__11739 (
            .O(N__47917),
            .I(N__47807));
    InMux I__11738 (
            .O(N__47916),
            .I(N__47787));
    InMux I__11737 (
            .O(N__47915),
            .I(N__47776));
    InMux I__11736 (
            .O(N__47914),
            .I(N__47776));
    InMux I__11735 (
            .O(N__47913),
            .I(N__47776));
    InMux I__11734 (
            .O(N__47912),
            .I(N__47776));
    InMux I__11733 (
            .O(N__47911),
            .I(N__47776));
    InMux I__11732 (
            .O(N__47910),
            .I(N__47771));
    InMux I__11731 (
            .O(N__47909),
            .I(N__47771));
    Span4Mux_h I__11730 (
            .O(N__47902),
            .I(N__47764));
    LocalMux I__11729 (
            .O(N__47895),
            .I(N__47764));
    LocalMux I__11728 (
            .O(N__47888),
            .I(N__47764));
    Span4Mux_v I__11727 (
            .O(N__47877),
            .I(N__47759));
    Span4Mux_h I__11726 (
            .O(N__47866),
            .I(N__47759));
    InMux I__11725 (
            .O(N__47865),
            .I(N__47754));
    InMux I__11724 (
            .O(N__47864),
            .I(N__47754));
    LocalMux I__11723 (
            .O(N__47861),
            .I(N__47751));
    InMux I__11722 (
            .O(N__47860),
            .I(N__47746));
    InMux I__11721 (
            .O(N__47859),
            .I(N__47746));
    Span4Mux_h I__11720 (
            .O(N__47856),
            .I(N__47738));
    InMux I__11719 (
            .O(N__47855),
            .I(N__47735));
    InMux I__11718 (
            .O(N__47854),
            .I(N__47732));
    InMux I__11717 (
            .O(N__47853),
            .I(N__47727));
    InMux I__11716 (
            .O(N__47852),
            .I(N__47727));
    Span4Mux_v I__11715 (
            .O(N__47849),
            .I(N__47722));
    Span4Mux_h I__11714 (
            .O(N__47844),
            .I(N__47722));
    LocalMux I__11713 (
            .O(N__47841),
            .I(N__47719));
    LocalMux I__11712 (
            .O(N__47838),
            .I(N__47716));
    Span4Mux_h I__11711 (
            .O(N__47835),
            .I(N__47711));
    LocalMux I__11710 (
            .O(N__47828),
            .I(N__47711));
    LocalMux I__11709 (
            .O(N__47825),
            .I(N__47708));
    InMux I__11708 (
            .O(N__47824),
            .I(N__47703));
    InMux I__11707 (
            .O(N__47823),
            .I(N__47703));
    InMux I__11706 (
            .O(N__47822),
            .I(N__47697));
    LocalMux I__11705 (
            .O(N__47817),
            .I(N__47694));
    InMux I__11704 (
            .O(N__47816),
            .I(N__47687));
    InMux I__11703 (
            .O(N__47815),
            .I(N__47687));
    InMux I__11702 (
            .O(N__47812),
            .I(N__47687));
    InMux I__11701 (
            .O(N__47811),
            .I(N__47684));
    InMux I__11700 (
            .O(N__47810),
            .I(N__47681));
    LocalMux I__11699 (
            .O(N__47807),
            .I(N__47678));
    InMux I__11698 (
            .O(N__47806),
            .I(N__47671));
    InMux I__11697 (
            .O(N__47805),
            .I(N__47671));
    InMux I__11696 (
            .O(N__47804),
            .I(N__47671));
    InMux I__11695 (
            .O(N__47803),
            .I(N__47667));
    InMux I__11694 (
            .O(N__47802),
            .I(N__47664));
    InMux I__11693 (
            .O(N__47801),
            .I(N__47659));
    InMux I__11692 (
            .O(N__47800),
            .I(N__47659));
    InMux I__11691 (
            .O(N__47799),
            .I(N__47654));
    InMux I__11690 (
            .O(N__47798),
            .I(N__47654));
    InMux I__11689 (
            .O(N__47797),
            .I(N__47647));
    InMux I__11688 (
            .O(N__47796),
            .I(N__47647));
    InMux I__11687 (
            .O(N__47795),
            .I(N__47647));
    InMux I__11686 (
            .O(N__47794),
            .I(N__47640));
    InMux I__11685 (
            .O(N__47793),
            .I(N__47640));
    InMux I__11684 (
            .O(N__47792),
            .I(N__47640));
    InMux I__11683 (
            .O(N__47791),
            .I(N__47637));
    CascadeMux I__11682 (
            .O(N__47790),
            .I(N__47633));
    LocalMux I__11681 (
            .O(N__47787),
            .I(N__47620));
    LocalMux I__11680 (
            .O(N__47776),
            .I(N__47620));
    LocalMux I__11679 (
            .O(N__47771),
            .I(N__47620));
    Span4Mux_v I__11678 (
            .O(N__47764),
            .I(N__47620));
    Span4Mux_h I__11677 (
            .O(N__47759),
            .I(N__47620));
    LocalMux I__11676 (
            .O(N__47754),
            .I(N__47620));
    Span4Mux_h I__11675 (
            .O(N__47751),
            .I(N__47615));
    LocalMux I__11674 (
            .O(N__47746),
            .I(N__47615));
    InMux I__11673 (
            .O(N__47745),
            .I(N__47606));
    InMux I__11672 (
            .O(N__47744),
            .I(N__47606));
    InMux I__11671 (
            .O(N__47743),
            .I(N__47606));
    InMux I__11670 (
            .O(N__47742),
            .I(N__47606));
    CascadeMux I__11669 (
            .O(N__47741),
            .I(N__47596));
    Span4Mux_h I__11668 (
            .O(N__47738),
            .I(N__47588));
    LocalMux I__11667 (
            .O(N__47735),
            .I(N__47588));
    LocalMux I__11666 (
            .O(N__47732),
            .I(N__47585));
    LocalMux I__11665 (
            .O(N__47727),
            .I(N__47580));
    Span4Mux_h I__11664 (
            .O(N__47722),
            .I(N__47580));
    Span4Mux_h I__11663 (
            .O(N__47719),
            .I(N__47577));
    Span4Mux_v I__11662 (
            .O(N__47716),
            .I(N__47572));
    Span4Mux_h I__11661 (
            .O(N__47711),
            .I(N__47572));
    Span4Mux_h I__11660 (
            .O(N__47708),
            .I(N__47567));
    LocalMux I__11659 (
            .O(N__47703),
            .I(N__47567));
    InMux I__11658 (
            .O(N__47702),
            .I(N__47564));
    InMux I__11657 (
            .O(N__47701),
            .I(N__47559));
    InMux I__11656 (
            .O(N__47700),
            .I(N__47559));
    LocalMux I__11655 (
            .O(N__47697),
            .I(N__47544));
    Span4Mux_h I__11654 (
            .O(N__47694),
            .I(N__47544));
    LocalMux I__11653 (
            .O(N__47687),
            .I(N__47544));
    LocalMux I__11652 (
            .O(N__47684),
            .I(N__47544));
    LocalMux I__11651 (
            .O(N__47681),
            .I(N__47544));
    Span4Mux_h I__11650 (
            .O(N__47678),
            .I(N__47544));
    LocalMux I__11649 (
            .O(N__47671),
            .I(N__47544));
    CascadeMux I__11648 (
            .O(N__47670),
            .I(N__47537));
    LocalMux I__11647 (
            .O(N__47667),
            .I(N__47522));
    LocalMux I__11646 (
            .O(N__47664),
            .I(N__47522));
    LocalMux I__11645 (
            .O(N__47659),
            .I(N__47522));
    LocalMux I__11644 (
            .O(N__47654),
            .I(N__47522));
    LocalMux I__11643 (
            .O(N__47647),
            .I(N__47522));
    LocalMux I__11642 (
            .O(N__47640),
            .I(N__47522));
    LocalMux I__11641 (
            .O(N__47637),
            .I(N__47522));
    InMux I__11640 (
            .O(N__47636),
            .I(N__47517));
    InMux I__11639 (
            .O(N__47633),
            .I(N__47517));
    Span4Mux_v I__11638 (
            .O(N__47620),
            .I(N__47510));
    Span4Mux_v I__11637 (
            .O(N__47615),
            .I(N__47510));
    LocalMux I__11636 (
            .O(N__47606),
            .I(N__47510));
    InMux I__11635 (
            .O(N__47605),
            .I(N__47504));
    InMux I__11634 (
            .O(N__47604),
            .I(N__47497));
    InMux I__11633 (
            .O(N__47603),
            .I(N__47497));
    InMux I__11632 (
            .O(N__47602),
            .I(N__47497));
    CascadeMux I__11631 (
            .O(N__47601),
            .I(N__47492));
    InMux I__11630 (
            .O(N__47600),
            .I(N__47485));
    InMux I__11629 (
            .O(N__47599),
            .I(N__47480));
    InMux I__11628 (
            .O(N__47596),
            .I(N__47480));
    InMux I__11627 (
            .O(N__47595),
            .I(N__47473));
    InMux I__11626 (
            .O(N__47594),
            .I(N__47473));
    InMux I__11625 (
            .O(N__47593),
            .I(N__47473));
    Span4Mux_h I__11624 (
            .O(N__47588),
            .I(N__47470));
    Span4Mux_h I__11623 (
            .O(N__47585),
            .I(N__47459));
    Span4Mux_h I__11622 (
            .O(N__47580),
            .I(N__47459));
    Span4Mux_v I__11621 (
            .O(N__47577),
            .I(N__47459));
    Span4Mux_v I__11620 (
            .O(N__47572),
            .I(N__47459));
    Span4Mux_h I__11619 (
            .O(N__47567),
            .I(N__47459));
    LocalMux I__11618 (
            .O(N__47564),
            .I(N__47452));
    LocalMux I__11617 (
            .O(N__47559),
            .I(N__47452));
    Span4Mux_v I__11616 (
            .O(N__47544),
            .I(N__47452));
    InMux I__11615 (
            .O(N__47543),
            .I(N__47447));
    InMux I__11614 (
            .O(N__47542),
            .I(N__47447));
    InMux I__11613 (
            .O(N__47541),
            .I(N__47440));
    InMux I__11612 (
            .O(N__47540),
            .I(N__47440));
    InMux I__11611 (
            .O(N__47537),
            .I(N__47440));
    Span4Mux_v I__11610 (
            .O(N__47522),
            .I(N__47433));
    LocalMux I__11609 (
            .O(N__47517),
            .I(N__47433));
    Span4Mux_h I__11608 (
            .O(N__47510),
            .I(N__47433));
    InMux I__11607 (
            .O(N__47509),
            .I(N__47426));
    InMux I__11606 (
            .O(N__47508),
            .I(N__47426));
    InMux I__11605 (
            .O(N__47507),
            .I(N__47426));
    LocalMux I__11604 (
            .O(N__47504),
            .I(N__47421));
    LocalMux I__11603 (
            .O(N__47497),
            .I(N__47421));
    InMux I__11602 (
            .O(N__47496),
            .I(N__47412));
    InMux I__11601 (
            .O(N__47495),
            .I(N__47412));
    InMux I__11600 (
            .O(N__47492),
            .I(N__47412));
    InMux I__11599 (
            .O(N__47491),
            .I(N__47412));
    InMux I__11598 (
            .O(N__47490),
            .I(N__47405));
    InMux I__11597 (
            .O(N__47489),
            .I(N__47405));
    InMux I__11596 (
            .O(N__47488),
            .I(N__47405));
    LocalMux I__11595 (
            .O(N__47485),
            .I(comm_cmd_0));
    LocalMux I__11594 (
            .O(N__47480),
            .I(comm_cmd_0));
    LocalMux I__11593 (
            .O(N__47473),
            .I(comm_cmd_0));
    Odrv4 I__11592 (
            .O(N__47470),
            .I(comm_cmd_0));
    Odrv4 I__11591 (
            .O(N__47459),
            .I(comm_cmd_0));
    Odrv4 I__11590 (
            .O(N__47452),
            .I(comm_cmd_0));
    LocalMux I__11589 (
            .O(N__47447),
            .I(comm_cmd_0));
    LocalMux I__11588 (
            .O(N__47440),
            .I(comm_cmd_0));
    Odrv4 I__11587 (
            .O(N__47433),
            .I(comm_cmd_0));
    LocalMux I__11586 (
            .O(N__47426),
            .I(comm_cmd_0));
    Odrv4 I__11585 (
            .O(N__47421),
            .I(comm_cmd_0));
    LocalMux I__11584 (
            .O(N__47412),
            .I(comm_cmd_0));
    LocalMux I__11583 (
            .O(N__47405),
            .I(comm_cmd_0));
    CascadeMux I__11582 (
            .O(N__47378),
            .I(N__47375));
    InMux I__11581 (
            .O(N__47375),
            .I(N__47372));
    LocalMux I__11580 (
            .O(N__47372),
            .I(N__47368));
    InMux I__11579 (
            .O(N__47371),
            .I(N__47365));
    Span4Mux_v I__11578 (
            .O(N__47368),
            .I(N__47360));
    LocalMux I__11577 (
            .O(N__47365),
            .I(N__47360));
    Span4Mux_v I__11576 (
            .O(N__47360),
            .I(N__47356));
    CascadeMux I__11575 (
            .O(N__47359),
            .I(N__47353));
    Span4Mux_h I__11574 (
            .O(N__47356),
            .I(N__47350));
    InMux I__11573 (
            .O(N__47353),
            .I(N__47347));
    Span4Mux_h I__11572 (
            .O(N__47350),
            .I(N__47344));
    LocalMux I__11571 (
            .O(N__47347),
            .I(buf_adcdata4_16));
    Odrv4 I__11570 (
            .O(N__47344),
            .I(buf_adcdata4_16));
    InMux I__11569 (
            .O(N__47339),
            .I(N__47330));
    InMux I__11568 (
            .O(N__47338),
            .I(N__47330));
    InMux I__11567 (
            .O(N__47337),
            .I(N__47327));
    CascadeMux I__11566 (
            .O(N__47336),
            .I(N__47316));
    InMux I__11565 (
            .O(N__47335),
            .I(N__47312));
    LocalMux I__11564 (
            .O(N__47330),
            .I(N__47304));
    LocalMux I__11563 (
            .O(N__47327),
            .I(N__47301));
    InMux I__11562 (
            .O(N__47326),
            .I(N__47294));
    InMux I__11561 (
            .O(N__47325),
            .I(N__47294));
    InMux I__11560 (
            .O(N__47324),
            .I(N__47294));
    InMux I__11559 (
            .O(N__47323),
            .I(N__47285));
    InMux I__11558 (
            .O(N__47322),
            .I(N__47285));
    InMux I__11557 (
            .O(N__47321),
            .I(N__47278));
    InMux I__11556 (
            .O(N__47320),
            .I(N__47278));
    InMux I__11555 (
            .O(N__47319),
            .I(N__47278));
    InMux I__11554 (
            .O(N__47316),
            .I(N__47275));
    CascadeMux I__11553 (
            .O(N__47315),
            .I(N__47269));
    LocalMux I__11552 (
            .O(N__47312),
            .I(N__47263));
    InMux I__11551 (
            .O(N__47311),
            .I(N__47257));
    InMux I__11550 (
            .O(N__47310),
            .I(N__47240));
    CascadeMux I__11549 (
            .O(N__47309),
            .I(N__47233));
    InMux I__11548 (
            .O(N__47308),
            .I(N__47227));
    CascadeMux I__11547 (
            .O(N__47307),
            .I(N__47224));
    Span4Mux_h I__11546 (
            .O(N__47304),
            .I(N__47217));
    Span4Mux_v I__11545 (
            .O(N__47301),
            .I(N__47217));
    LocalMux I__11544 (
            .O(N__47294),
            .I(N__47217));
    InMux I__11543 (
            .O(N__47293),
            .I(N__47214));
    InMux I__11542 (
            .O(N__47292),
            .I(N__47209));
    InMux I__11541 (
            .O(N__47291),
            .I(N__47209));
    InMux I__11540 (
            .O(N__47290),
            .I(N__47206));
    LocalMux I__11539 (
            .O(N__47285),
            .I(N__47199));
    LocalMux I__11538 (
            .O(N__47278),
            .I(N__47199));
    LocalMux I__11537 (
            .O(N__47275),
            .I(N__47199));
    InMux I__11536 (
            .O(N__47274),
            .I(N__47196));
    InMux I__11535 (
            .O(N__47273),
            .I(N__47191));
    InMux I__11534 (
            .O(N__47272),
            .I(N__47191));
    InMux I__11533 (
            .O(N__47269),
            .I(N__47188));
    InMux I__11532 (
            .O(N__47268),
            .I(N__47185));
    InMux I__11531 (
            .O(N__47267),
            .I(N__47178));
    InMux I__11530 (
            .O(N__47266),
            .I(N__47175));
    Span4Mux_v I__11529 (
            .O(N__47263),
            .I(N__47170));
    InMux I__11528 (
            .O(N__47262),
            .I(N__47163));
    InMux I__11527 (
            .O(N__47261),
            .I(N__47163));
    InMux I__11526 (
            .O(N__47260),
            .I(N__47163));
    LocalMux I__11525 (
            .O(N__47257),
            .I(N__47160));
    InMux I__11524 (
            .O(N__47256),
            .I(N__47153));
    InMux I__11523 (
            .O(N__47255),
            .I(N__47153));
    InMux I__11522 (
            .O(N__47254),
            .I(N__47153));
    InMux I__11521 (
            .O(N__47253),
            .I(N__47143));
    InMux I__11520 (
            .O(N__47252),
            .I(N__47143));
    InMux I__11519 (
            .O(N__47251),
            .I(N__47143));
    InMux I__11518 (
            .O(N__47250),
            .I(N__47134));
    InMux I__11517 (
            .O(N__47249),
            .I(N__47127));
    InMux I__11516 (
            .O(N__47248),
            .I(N__47127));
    InMux I__11515 (
            .O(N__47247),
            .I(N__47127));
    InMux I__11514 (
            .O(N__47246),
            .I(N__47124));
    InMux I__11513 (
            .O(N__47245),
            .I(N__47121));
    InMux I__11512 (
            .O(N__47244),
            .I(N__47116));
    InMux I__11511 (
            .O(N__47243),
            .I(N__47116));
    LocalMux I__11510 (
            .O(N__47240),
            .I(N__47113));
    InMux I__11509 (
            .O(N__47239),
            .I(N__47110));
    InMux I__11508 (
            .O(N__47238),
            .I(N__47107));
    InMux I__11507 (
            .O(N__47237),
            .I(N__47102));
    InMux I__11506 (
            .O(N__47236),
            .I(N__47102));
    InMux I__11505 (
            .O(N__47233),
            .I(N__47099));
    CascadeMux I__11504 (
            .O(N__47232),
            .I(N__47096));
    InMux I__11503 (
            .O(N__47231),
            .I(N__47089));
    InMux I__11502 (
            .O(N__47230),
            .I(N__47089));
    LocalMux I__11501 (
            .O(N__47227),
            .I(N__47081));
    InMux I__11500 (
            .O(N__47224),
            .I(N__47078));
    Span4Mux_h I__11499 (
            .O(N__47217),
            .I(N__47072));
    LocalMux I__11498 (
            .O(N__47214),
            .I(N__47072));
    LocalMux I__11497 (
            .O(N__47209),
            .I(N__47065));
    LocalMux I__11496 (
            .O(N__47206),
            .I(N__47065));
    Span4Mux_v I__11495 (
            .O(N__47199),
            .I(N__47065));
    LocalMux I__11494 (
            .O(N__47196),
            .I(N__47060));
    LocalMux I__11493 (
            .O(N__47191),
            .I(N__47060));
    LocalMux I__11492 (
            .O(N__47188),
            .I(N__47055));
    LocalMux I__11491 (
            .O(N__47185),
            .I(N__47055));
    CascadeMux I__11490 (
            .O(N__47184),
            .I(N__47052));
    CascadeMux I__11489 (
            .O(N__47183),
            .I(N__47049));
    CascadeMux I__11488 (
            .O(N__47182),
            .I(N__47043));
    CascadeMux I__11487 (
            .O(N__47181),
            .I(N__47040));
    LocalMux I__11486 (
            .O(N__47178),
            .I(N__47037));
    LocalMux I__11485 (
            .O(N__47175),
            .I(N__47034));
    InMux I__11484 (
            .O(N__47174),
            .I(N__47031));
    InMux I__11483 (
            .O(N__47173),
            .I(N__47028));
    Span4Mux_v I__11482 (
            .O(N__47170),
            .I(N__47018));
    LocalMux I__11481 (
            .O(N__47163),
            .I(N__47018));
    Span4Mux_v I__11480 (
            .O(N__47160),
            .I(N__47018));
    LocalMux I__11479 (
            .O(N__47153),
            .I(N__47018));
    InMux I__11478 (
            .O(N__47152),
            .I(N__47011));
    InMux I__11477 (
            .O(N__47151),
            .I(N__47011));
    InMux I__11476 (
            .O(N__47150),
            .I(N__47011));
    LocalMux I__11475 (
            .O(N__47143),
            .I(N__47008));
    InMux I__11474 (
            .O(N__47142),
            .I(N__47001));
    InMux I__11473 (
            .O(N__47141),
            .I(N__47001));
    InMux I__11472 (
            .O(N__47140),
            .I(N__47001));
    InMux I__11471 (
            .O(N__47139),
            .I(N__46994));
    InMux I__11470 (
            .O(N__47138),
            .I(N__46994));
    InMux I__11469 (
            .O(N__47137),
            .I(N__46994));
    LocalMux I__11468 (
            .O(N__47134),
            .I(N__46977));
    LocalMux I__11467 (
            .O(N__47127),
            .I(N__46977));
    LocalMux I__11466 (
            .O(N__47124),
            .I(N__46977));
    LocalMux I__11465 (
            .O(N__47121),
            .I(N__46977));
    LocalMux I__11464 (
            .O(N__47116),
            .I(N__46977));
    Span4Mux_v I__11463 (
            .O(N__47113),
            .I(N__46977));
    LocalMux I__11462 (
            .O(N__47110),
            .I(N__46977));
    LocalMux I__11461 (
            .O(N__47107),
            .I(N__46977));
    LocalMux I__11460 (
            .O(N__47102),
            .I(N__46972));
    LocalMux I__11459 (
            .O(N__47099),
            .I(N__46972));
    InMux I__11458 (
            .O(N__47096),
            .I(N__46967));
    InMux I__11457 (
            .O(N__47095),
            .I(N__46967));
    InMux I__11456 (
            .O(N__47094),
            .I(N__46960));
    LocalMux I__11455 (
            .O(N__47089),
            .I(N__46957));
    InMux I__11454 (
            .O(N__47088),
            .I(N__46952));
    InMux I__11453 (
            .O(N__47087),
            .I(N__46952));
    InMux I__11452 (
            .O(N__47086),
            .I(N__46947));
    InMux I__11451 (
            .O(N__47085),
            .I(N__46947));
    InMux I__11450 (
            .O(N__47084),
            .I(N__46943));
    Span4Mux_v I__11449 (
            .O(N__47081),
            .I(N__46938));
    LocalMux I__11448 (
            .O(N__47078),
            .I(N__46938));
    InMux I__11447 (
            .O(N__47077),
            .I(N__46935));
    Span4Mux_h I__11446 (
            .O(N__47072),
            .I(N__46932));
    Span4Mux_h I__11445 (
            .O(N__47065),
            .I(N__46924));
    Span4Mux_v I__11444 (
            .O(N__47060),
            .I(N__46924));
    Span4Mux_v I__11443 (
            .O(N__47055),
            .I(N__46924));
    InMux I__11442 (
            .O(N__47052),
            .I(N__46917));
    InMux I__11441 (
            .O(N__47049),
            .I(N__46917));
    InMux I__11440 (
            .O(N__47048),
            .I(N__46917));
    InMux I__11439 (
            .O(N__47047),
            .I(N__46912));
    InMux I__11438 (
            .O(N__47046),
            .I(N__46912));
    InMux I__11437 (
            .O(N__47043),
            .I(N__46905));
    InMux I__11436 (
            .O(N__47040),
            .I(N__46902));
    Span4Mux_h I__11435 (
            .O(N__47037),
            .I(N__46899));
    Span4Mux_h I__11434 (
            .O(N__47034),
            .I(N__46891));
    LocalMux I__11433 (
            .O(N__47031),
            .I(N__46891));
    LocalMux I__11432 (
            .O(N__47028),
            .I(N__46891));
    InMux I__11431 (
            .O(N__47027),
            .I(N__46888));
    Span4Mux_h I__11430 (
            .O(N__47018),
            .I(N__46875));
    LocalMux I__11429 (
            .O(N__47011),
            .I(N__46875));
    Span4Mux_v I__11428 (
            .O(N__47008),
            .I(N__46875));
    LocalMux I__11427 (
            .O(N__47001),
            .I(N__46875));
    LocalMux I__11426 (
            .O(N__46994),
            .I(N__46875));
    Span4Mux_v I__11425 (
            .O(N__46977),
            .I(N__46875));
    Span4Mux_v I__11424 (
            .O(N__46972),
            .I(N__46870));
    LocalMux I__11423 (
            .O(N__46967),
            .I(N__46870));
    InMux I__11422 (
            .O(N__46966),
            .I(N__46867));
    InMux I__11421 (
            .O(N__46965),
            .I(N__46864));
    InMux I__11420 (
            .O(N__46964),
            .I(N__46861));
    InMux I__11419 (
            .O(N__46963),
            .I(N__46858));
    LocalMux I__11418 (
            .O(N__46960),
            .I(N__46855));
    Sp12to4 I__11417 (
            .O(N__46957),
            .I(N__46848));
    LocalMux I__11416 (
            .O(N__46952),
            .I(N__46848));
    LocalMux I__11415 (
            .O(N__46947),
            .I(N__46848));
    InMux I__11414 (
            .O(N__46946),
            .I(N__46845));
    LocalMux I__11413 (
            .O(N__46943),
            .I(N__46842));
    Sp12to4 I__11412 (
            .O(N__46938),
            .I(N__46839));
    LocalMux I__11411 (
            .O(N__46935),
            .I(N__46836));
    Span4Mux_h I__11410 (
            .O(N__46932),
            .I(N__46830));
    InMux I__11409 (
            .O(N__46931),
            .I(N__46827));
    Span4Mux_h I__11408 (
            .O(N__46924),
            .I(N__46820));
    LocalMux I__11407 (
            .O(N__46917),
            .I(N__46820));
    LocalMux I__11406 (
            .O(N__46912),
            .I(N__46820));
    InMux I__11405 (
            .O(N__46911),
            .I(N__46814));
    InMux I__11404 (
            .O(N__46910),
            .I(N__46811));
    InMux I__11403 (
            .O(N__46909),
            .I(N__46806));
    InMux I__11402 (
            .O(N__46908),
            .I(N__46806));
    LocalMux I__11401 (
            .O(N__46905),
            .I(N__46799));
    LocalMux I__11400 (
            .O(N__46902),
            .I(N__46799));
    Span4Mux_v I__11399 (
            .O(N__46899),
            .I(N__46799));
    InMux I__11398 (
            .O(N__46898),
            .I(N__46796));
    Span4Mux_v I__11397 (
            .O(N__46891),
            .I(N__46787));
    LocalMux I__11396 (
            .O(N__46888),
            .I(N__46787));
    Span4Mux_h I__11395 (
            .O(N__46875),
            .I(N__46787));
    Span4Mux_v I__11394 (
            .O(N__46870),
            .I(N__46787));
    LocalMux I__11393 (
            .O(N__46867),
            .I(N__46772));
    LocalMux I__11392 (
            .O(N__46864),
            .I(N__46772));
    LocalMux I__11391 (
            .O(N__46861),
            .I(N__46772));
    LocalMux I__11390 (
            .O(N__46858),
            .I(N__46772));
    Span12Mux_s10_h I__11389 (
            .O(N__46855),
            .I(N__46772));
    Span12Mux_h I__11388 (
            .O(N__46848),
            .I(N__46772));
    LocalMux I__11387 (
            .O(N__46845),
            .I(N__46772));
    Span12Mux_v I__11386 (
            .O(N__46842),
            .I(N__46765));
    Span12Mux_v I__11385 (
            .O(N__46839),
            .I(N__46765));
    Span12Mux_h I__11384 (
            .O(N__46836),
            .I(N__46765));
    InMux I__11383 (
            .O(N__46835),
            .I(N__46758));
    InMux I__11382 (
            .O(N__46834),
            .I(N__46758));
    InMux I__11381 (
            .O(N__46833),
            .I(N__46758));
    Span4Mux_v I__11380 (
            .O(N__46830),
            .I(N__46751));
    LocalMux I__11379 (
            .O(N__46827),
            .I(N__46751));
    Span4Mux_h I__11378 (
            .O(N__46820),
            .I(N__46751));
    InMux I__11377 (
            .O(N__46819),
            .I(N__46748));
    InMux I__11376 (
            .O(N__46818),
            .I(N__46743));
    InMux I__11375 (
            .O(N__46817),
            .I(N__46743));
    LocalMux I__11374 (
            .O(N__46814),
            .I(comm_cmd_3));
    LocalMux I__11373 (
            .O(N__46811),
            .I(comm_cmd_3));
    LocalMux I__11372 (
            .O(N__46806),
            .I(comm_cmd_3));
    Odrv4 I__11371 (
            .O(N__46799),
            .I(comm_cmd_3));
    LocalMux I__11370 (
            .O(N__46796),
            .I(comm_cmd_3));
    Odrv4 I__11369 (
            .O(N__46787),
            .I(comm_cmd_3));
    Odrv12 I__11368 (
            .O(N__46772),
            .I(comm_cmd_3));
    Odrv12 I__11367 (
            .O(N__46765),
            .I(comm_cmd_3));
    LocalMux I__11366 (
            .O(N__46758),
            .I(comm_cmd_3));
    Odrv4 I__11365 (
            .O(N__46751),
            .I(comm_cmd_3));
    LocalMux I__11364 (
            .O(N__46748),
            .I(comm_cmd_3));
    LocalMux I__11363 (
            .O(N__46743),
            .I(comm_cmd_3));
    InMux I__11362 (
            .O(N__46718),
            .I(N__46715));
    LocalMux I__11361 (
            .O(N__46715),
            .I(N__46712));
    Span12Mux_h I__11360 (
            .O(N__46712),
            .I(N__46709));
    Odrv12 I__11359 (
            .O(N__46709),
            .I(n4108));
    CascadeMux I__11358 (
            .O(N__46706),
            .I(N__46703));
    InMux I__11357 (
            .O(N__46703),
            .I(N__46700));
    LocalMux I__11356 (
            .O(N__46700),
            .I(N__46697));
    Span4Mux_v I__11355 (
            .O(N__46697),
            .I(N__46692));
    CascadeMux I__11354 (
            .O(N__46696),
            .I(N__46689));
    InMux I__11353 (
            .O(N__46695),
            .I(N__46686));
    Sp12to4 I__11352 (
            .O(N__46692),
            .I(N__46683));
    InMux I__11351 (
            .O(N__46689),
            .I(N__46680));
    LocalMux I__11350 (
            .O(N__46686),
            .I(N__46677));
    Span12Mux_h I__11349 (
            .O(N__46683),
            .I(N__46674));
    LocalMux I__11348 (
            .O(N__46680),
            .I(cmd_rdadctmp_10_adj_1066));
    Odrv4 I__11347 (
            .O(N__46677),
            .I(cmd_rdadctmp_10_adj_1066));
    Odrv12 I__11346 (
            .O(N__46674),
            .I(cmd_rdadctmp_10_adj_1066));
    InMux I__11345 (
            .O(N__46667),
            .I(N__46663));
    InMux I__11344 (
            .O(N__46666),
            .I(N__46660));
    LocalMux I__11343 (
            .O(N__46663),
            .I(buf_adcdata2_2));
    LocalMux I__11342 (
            .O(N__46660),
            .I(buf_adcdata2_2));
    SRMux I__11341 (
            .O(N__46655),
            .I(N__46652));
    LocalMux I__11340 (
            .O(N__46652),
            .I(N__46649));
    Span4Mux_h I__11339 (
            .O(N__46649),
            .I(N__46646));
    Span4Mux_v I__11338 (
            .O(N__46646),
            .I(N__46643));
    Odrv4 I__11337 (
            .O(N__46643),
            .I(\comm_spi.data_tx_7__N_808 ));
    InMux I__11336 (
            .O(N__46640),
            .I(N__46635));
    InMux I__11335 (
            .O(N__46639),
            .I(N__46630));
    InMux I__11334 (
            .O(N__46638),
            .I(N__46630));
    LocalMux I__11333 (
            .O(N__46635),
            .I(N__46627));
    LocalMux I__11332 (
            .O(N__46630),
            .I(N__46624));
    Span4Mux_v I__11331 (
            .O(N__46627),
            .I(N__46621));
    Span12Mux_h I__11330 (
            .O(N__46624),
            .I(N__46618));
    Span4Mux_v I__11329 (
            .O(N__46621),
            .I(N__46615));
    Odrv12 I__11328 (
            .O(N__46618),
            .I(comm_tx_buf_4));
    Odrv4 I__11327 (
            .O(N__46615),
            .I(comm_tx_buf_4));
    InMux I__11326 (
            .O(N__46610),
            .I(N__46588));
    InMux I__11325 (
            .O(N__46609),
            .I(N__46588));
    InMux I__11324 (
            .O(N__46608),
            .I(N__46588));
    InMux I__11323 (
            .O(N__46607),
            .I(N__46588));
    InMux I__11322 (
            .O(N__46606),
            .I(N__46588));
    InMux I__11321 (
            .O(N__46605),
            .I(N__46585));
    InMux I__11320 (
            .O(N__46604),
            .I(N__46571));
    InMux I__11319 (
            .O(N__46603),
            .I(N__46562));
    InMux I__11318 (
            .O(N__46602),
            .I(N__46562));
    InMux I__11317 (
            .O(N__46601),
            .I(N__46562));
    InMux I__11316 (
            .O(N__46600),
            .I(N__46562));
    InMux I__11315 (
            .O(N__46599),
            .I(N__46557));
    LocalMux I__11314 (
            .O(N__46588),
            .I(N__46550));
    LocalMux I__11313 (
            .O(N__46585),
            .I(N__46550));
    SRMux I__11312 (
            .O(N__46584),
            .I(N__46547));
    InMux I__11311 (
            .O(N__46583),
            .I(N__46540));
    InMux I__11310 (
            .O(N__46582),
            .I(N__46540));
    InMux I__11309 (
            .O(N__46581),
            .I(N__46540));
    SRMux I__11308 (
            .O(N__46580),
            .I(N__46537));
    InMux I__11307 (
            .O(N__46579),
            .I(N__46524));
    InMux I__11306 (
            .O(N__46578),
            .I(N__46524));
    InMux I__11305 (
            .O(N__46577),
            .I(N__46524));
    InMux I__11304 (
            .O(N__46576),
            .I(N__46524));
    InMux I__11303 (
            .O(N__46575),
            .I(N__46524));
    InMux I__11302 (
            .O(N__46574),
            .I(N__46524));
    LocalMux I__11301 (
            .O(N__46571),
            .I(N__46519));
    LocalMux I__11300 (
            .O(N__46562),
            .I(N__46519));
    InMux I__11299 (
            .O(N__46561),
            .I(N__46516));
    InMux I__11298 (
            .O(N__46560),
            .I(N__46513));
    LocalMux I__11297 (
            .O(N__46557),
            .I(N__46510));
    InMux I__11296 (
            .O(N__46556),
            .I(N__46507));
    SRMux I__11295 (
            .O(N__46555),
            .I(N__46504));
    Span4Mux_v I__11294 (
            .O(N__46550),
            .I(N__46498));
    LocalMux I__11293 (
            .O(N__46547),
            .I(N__46495));
    LocalMux I__11292 (
            .O(N__46540),
            .I(N__46490));
    LocalMux I__11291 (
            .O(N__46537),
            .I(N__46490));
    LocalMux I__11290 (
            .O(N__46524),
            .I(N__46487));
    Span4Mux_v I__11289 (
            .O(N__46519),
            .I(N__46484));
    LocalMux I__11288 (
            .O(N__46516),
            .I(N__46481));
    LocalMux I__11287 (
            .O(N__46513),
            .I(N__46478));
    Span4Mux_v I__11286 (
            .O(N__46510),
            .I(N__46471));
    LocalMux I__11285 (
            .O(N__46507),
            .I(N__46471));
    LocalMux I__11284 (
            .O(N__46504),
            .I(N__46471));
    InMux I__11283 (
            .O(N__46503),
            .I(N__46466));
    InMux I__11282 (
            .O(N__46502),
            .I(N__46457));
    InMux I__11281 (
            .O(N__46501),
            .I(N__46457));
    Span4Mux_h I__11280 (
            .O(N__46498),
            .I(N__46450));
    Span4Mux_v I__11279 (
            .O(N__46495),
            .I(N__46450));
    Span4Mux_v I__11278 (
            .O(N__46490),
            .I(N__46450));
    Span4Mux_v I__11277 (
            .O(N__46487),
            .I(N__46447));
    Span4Mux_h I__11276 (
            .O(N__46484),
            .I(N__46442));
    Span4Mux_v I__11275 (
            .O(N__46481),
            .I(N__46442));
    Span4Mux_v I__11274 (
            .O(N__46478),
            .I(N__46437));
    Span4Mux_h I__11273 (
            .O(N__46471),
            .I(N__46437));
    InMux I__11272 (
            .O(N__46470),
            .I(N__46434));
    InMux I__11271 (
            .O(N__46469),
            .I(N__46431));
    LocalMux I__11270 (
            .O(N__46466),
            .I(N__46428));
    InMux I__11269 (
            .O(N__46465),
            .I(N__46419));
    InMux I__11268 (
            .O(N__46464),
            .I(N__46419));
    InMux I__11267 (
            .O(N__46463),
            .I(N__46419));
    InMux I__11266 (
            .O(N__46462),
            .I(N__46419));
    LocalMux I__11265 (
            .O(N__46457),
            .I(N__46412));
    Span4Mux_h I__11264 (
            .O(N__46450),
            .I(N__46412));
    Span4Mux_h I__11263 (
            .O(N__46447),
            .I(N__46412));
    Odrv4 I__11262 (
            .O(N__46442),
            .I(comm_clear));
    Odrv4 I__11261 (
            .O(N__46437),
            .I(comm_clear));
    LocalMux I__11260 (
            .O(N__46434),
            .I(comm_clear));
    LocalMux I__11259 (
            .O(N__46431),
            .I(comm_clear));
    Odrv4 I__11258 (
            .O(N__46428),
            .I(comm_clear));
    LocalMux I__11257 (
            .O(N__46419),
            .I(comm_clear));
    Odrv4 I__11256 (
            .O(N__46412),
            .I(comm_clear));
    InMux I__11255 (
            .O(N__46397),
            .I(N__46393));
    InMux I__11254 (
            .O(N__46396),
            .I(N__46390));
    LocalMux I__11253 (
            .O(N__46393),
            .I(N__46387));
    LocalMux I__11252 (
            .O(N__46390),
            .I(N__46384));
    Span4Mux_h I__11251 (
            .O(N__46387),
            .I(N__46381));
    Span4Mux_h I__11250 (
            .O(N__46384),
            .I(N__46378));
    Span4Mux_h I__11249 (
            .O(N__46381),
            .I(N__46374));
    Span4Mux_h I__11248 (
            .O(N__46378),
            .I(N__46371));
    InMux I__11247 (
            .O(N__46377),
            .I(N__46368));
    Odrv4 I__11246 (
            .O(N__46374),
            .I(\comm_spi.n16899 ));
    Odrv4 I__11245 (
            .O(N__46371),
            .I(\comm_spi.n16899 ));
    LocalMux I__11244 (
            .O(N__46368),
            .I(\comm_spi.n16899 ));
    CascadeMux I__11243 (
            .O(N__46361),
            .I(N__46358));
    InMux I__11242 (
            .O(N__46358),
            .I(N__46354));
    CascadeMux I__11241 (
            .O(N__46357),
            .I(N__46350));
    LocalMux I__11240 (
            .O(N__46354),
            .I(N__46347));
    InMux I__11239 (
            .O(N__46353),
            .I(N__46344));
    InMux I__11238 (
            .O(N__46350),
            .I(N__46341));
    Span4Mux_v I__11237 (
            .O(N__46347),
            .I(N__46338));
    LocalMux I__11236 (
            .O(N__46344),
            .I(cmd_rdadctmp_29_adj_1047));
    LocalMux I__11235 (
            .O(N__46341),
            .I(cmd_rdadctmp_29_adj_1047));
    Odrv4 I__11234 (
            .O(N__46338),
            .I(cmd_rdadctmp_29_adj_1047));
    InMux I__11233 (
            .O(N__46331),
            .I(N__46328));
    LocalMux I__11232 (
            .O(N__46328),
            .I(N__46324));
    InMux I__11231 (
            .O(N__46327),
            .I(N__46321));
    Span4Mux_v I__11230 (
            .O(N__46324),
            .I(N__46318));
    LocalMux I__11229 (
            .O(N__46321),
            .I(buf_adcdata2_21));
    Odrv4 I__11228 (
            .O(N__46318),
            .I(buf_adcdata2_21));
    IoInMux I__11227 (
            .O(N__46313),
            .I(N__46310));
    LocalMux I__11226 (
            .O(N__46310),
            .I(N__46307));
    IoSpan4Mux I__11225 (
            .O(N__46307),
            .I(N__46304));
    IoSpan4Mux I__11224 (
            .O(N__46304),
            .I(N__46301));
    Span4Mux_s3_h I__11223 (
            .O(N__46301),
            .I(N__46298));
    Span4Mux_h I__11222 (
            .O(N__46298),
            .I(N__46295));
    Odrv4 I__11221 (
            .O(N__46295),
            .I(ICE_GPMI_0));
    CascadeMux I__11220 (
            .O(N__46292),
            .I(N__46289));
    InMux I__11219 (
            .O(N__46289),
            .I(N__46286));
    LocalMux I__11218 (
            .O(N__46286),
            .I(N__46282));
    CascadeMux I__11217 (
            .O(N__46285),
            .I(N__46279));
    Span4Mux_v I__11216 (
            .O(N__46282),
            .I(N__46276));
    InMux I__11215 (
            .O(N__46279),
            .I(N__46273));
    Span4Mux_h I__11214 (
            .O(N__46276),
            .I(N__46269));
    LocalMux I__11213 (
            .O(N__46273),
            .I(N__46266));
    InMux I__11212 (
            .O(N__46272),
            .I(N__46263));
    Odrv4 I__11211 (
            .O(N__46269),
            .I(cmd_rdadctmp_20));
    Odrv4 I__11210 (
            .O(N__46266),
            .I(cmd_rdadctmp_20));
    LocalMux I__11209 (
            .O(N__46263),
            .I(cmd_rdadctmp_20));
    InMux I__11208 (
            .O(N__46256),
            .I(N__46253));
    LocalMux I__11207 (
            .O(N__46253),
            .I(N__46249));
    InMux I__11206 (
            .O(N__46252),
            .I(N__46246));
    Span4Mux_h I__11205 (
            .O(N__46249),
            .I(N__46243));
    LocalMux I__11204 (
            .O(N__46246),
            .I(buf_adcdata1_12));
    Odrv4 I__11203 (
            .O(N__46243),
            .I(buf_adcdata1_12));
    CascadeMux I__11202 (
            .O(N__46238),
            .I(N__46235));
    InMux I__11201 (
            .O(N__46235),
            .I(N__46232));
    LocalMux I__11200 (
            .O(N__46232),
            .I(N__46229));
    Span12Mux_s11_v I__11199 (
            .O(N__46229),
            .I(N__46224));
    InMux I__11198 (
            .O(N__46228),
            .I(N__46221));
    CascadeMux I__11197 (
            .O(N__46227),
            .I(N__46218));
    Span12Mux_h I__11196 (
            .O(N__46224),
            .I(N__46215));
    LocalMux I__11195 (
            .O(N__46221),
            .I(N__46212));
    InMux I__11194 (
            .O(N__46218),
            .I(N__46209));
    Odrv12 I__11193 (
            .O(N__46215),
            .I(cmd_rdadctmp_17_adj_1059));
    Odrv12 I__11192 (
            .O(N__46212),
            .I(cmd_rdadctmp_17_adj_1059));
    LocalMux I__11191 (
            .O(N__46209),
            .I(cmd_rdadctmp_17_adj_1059));
    InMux I__11190 (
            .O(N__46202),
            .I(N__46199));
    LocalMux I__11189 (
            .O(N__46199),
            .I(N__46196));
    Span4Mux_v I__11188 (
            .O(N__46196),
            .I(N__46192));
    InMux I__11187 (
            .O(N__46195),
            .I(N__46189));
    Span4Mux_h I__11186 (
            .O(N__46192),
            .I(N__46186));
    LocalMux I__11185 (
            .O(N__46189),
            .I(buf_adcdata2_9));
    Odrv4 I__11184 (
            .O(N__46186),
            .I(buf_adcdata2_9));
    CascadeMux I__11183 (
            .O(N__46181),
            .I(N__46178));
    InMux I__11182 (
            .O(N__46178),
            .I(N__46174));
    InMux I__11181 (
            .O(N__46177),
            .I(N__46171));
    LocalMux I__11180 (
            .O(N__46174),
            .I(N__46168));
    LocalMux I__11179 (
            .O(N__46171),
            .I(N__46165));
    Span4Mux_v I__11178 (
            .O(N__46168),
            .I(N__46159));
    Span4Mux_h I__11177 (
            .O(N__46165),
            .I(N__46159));
    CascadeMux I__11176 (
            .O(N__46164),
            .I(N__46156));
    Span4Mux_h I__11175 (
            .O(N__46159),
            .I(N__46153));
    InMux I__11174 (
            .O(N__46156),
            .I(N__46150));
    Odrv4 I__11173 (
            .O(N__46153),
            .I(cmd_rdadctmp_19_adj_1057));
    LocalMux I__11172 (
            .O(N__46150),
            .I(cmd_rdadctmp_19_adj_1057));
    CascadeMux I__11171 (
            .O(N__46145),
            .I(N__46142));
    InMux I__11170 (
            .O(N__46142),
            .I(N__46138));
    CascadeMux I__11169 (
            .O(N__46141),
            .I(N__46134));
    LocalMux I__11168 (
            .O(N__46138),
            .I(N__46131));
    InMux I__11167 (
            .O(N__46137),
            .I(N__46126));
    InMux I__11166 (
            .O(N__46134),
            .I(N__46126));
    Odrv4 I__11165 (
            .O(N__46131),
            .I(cmd_rdadctmp_20_adj_1056));
    LocalMux I__11164 (
            .O(N__46126),
            .I(cmd_rdadctmp_20_adj_1056));
    CascadeMux I__11163 (
            .O(N__46121),
            .I(N__46112));
    CascadeMux I__11162 (
            .O(N__46120),
            .I(N__46109));
    InMux I__11161 (
            .O(N__46119),
            .I(N__46097));
    InMux I__11160 (
            .O(N__46118),
            .I(N__46097));
    InMux I__11159 (
            .O(N__46117),
            .I(N__46097));
    InMux I__11158 (
            .O(N__46116),
            .I(N__46097));
    InMux I__11157 (
            .O(N__46115),
            .I(N__46097));
    InMux I__11156 (
            .O(N__46112),
            .I(N__46090));
    InMux I__11155 (
            .O(N__46109),
            .I(N__46090));
    InMux I__11154 (
            .O(N__46108),
            .I(N__46090));
    LocalMux I__11153 (
            .O(N__46097),
            .I(N__46086));
    LocalMux I__11152 (
            .O(N__46090),
            .I(N__46083));
    InMux I__11151 (
            .O(N__46089),
            .I(N__46073));
    Span4Mux_v I__11150 (
            .O(N__46086),
            .I(N__46067));
    Span4Mux_v I__11149 (
            .O(N__46083),
            .I(N__46067));
    InMux I__11148 (
            .O(N__46082),
            .I(N__46064));
    InMux I__11147 (
            .O(N__46081),
            .I(N__46059));
    InMux I__11146 (
            .O(N__46080),
            .I(N__46053));
    InMux I__11145 (
            .O(N__46079),
            .I(N__46053));
    InMux I__11144 (
            .O(N__46078),
            .I(N__46046));
    InMux I__11143 (
            .O(N__46077),
            .I(N__46046));
    InMux I__11142 (
            .O(N__46076),
            .I(N__46046));
    LocalMux I__11141 (
            .O(N__46073),
            .I(N__46043));
    InMux I__11140 (
            .O(N__46072),
            .I(N__46040));
    Span4Mux_h I__11139 (
            .O(N__46067),
            .I(N__46034));
    LocalMux I__11138 (
            .O(N__46064),
            .I(N__46031));
    InMux I__11137 (
            .O(N__46063),
            .I(N__46028));
    InMux I__11136 (
            .O(N__46062),
            .I(N__46025));
    LocalMux I__11135 (
            .O(N__46059),
            .I(N__46022));
    InMux I__11134 (
            .O(N__46058),
            .I(N__46019));
    LocalMux I__11133 (
            .O(N__46053),
            .I(N__46014));
    LocalMux I__11132 (
            .O(N__46046),
            .I(N__46014));
    Span4Mux_v I__11131 (
            .O(N__46043),
            .I(N__46011));
    LocalMux I__11130 (
            .O(N__46040),
            .I(N__46008));
    InMux I__11129 (
            .O(N__46039),
            .I(N__46005));
    CascadeMux I__11128 (
            .O(N__46038),
            .I(N__45998));
    CascadeMux I__11127 (
            .O(N__46037),
            .I(N__45994));
    Sp12to4 I__11126 (
            .O(N__46034),
            .I(N__45986));
    Span12Mux_v I__11125 (
            .O(N__46031),
            .I(N__45986));
    LocalMux I__11124 (
            .O(N__46028),
            .I(N__45986));
    LocalMux I__11123 (
            .O(N__46025),
            .I(N__45983));
    Span4Mux_h I__11122 (
            .O(N__46022),
            .I(N__45978));
    LocalMux I__11121 (
            .O(N__46019),
            .I(N__45978));
    Span4Mux_v I__11120 (
            .O(N__46014),
            .I(N__45975));
    Span4Mux_h I__11119 (
            .O(N__46011),
            .I(N__45968));
    Span4Mux_v I__11118 (
            .O(N__46008),
            .I(N__45968));
    LocalMux I__11117 (
            .O(N__46005),
            .I(N__45968));
    InMux I__11116 (
            .O(N__46004),
            .I(N__45959));
    InMux I__11115 (
            .O(N__46003),
            .I(N__45959));
    InMux I__11114 (
            .O(N__46002),
            .I(N__45959));
    InMux I__11113 (
            .O(N__46001),
            .I(N__45959));
    InMux I__11112 (
            .O(N__45998),
            .I(N__45950));
    InMux I__11111 (
            .O(N__45997),
            .I(N__45950));
    InMux I__11110 (
            .O(N__45994),
            .I(N__45950));
    InMux I__11109 (
            .O(N__45993),
            .I(N__45950));
    Span12Mux_h I__11108 (
            .O(N__45986),
            .I(N__45945));
    Span4Mux_v I__11107 (
            .O(N__45983),
            .I(N__45942));
    Span4Mux_h I__11106 (
            .O(N__45978),
            .I(N__45939));
    Span4Mux_v I__11105 (
            .O(N__45975),
            .I(N__45934));
    Span4Mux_h I__11104 (
            .O(N__45968),
            .I(N__45934));
    LocalMux I__11103 (
            .O(N__45959),
            .I(N__45931));
    LocalMux I__11102 (
            .O(N__45950),
            .I(N__45928));
    InMux I__11101 (
            .O(N__45949),
            .I(N__45923));
    InMux I__11100 (
            .O(N__45948),
            .I(N__45923));
    Odrv12 I__11099 (
            .O(N__45945),
            .I(n8302));
    Odrv4 I__11098 (
            .O(N__45942),
            .I(n8302));
    Odrv4 I__11097 (
            .O(N__45939),
            .I(n8302));
    Odrv4 I__11096 (
            .O(N__45934),
            .I(n8302));
    Odrv12 I__11095 (
            .O(N__45931),
            .I(n8302));
    Odrv4 I__11094 (
            .O(N__45928),
            .I(n8302));
    LocalMux I__11093 (
            .O(N__45923),
            .I(n8302));
    CascadeMux I__11092 (
            .O(N__45908),
            .I(N__45905));
    InMux I__11091 (
            .O(N__45905),
            .I(N__45900));
    InMux I__11090 (
            .O(N__45904),
            .I(N__45895));
    InMux I__11089 (
            .O(N__45903),
            .I(N__45895));
    LocalMux I__11088 (
            .O(N__45900),
            .I(cmd_rdadctmp_21_adj_1055));
    LocalMux I__11087 (
            .O(N__45895),
            .I(cmd_rdadctmp_21_adj_1055));
    InMux I__11086 (
            .O(N__45890),
            .I(N__45887));
    LocalMux I__11085 (
            .O(N__45887),
            .I(N__45884));
    Span4Mux_h I__11084 (
            .O(N__45884),
            .I(N__45881));
    Odrv4 I__11083 (
            .O(N__45881),
            .I(buf_data2_23));
    InMux I__11082 (
            .O(N__45878),
            .I(N__45874));
    CascadeMux I__11081 (
            .O(N__45877),
            .I(N__45871));
    LocalMux I__11080 (
            .O(N__45874),
            .I(N__45868));
    InMux I__11079 (
            .O(N__45871),
            .I(N__45864));
    Span4Mux_h I__11078 (
            .O(N__45868),
            .I(N__45861));
    CascadeMux I__11077 (
            .O(N__45867),
            .I(N__45858));
    LocalMux I__11076 (
            .O(N__45864),
            .I(N__45855));
    Span4Mux_v I__11075 (
            .O(N__45861),
            .I(N__45852));
    InMux I__11074 (
            .O(N__45858),
            .I(N__45849));
    Span12Mux_s10_v I__11073 (
            .O(N__45855),
            .I(N__45846));
    Span4Mux_h I__11072 (
            .O(N__45852),
            .I(N__45843));
    LocalMux I__11071 (
            .O(N__45849),
            .I(buf_adcdata4_23));
    Odrv12 I__11070 (
            .O(N__45846),
            .I(buf_adcdata4_23));
    Odrv4 I__11069 (
            .O(N__45843),
            .I(buf_adcdata4_23));
    InMux I__11068 (
            .O(N__45836),
            .I(N__45833));
    LocalMux I__11067 (
            .O(N__45833),
            .I(N__45830));
    Span4Mux_v I__11066 (
            .O(N__45830),
            .I(N__45827));
    Span4Mux_h I__11065 (
            .O(N__45827),
            .I(N__45824));
    Sp12to4 I__11064 (
            .O(N__45824),
            .I(N__45821));
    Odrv12 I__11063 (
            .O(N__45821),
            .I(n4101));
    InMux I__11062 (
            .O(N__45818),
            .I(N__45815));
    LocalMux I__11061 (
            .O(N__45815),
            .I(N__45810));
    InMux I__11060 (
            .O(N__45814),
            .I(N__45807));
    InMux I__11059 (
            .O(N__45813),
            .I(N__45804));
    Odrv12 I__11058 (
            .O(N__45810),
            .I(\comm_spi.n10442 ));
    LocalMux I__11057 (
            .O(N__45807),
            .I(\comm_spi.n10442 ));
    LocalMux I__11056 (
            .O(N__45804),
            .I(\comm_spi.n10442 ));
    InMux I__11055 (
            .O(N__45797),
            .I(N__45789));
    InMux I__11054 (
            .O(N__45796),
            .I(N__45789));
    InMux I__11053 (
            .O(N__45795),
            .I(N__45786));
    InMux I__11052 (
            .O(N__45794),
            .I(N__45783));
    LocalMux I__11051 (
            .O(N__45789),
            .I(N__45778));
    LocalMux I__11050 (
            .O(N__45786),
            .I(N__45778));
    LocalMux I__11049 (
            .O(N__45783),
            .I(N__45774));
    Span4Mux_v I__11048 (
            .O(N__45778),
            .I(N__45771));
    InMux I__11047 (
            .O(N__45777),
            .I(N__45768));
    Span4Mux_v I__11046 (
            .O(N__45774),
            .I(N__45765));
    Span4Mux_h I__11045 (
            .O(N__45771),
            .I(N__45762));
    LocalMux I__11044 (
            .O(N__45768),
            .I(N__45759));
    Sp12to4 I__11043 (
            .O(N__45765),
            .I(N__45754));
    Sp12to4 I__11042 (
            .O(N__45762),
            .I(N__45754));
    Span4Mux_h I__11041 (
            .O(N__45759),
            .I(N__45751));
    Span12Mux_s6_h I__11040 (
            .O(N__45754),
            .I(N__45746));
    Sp12to4 I__11039 (
            .O(N__45751),
            .I(N__45746));
    Span12Mux_v I__11038 (
            .O(N__45746),
            .I(N__45743));
    Odrv12 I__11037 (
            .O(N__45743),
            .I(ICE_SPI_MOSI));
    SRMux I__11036 (
            .O(N__45740),
            .I(N__45737));
    LocalMux I__11035 (
            .O(N__45737),
            .I(\comm_spi.imosi_N_792 ));
    CascadeMux I__11034 (
            .O(N__45734),
            .I(N__45731));
    InMux I__11033 (
            .O(N__45731),
            .I(N__45727));
    CascadeMux I__11032 (
            .O(N__45730),
            .I(N__45723));
    LocalMux I__11031 (
            .O(N__45727),
            .I(N__45720));
    InMux I__11030 (
            .O(N__45726),
            .I(N__45715));
    InMux I__11029 (
            .O(N__45723),
            .I(N__45715));
    Span4Mux_v I__11028 (
            .O(N__45720),
            .I(N__45712));
    LocalMux I__11027 (
            .O(N__45715),
            .I(cmd_rdadctmp_28_adj_1048));
    Odrv4 I__11026 (
            .O(N__45712),
            .I(cmd_rdadctmp_28_adj_1048));
    InMux I__11025 (
            .O(N__45707),
            .I(N__45704));
    LocalMux I__11024 (
            .O(N__45704),
            .I(N__45700));
    InMux I__11023 (
            .O(N__45703),
            .I(N__45697));
    Span4Mux_h I__11022 (
            .O(N__45700),
            .I(N__45694));
    LocalMux I__11021 (
            .O(N__45697),
            .I(buf_adcdata2_20));
    Odrv4 I__11020 (
            .O(N__45694),
            .I(buf_adcdata2_20));
    InMux I__11019 (
            .O(N__45689),
            .I(N__45686));
    LocalMux I__11018 (
            .O(N__45686),
            .I(N__45683));
    Odrv12 I__11017 (
            .O(N__45683),
            .I(n4_adj_1250));
    InMux I__11016 (
            .O(N__45680),
            .I(N__45677));
    LocalMux I__11015 (
            .O(N__45677),
            .I(N__45673));
    InMux I__11014 (
            .O(N__45676),
            .I(N__45670));
    Span4Mux_h I__11013 (
            .O(N__45673),
            .I(N__45667));
    LocalMux I__11012 (
            .O(N__45670),
            .I(buf_adcdata2_12));
    Odrv4 I__11011 (
            .O(N__45667),
            .I(buf_adcdata2_12));
    InMux I__11010 (
            .O(N__45662),
            .I(N__45640));
    InMux I__11009 (
            .O(N__45661),
            .I(N__45640));
    InMux I__11008 (
            .O(N__45660),
            .I(N__45636));
    InMux I__11007 (
            .O(N__45659),
            .I(N__45633));
    InMux I__11006 (
            .O(N__45658),
            .I(N__45630));
    InMux I__11005 (
            .O(N__45657),
            .I(N__45627));
    InMux I__11004 (
            .O(N__45656),
            .I(N__45622));
    InMux I__11003 (
            .O(N__45655),
            .I(N__45622));
    InMux I__11002 (
            .O(N__45654),
            .I(N__45619));
    CascadeMux I__11001 (
            .O(N__45653),
            .I(N__45616));
    InMux I__11000 (
            .O(N__45652),
            .I(N__45613));
    InMux I__10999 (
            .O(N__45651),
            .I(N__45608));
    InMux I__10998 (
            .O(N__45650),
            .I(N__45608));
    InMux I__10997 (
            .O(N__45649),
            .I(N__45599));
    InMux I__10996 (
            .O(N__45648),
            .I(N__45592));
    InMux I__10995 (
            .O(N__45647),
            .I(N__45592));
    InMux I__10994 (
            .O(N__45646),
            .I(N__45589));
    InMux I__10993 (
            .O(N__45645),
            .I(N__45586));
    LocalMux I__10992 (
            .O(N__45640),
            .I(N__45583));
    InMux I__10991 (
            .O(N__45639),
            .I(N__45580));
    LocalMux I__10990 (
            .O(N__45636),
            .I(N__45575));
    LocalMux I__10989 (
            .O(N__45633),
            .I(N__45575));
    LocalMux I__10988 (
            .O(N__45630),
            .I(N__45572));
    LocalMux I__10987 (
            .O(N__45627),
            .I(N__45569));
    LocalMux I__10986 (
            .O(N__45622),
            .I(N__45566));
    LocalMux I__10985 (
            .O(N__45619),
            .I(N__45563));
    InMux I__10984 (
            .O(N__45616),
            .I(N__45560));
    LocalMux I__10983 (
            .O(N__45613),
            .I(N__45557));
    LocalMux I__10982 (
            .O(N__45608),
            .I(N__45554));
    InMux I__10981 (
            .O(N__45607),
            .I(N__45551));
    InMux I__10980 (
            .O(N__45606),
            .I(N__45546));
    InMux I__10979 (
            .O(N__45605),
            .I(N__45546));
    InMux I__10978 (
            .O(N__45604),
            .I(N__45531));
    InMux I__10977 (
            .O(N__45603),
            .I(N__45531));
    InMux I__10976 (
            .O(N__45602),
            .I(N__45528));
    LocalMux I__10975 (
            .O(N__45599),
            .I(N__45525));
    InMux I__10974 (
            .O(N__45598),
            .I(N__45522));
    InMux I__10973 (
            .O(N__45597),
            .I(N__45519));
    LocalMux I__10972 (
            .O(N__45592),
            .I(N__45506));
    LocalMux I__10971 (
            .O(N__45589),
            .I(N__45506));
    LocalMux I__10970 (
            .O(N__45586),
            .I(N__45506));
    Span4Mux_v I__10969 (
            .O(N__45583),
            .I(N__45506));
    LocalMux I__10968 (
            .O(N__45580),
            .I(N__45506));
    Span4Mux_h I__10967 (
            .O(N__45575),
            .I(N__45506));
    Span4Mux_v I__10966 (
            .O(N__45572),
            .I(N__45501));
    Span4Mux_v I__10965 (
            .O(N__45569),
            .I(N__45501));
    Span4Mux_h I__10964 (
            .O(N__45566),
            .I(N__45497));
    Span4Mux_h I__10963 (
            .O(N__45563),
            .I(N__45488));
    LocalMux I__10962 (
            .O(N__45560),
            .I(N__45488));
    Span4Mux_v I__10961 (
            .O(N__45557),
            .I(N__45488));
    Span4Mux_v I__10960 (
            .O(N__45554),
            .I(N__45488));
    LocalMux I__10959 (
            .O(N__45551),
            .I(N__45483));
    LocalMux I__10958 (
            .O(N__45546),
            .I(N__45483));
    InMux I__10957 (
            .O(N__45545),
            .I(N__45478));
    InMux I__10956 (
            .O(N__45544),
            .I(N__45478));
    InMux I__10955 (
            .O(N__45543),
            .I(N__45471));
    InMux I__10954 (
            .O(N__45542),
            .I(N__45471));
    InMux I__10953 (
            .O(N__45541),
            .I(N__45471));
    InMux I__10952 (
            .O(N__45540),
            .I(N__45466));
    InMux I__10951 (
            .O(N__45539),
            .I(N__45466));
    InMux I__10950 (
            .O(N__45538),
            .I(N__45461));
    InMux I__10949 (
            .O(N__45537),
            .I(N__45456));
    InMux I__10948 (
            .O(N__45536),
            .I(N__45456));
    LocalMux I__10947 (
            .O(N__45531),
            .I(N__45451));
    LocalMux I__10946 (
            .O(N__45528),
            .I(N__45446));
    Span4Mux_h I__10945 (
            .O(N__45525),
            .I(N__45446));
    LocalMux I__10944 (
            .O(N__45522),
            .I(N__45441));
    LocalMux I__10943 (
            .O(N__45519),
            .I(N__45441));
    Span4Mux_h I__10942 (
            .O(N__45506),
            .I(N__45438));
    Span4Mux_h I__10941 (
            .O(N__45501),
            .I(N__45432));
    InMux I__10940 (
            .O(N__45500),
            .I(N__45429));
    Span4Mux_h I__10939 (
            .O(N__45497),
            .I(N__45416));
    Span4Mux_h I__10938 (
            .O(N__45488),
            .I(N__45416));
    Span4Mux_v I__10937 (
            .O(N__45483),
            .I(N__45416));
    LocalMux I__10936 (
            .O(N__45478),
            .I(N__45416));
    LocalMux I__10935 (
            .O(N__45471),
            .I(N__45416));
    LocalMux I__10934 (
            .O(N__45466),
            .I(N__45416));
    CascadeMux I__10933 (
            .O(N__45465),
            .I(N__45406));
    InMux I__10932 (
            .O(N__45464),
            .I(N__45402));
    LocalMux I__10931 (
            .O(N__45461),
            .I(N__45397));
    LocalMux I__10930 (
            .O(N__45456),
            .I(N__45397));
    InMux I__10929 (
            .O(N__45455),
            .I(N__45394));
    InMux I__10928 (
            .O(N__45454),
            .I(N__45391));
    Span4Mux_h I__10927 (
            .O(N__45451),
            .I(N__45382));
    Span4Mux_v I__10926 (
            .O(N__45446),
            .I(N__45382));
    Span4Mux_h I__10925 (
            .O(N__45441),
            .I(N__45382));
    Span4Mux_h I__10924 (
            .O(N__45438),
            .I(N__45382));
    InMux I__10923 (
            .O(N__45437),
            .I(N__45379));
    InMux I__10922 (
            .O(N__45436),
            .I(N__45374));
    InMux I__10921 (
            .O(N__45435),
            .I(N__45374));
    Span4Mux_h I__10920 (
            .O(N__45432),
            .I(N__45369));
    LocalMux I__10919 (
            .O(N__45429),
            .I(N__45369));
    Span4Mux_v I__10918 (
            .O(N__45416),
            .I(N__45366));
    InMux I__10917 (
            .O(N__45415),
            .I(N__45361));
    InMux I__10916 (
            .O(N__45414),
            .I(N__45361));
    InMux I__10915 (
            .O(N__45413),
            .I(N__45352));
    InMux I__10914 (
            .O(N__45412),
            .I(N__45352));
    InMux I__10913 (
            .O(N__45411),
            .I(N__45352));
    InMux I__10912 (
            .O(N__45410),
            .I(N__45352));
    InMux I__10911 (
            .O(N__45409),
            .I(N__45349));
    InMux I__10910 (
            .O(N__45406),
            .I(N__45344));
    InMux I__10909 (
            .O(N__45405),
            .I(N__45344));
    LocalMux I__10908 (
            .O(N__45402),
            .I(comm_cmd_2));
    Odrv12 I__10907 (
            .O(N__45397),
            .I(comm_cmd_2));
    LocalMux I__10906 (
            .O(N__45394),
            .I(comm_cmd_2));
    LocalMux I__10905 (
            .O(N__45391),
            .I(comm_cmd_2));
    Odrv4 I__10904 (
            .O(N__45382),
            .I(comm_cmd_2));
    LocalMux I__10903 (
            .O(N__45379),
            .I(comm_cmd_2));
    LocalMux I__10902 (
            .O(N__45374),
            .I(comm_cmd_2));
    Odrv4 I__10901 (
            .O(N__45369),
            .I(comm_cmd_2));
    Odrv4 I__10900 (
            .O(N__45366),
            .I(comm_cmd_2));
    LocalMux I__10899 (
            .O(N__45361),
            .I(comm_cmd_2));
    LocalMux I__10898 (
            .O(N__45352),
            .I(comm_cmd_2));
    LocalMux I__10897 (
            .O(N__45349),
            .I(comm_cmd_2));
    LocalMux I__10896 (
            .O(N__45344),
            .I(comm_cmd_2));
    CascadeMux I__10895 (
            .O(N__45317),
            .I(N__45314));
    InMux I__10894 (
            .O(N__45314),
            .I(N__45310));
    CascadeMux I__10893 (
            .O(N__45313),
            .I(N__45303));
    LocalMux I__10892 (
            .O(N__45310),
            .I(N__45299));
    InMux I__10891 (
            .O(N__45309),
            .I(N__45290));
    InMux I__10890 (
            .O(N__45308),
            .I(N__45286));
    InMux I__10889 (
            .O(N__45307),
            .I(N__45280));
    InMux I__10888 (
            .O(N__45306),
            .I(N__45280));
    InMux I__10887 (
            .O(N__45303),
            .I(N__45273));
    InMux I__10886 (
            .O(N__45302),
            .I(N__45273));
    Span4Mux_v I__10885 (
            .O(N__45299),
            .I(N__45270));
    InMux I__10884 (
            .O(N__45298),
            .I(N__45265));
    InMux I__10883 (
            .O(N__45297),
            .I(N__45265));
    InMux I__10882 (
            .O(N__45296),
            .I(N__45256));
    InMux I__10881 (
            .O(N__45295),
            .I(N__45256));
    InMux I__10880 (
            .O(N__45294),
            .I(N__45253));
    InMux I__10879 (
            .O(N__45293),
            .I(N__45250));
    LocalMux I__10878 (
            .O(N__45290),
            .I(N__45247));
    InMux I__10877 (
            .O(N__45289),
            .I(N__45244));
    LocalMux I__10876 (
            .O(N__45286),
            .I(N__45241));
    InMux I__10875 (
            .O(N__45285),
            .I(N__45226));
    LocalMux I__10874 (
            .O(N__45280),
            .I(N__45212));
    InMux I__10873 (
            .O(N__45279),
            .I(N__45207));
    InMux I__10872 (
            .O(N__45278),
            .I(N__45207));
    LocalMux I__10871 (
            .O(N__45273),
            .I(N__45200));
    Span4Mux_h I__10870 (
            .O(N__45270),
            .I(N__45200));
    LocalMux I__10869 (
            .O(N__45265),
            .I(N__45200));
    InMux I__10868 (
            .O(N__45264),
            .I(N__45197));
    InMux I__10867 (
            .O(N__45263),
            .I(N__45190));
    InMux I__10866 (
            .O(N__45262),
            .I(N__45190));
    InMux I__10865 (
            .O(N__45261),
            .I(N__45190));
    LocalMux I__10864 (
            .O(N__45256),
            .I(N__45185));
    LocalMux I__10863 (
            .O(N__45253),
            .I(N__45185));
    LocalMux I__10862 (
            .O(N__45250),
            .I(N__45173));
    Span4Mux_h I__10861 (
            .O(N__45247),
            .I(N__45173));
    LocalMux I__10860 (
            .O(N__45244),
            .I(N__45173));
    Span4Mux_v I__10859 (
            .O(N__45241),
            .I(N__45173));
    InMux I__10858 (
            .O(N__45240),
            .I(N__45170));
    InMux I__10857 (
            .O(N__45239),
            .I(N__45167));
    InMux I__10856 (
            .O(N__45238),
            .I(N__45160));
    InMux I__10855 (
            .O(N__45237),
            .I(N__45160));
    InMux I__10854 (
            .O(N__45236),
            .I(N__45160));
    InMux I__10853 (
            .O(N__45235),
            .I(N__45155));
    InMux I__10852 (
            .O(N__45234),
            .I(N__45155));
    InMux I__10851 (
            .O(N__45233),
            .I(N__45142));
    InMux I__10850 (
            .O(N__45232),
            .I(N__45142));
    InMux I__10849 (
            .O(N__45231),
            .I(N__45142));
    InMux I__10848 (
            .O(N__45230),
            .I(N__45142));
    InMux I__10847 (
            .O(N__45229),
            .I(N__45139));
    LocalMux I__10846 (
            .O(N__45226),
            .I(N__45136));
    InMux I__10845 (
            .O(N__45225),
            .I(N__45133));
    InMux I__10844 (
            .O(N__45224),
            .I(N__45128));
    InMux I__10843 (
            .O(N__45223),
            .I(N__45128));
    InMux I__10842 (
            .O(N__45222),
            .I(N__45123));
    InMux I__10841 (
            .O(N__45221),
            .I(N__45123));
    InMux I__10840 (
            .O(N__45220),
            .I(N__45120));
    InMux I__10839 (
            .O(N__45219),
            .I(N__45117));
    InMux I__10838 (
            .O(N__45218),
            .I(N__45114));
    InMux I__10837 (
            .O(N__45217),
            .I(N__45109));
    InMux I__10836 (
            .O(N__45216),
            .I(N__45109));
    CascadeMux I__10835 (
            .O(N__45215),
            .I(N__45106));
    Span4Mux_h I__10834 (
            .O(N__45212),
            .I(N__45096));
    LocalMux I__10833 (
            .O(N__45207),
            .I(N__45096));
    Span4Mux_h I__10832 (
            .O(N__45200),
            .I(N__45096));
    LocalMux I__10831 (
            .O(N__45197),
            .I(N__45096));
    LocalMux I__10830 (
            .O(N__45190),
            .I(N__45091));
    Span4Mux_h I__10829 (
            .O(N__45185),
            .I(N__45091));
    InMux I__10828 (
            .O(N__45184),
            .I(N__45084));
    InMux I__10827 (
            .O(N__45183),
            .I(N__45084));
    InMux I__10826 (
            .O(N__45182),
            .I(N__45084));
    Span4Mux_h I__10825 (
            .O(N__45173),
            .I(N__45079));
    LocalMux I__10824 (
            .O(N__45170),
            .I(N__45079));
    LocalMux I__10823 (
            .O(N__45167),
            .I(N__45076));
    LocalMux I__10822 (
            .O(N__45160),
            .I(N__45071));
    LocalMux I__10821 (
            .O(N__45155),
            .I(N__45071));
    InMux I__10820 (
            .O(N__45154),
            .I(N__45066));
    InMux I__10819 (
            .O(N__45153),
            .I(N__45066));
    InMux I__10818 (
            .O(N__45152),
            .I(N__45063));
    InMux I__10817 (
            .O(N__45151),
            .I(N__45060));
    LocalMux I__10816 (
            .O(N__45142),
            .I(N__45055));
    LocalMux I__10815 (
            .O(N__45139),
            .I(N__45044));
    Span4Mux_v I__10814 (
            .O(N__45136),
            .I(N__45044));
    LocalMux I__10813 (
            .O(N__45133),
            .I(N__45044));
    LocalMux I__10812 (
            .O(N__45128),
            .I(N__45044));
    LocalMux I__10811 (
            .O(N__45123),
            .I(N__45044));
    LocalMux I__10810 (
            .O(N__45120),
            .I(N__45031));
    LocalMux I__10809 (
            .O(N__45117),
            .I(N__45031));
    LocalMux I__10808 (
            .O(N__45114),
            .I(N__45031));
    LocalMux I__10807 (
            .O(N__45109),
            .I(N__45031));
    InMux I__10806 (
            .O(N__45106),
            .I(N__45026));
    InMux I__10805 (
            .O(N__45105),
            .I(N__45026));
    Span4Mux_v I__10804 (
            .O(N__45096),
            .I(N__45019));
    Span4Mux_v I__10803 (
            .O(N__45091),
            .I(N__45019));
    LocalMux I__10802 (
            .O(N__45084),
            .I(N__45019));
    Span4Mux_h I__10801 (
            .O(N__45079),
            .I(N__45006));
    Span4Mux_h I__10800 (
            .O(N__45076),
            .I(N__45006));
    Span4Mux_v I__10799 (
            .O(N__45071),
            .I(N__45006));
    LocalMux I__10798 (
            .O(N__45066),
            .I(N__45006));
    LocalMux I__10797 (
            .O(N__45063),
            .I(N__45006));
    LocalMux I__10796 (
            .O(N__45060),
            .I(N__45006));
    InMux I__10795 (
            .O(N__45059),
            .I(N__45001));
    InMux I__10794 (
            .O(N__45058),
            .I(N__45001));
    Span4Mux_h I__10793 (
            .O(N__45055),
            .I(N__44996));
    Span4Mux_h I__10792 (
            .O(N__45044),
            .I(N__44996));
    InMux I__10791 (
            .O(N__45043),
            .I(N__44991));
    InMux I__10790 (
            .O(N__45042),
            .I(N__44991));
    InMux I__10789 (
            .O(N__45041),
            .I(N__44986));
    InMux I__10788 (
            .O(N__45040),
            .I(N__44986));
    Odrv12 I__10787 (
            .O(N__45031),
            .I(comm_cmd_1));
    LocalMux I__10786 (
            .O(N__45026),
            .I(comm_cmd_1));
    Odrv4 I__10785 (
            .O(N__45019),
            .I(comm_cmd_1));
    Odrv4 I__10784 (
            .O(N__45006),
            .I(comm_cmd_1));
    LocalMux I__10783 (
            .O(N__45001),
            .I(comm_cmd_1));
    Odrv4 I__10782 (
            .O(N__44996),
            .I(comm_cmd_1));
    LocalMux I__10781 (
            .O(N__44991),
            .I(comm_cmd_1));
    LocalMux I__10780 (
            .O(N__44986),
            .I(comm_cmd_1));
    InMux I__10779 (
            .O(N__44969),
            .I(N__44964));
    InMux I__10778 (
            .O(N__44968),
            .I(N__44960));
    InMux I__10777 (
            .O(N__44967),
            .I(N__44957));
    LocalMux I__10776 (
            .O(N__44964),
            .I(N__44954));
    InMux I__10775 (
            .O(N__44963),
            .I(N__44951));
    LocalMux I__10774 (
            .O(N__44960),
            .I(N__44948));
    LocalMux I__10773 (
            .O(N__44957),
            .I(N__44945));
    Span4Mux_h I__10772 (
            .O(N__44954),
            .I(N__44942));
    LocalMux I__10771 (
            .O(N__44951),
            .I(N__44939));
    Span4Mux_h I__10770 (
            .O(N__44948),
            .I(N__44934));
    Span4Mux_h I__10769 (
            .O(N__44945),
            .I(N__44934));
    Span4Mux_v I__10768 (
            .O(N__44942),
            .I(N__44931));
    Span4Mux_h I__10767 (
            .O(N__44939),
            .I(N__44926));
    Span4Mux_v I__10766 (
            .O(N__44934),
            .I(N__44926));
    Odrv4 I__10765 (
            .O(N__44931),
            .I(n9));
    Odrv4 I__10764 (
            .O(N__44926),
            .I(n9));
    InMux I__10763 (
            .O(N__44921),
            .I(N__44918));
    LocalMux I__10762 (
            .O(N__44918),
            .I(N__44914));
    InMux I__10761 (
            .O(N__44917),
            .I(N__44911));
    Span4Mux_v I__10760 (
            .O(N__44914),
            .I(N__44904));
    LocalMux I__10759 (
            .O(N__44911),
            .I(N__44901));
    InMux I__10758 (
            .O(N__44910),
            .I(N__44898));
    InMux I__10757 (
            .O(N__44909),
            .I(N__44895));
    InMux I__10756 (
            .O(N__44908),
            .I(N__44892));
    InMux I__10755 (
            .O(N__44907),
            .I(N__44889));
    Span4Mux_h I__10754 (
            .O(N__44904),
            .I(N__44874));
    Span4Mux_v I__10753 (
            .O(N__44901),
            .I(N__44874));
    LocalMux I__10752 (
            .O(N__44898),
            .I(N__44874));
    LocalMux I__10751 (
            .O(N__44895),
            .I(N__44874));
    LocalMux I__10750 (
            .O(N__44892),
            .I(N__44869));
    LocalMux I__10749 (
            .O(N__44889),
            .I(N__44869));
    InMux I__10748 (
            .O(N__44888),
            .I(N__44866));
    InMux I__10747 (
            .O(N__44887),
            .I(N__44863));
    InMux I__10746 (
            .O(N__44886),
            .I(N__44860));
    InMux I__10745 (
            .O(N__44885),
            .I(N__44857));
    InMux I__10744 (
            .O(N__44884),
            .I(N__44853));
    CascadeMux I__10743 (
            .O(N__44883),
            .I(N__44850));
    Span4Mux_v I__10742 (
            .O(N__44874),
            .I(N__44847));
    Span4Mux_v I__10741 (
            .O(N__44869),
            .I(N__44844));
    LocalMux I__10740 (
            .O(N__44866),
            .I(N__44839));
    LocalMux I__10739 (
            .O(N__44863),
            .I(N__44839));
    LocalMux I__10738 (
            .O(N__44860),
            .I(N__44834));
    LocalMux I__10737 (
            .O(N__44857),
            .I(N__44834));
    InMux I__10736 (
            .O(N__44856),
            .I(N__44831));
    LocalMux I__10735 (
            .O(N__44853),
            .I(N__44828));
    InMux I__10734 (
            .O(N__44850),
            .I(N__44825));
    Span4Mux_h I__10733 (
            .O(N__44847),
            .I(N__44822));
    Span4Mux_h I__10732 (
            .O(N__44844),
            .I(N__44813));
    Span4Mux_v I__10731 (
            .O(N__44839),
            .I(N__44813));
    Span4Mux_v I__10730 (
            .O(N__44834),
            .I(N__44813));
    LocalMux I__10729 (
            .O(N__44831),
            .I(N__44813));
    Span4Mux_v I__10728 (
            .O(N__44828),
            .I(N__44808));
    LocalMux I__10727 (
            .O(N__44825),
            .I(N__44808));
    Span4Mux_h I__10726 (
            .O(N__44822),
            .I(N__44804));
    Span4Mux_h I__10725 (
            .O(N__44813),
            .I(N__44801));
    Span4Mux_v I__10724 (
            .O(N__44808),
            .I(N__44798));
    InMux I__10723 (
            .O(N__44807),
            .I(N__44795));
    Odrv4 I__10722 (
            .O(N__44804),
            .I(comm_rx_buf_3));
    Odrv4 I__10721 (
            .O(N__44801),
            .I(comm_rx_buf_3));
    Odrv4 I__10720 (
            .O(N__44798),
            .I(comm_rx_buf_3));
    LocalMux I__10719 (
            .O(N__44795),
            .I(comm_rx_buf_3));
    InMux I__10718 (
            .O(N__44786),
            .I(N__44783));
    LocalMux I__10717 (
            .O(N__44783),
            .I(N__44780));
    Odrv4 I__10716 (
            .O(N__44780),
            .I(n4261));
    CascadeMux I__10715 (
            .O(N__44777),
            .I(N__44771));
    InMux I__10714 (
            .O(N__44776),
            .I(N__44768));
    CascadeMux I__10713 (
            .O(N__44775),
            .I(N__44765));
    InMux I__10712 (
            .O(N__44774),
            .I(N__44761));
    InMux I__10711 (
            .O(N__44771),
            .I(N__44758));
    LocalMux I__10710 (
            .O(N__44768),
            .I(N__44755));
    InMux I__10709 (
            .O(N__44765),
            .I(N__44752));
    InMux I__10708 (
            .O(N__44764),
            .I(N__44749));
    LocalMux I__10707 (
            .O(N__44761),
            .I(N__44746));
    LocalMux I__10706 (
            .O(N__44758),
            .I(N__44743));
    Span4Mux_h I__10705 (
            .O(N__44755),
            .I(N__44740));
    LocalMux I__10704 (
            .O(N__44752),
            .I(N__44737));
    LocalMux I__10703 (
            .O(N__44749),
            .I(N__44732));
    Span4Mux_h I__10702 (
            .O(N__44746),
            .I(N__44732));
    Span4Mux_h I__10701 (
            .O(N__44743),
            .I(N__44727));
    Span4Mux_h I__10700 (
            .O(N__44740),
            .I(N__44727));
    Span4Mux_h I__10699 (
            .O(N__44737),
            .I(N__44722));
    Span4Mux_v I__10698 (
            .O(N__44732),
            .I(N__44722));
    Odrv4 I__10697 (
            .O(N__44727),
            .I(comm_buf_1_3));
    Odrv4 I__10696 (
            .O(N__44722),
            .I(comm_buf_1_3));
    CEMux I__10695 (
            .O(N__44717),
            .I(N__44713));
    CEMux I__10694 (
            .O(N__44716),
            .I(N__44708));
    LocalMux I__10693 (
            .O(N__44713),
            .I(N__44705));
    CEMux I__10692 (
            .O(N__44712),
            .I(N__44702));
    CEMux I__10691 (
            .O(N__44711),
            .I(N__44699));
    LocalMux I__10690 (
            .O(N__44708),
            .I(N__44695));
    Span4Mux_v I__10689 (
            .O(N__44705),
            .I(N__44690));
    LocalMux I__10688 (
            .O(N__44702),
            .I(N__44690));
    LocalMux I__10687 (
            .O(N__44699),
            .I(N__44687));
    CEMux I__10686 (
            .O(N__44698),
            .I(N__44684));
    Span4Mux_v I__10685 (
            .O(N__44695),
            .I(N__44681));
    Span4Mux_h I__10684 (
            .O(N__44690),
            .I(N__44678));
    Span4Mux_h I__10683 (
            .O(N__44687),
            .I(N__44673));
    LocalMux I__10682 (
            .O(N__44684),
            .I(N__44673));
    Span4Mux_h I__10681 (
            .O(N__44681),
            .I(N__44670));
    Span4Mux_h I__10680 (
            .O(N__44678),
            .I(N__44667));
    Span4Mux_v I__10679 (
            .O(N__44673),
            .I(N__44664));
    Odrv4 I__10678 (
            .O(N__44670),
            .I(n8702));
    Odrv4 I__10677 (
            .O(N__44667),
            .I(n8702));
    Odrv4 I__10676 (
            .O(N__44664),
            .I(n8702));
    SRMux I__10675 (
            .O(N__44657),
            .I(N__44654));
    LocalMux I__10674 (
            .O(N__44654),
            .I(N__44649));
    SRMux I__10673 (
            .O(N__44653),
            .I(N__44646));
    SRMux I__10672 (
            .O(N__44652),
            .I(N__44642));
    Span4Mux_v I__10671 (
            .O(N__44649),
            .I(N__44636));
    LocalMux I__10670 (
            .O(N__44646),
            .I(N__44636));
    SRMux I__10669 (
            .O(N__44645),
            .I(N__44633));
    LocalMux I__10668 (
            .O(N__44642),
            .I(N__44630));
    SRMux I__10667 (
            .O(N__44641),
            .I(N__44627));
    Span4Mux_h I__10666 (
            .O(N__44636),
            .I(N__44622));
    LocalMux I__10665 (
            .O(N__44633),
            .I(N__44622));
    Span4Mux_v I__10664 (
            .O(N__44630),
            .I(N__44617));
    LocalMux I__10663 (
            .O(N__44627),
            .I(N__44617));
    Span4Mux_h I__10662 (
            .O(N__44622),
            .I(N__44614));
    Span4Mux_h I__10661 (
            .O(N__44617),
            .I(N__44611));
    Span4Mux_h I__10660 (
            .O(N__44614),
            .I(N__44608));
    Odrv4 I__10659 (
            .O(N__44611),
            .I(n10583));
    Odrv4 I__10658 (
            .O(N__44608),
            .I(n10583));
    InMux I__10657 (
            .O(N__44603),
            .I(N__44599));
    CascadeMux I__10656 (
            .O(N__44602),
            .I(N__44596));
    LocalMux I__10655 (
            .O(N__44599),
            .I(N__44593));
    InMux I__10654 (
            .O(N__44596),
            .I(N__44590));
    Span4Mux_h I__10653 (
            .O(N__44593),
            .I(N__44587));
    LocalMux I__10652 (
            .O(N__44590),
            .I(N__44584));
    Span4Mux_h I__10651 (
            .O(N__44587),
            .I(N__44580));
    Span4Mux_v I__10650 (
            .O(N__44584),
            .I(N__44577));
    InMux I__10649 (
            .O(N__44583),
            .I(N__44574));
    Odrv4 I__10648 (
            .O(N__44580),
            .I(cmd_rdadctmp_21));
    Odrv4 I__10647 (
            .O(N__44577),
            .I(cmd_rdadctmp_21));
    LocalMux I__10646 (
            .O(N__44574),
            .I(cmd_rdadctmp_21));
    CascadeMux I__10645 (
            .O(N__44567),
            .I(N__44564));
    InMux I__10644 (
            .O(N__44564),
            .I(N__44560));
    InMux I__10643 (
            .O(N__44563),
            .I(N__44557));
    LocalMux I__10642 (
            .O(N__44560),
            .I(N__44552));
    LocalMux I__10641 (
            .O(N__44557),
            .I(N__44552));
    Odrv4 I__10640 (
            .O(N__44552),
            .I(buf_adcdata1_13));
    CascadeMux I__10639 (
            .O(N__44549),
            .I(N__44546));
    InMux I__10638 (
            .O(N__44546),
            .I(N__44543));
    LocalMux I__10637 (
            .O(N__44543),
            .I(N__44539));
    InMux I__10636 (
            .O(N__44542),
            .I(N__44536));
    Span4Mux_h I__10635 (
            .O(N__44539),
            .I(N__44532));
    LocalMux I__10634 (
            .O(N__44536),
            .I(N__44529));
    CascadeMux I__10633 (
            .O(N__44535),
            .I(N__44526));
    Span4Mux_h I__10632 (
            .O(N__44532),
            .I(N__44523));
    Span4Mux_h I__10631 (
            .O(N__44529),
            .I(N__44520));
    InMux I__10630 (
            .O(N__44526),
            .I(N__44517));
    Odrv4 I__10629 (
            .O(N__44523),
            .I(cmd_rdadctmp_17_adj_1095));
    Odrv4 I__10628 (
            .O(N__44520),
            .I(cmd_rdadctmp_17_adj_1095));
    LocalMux I__10627 (
            .O(N__44517),
            .I(cmd_rdadctmp_17_adj_1095));
    InMux I__10626 (
            .O(N__44510),
            .I(N__44505));
    InMux I__10625 (
            .O(N__44509),
            .I(N__44502));
    CascadeMux I__10624 (
            .O(N__44508),
            .I(N__44499));
    LocalMux I__10623 (
            .O(N__44505),
            .I(N__44494));
    LocalMux I__10622 (
            .O(N__44502),
            .I(N__44494));
    InMux I__10621 (
            .O(N__44499),
            .I(N__44491));
    Odrv12 I__10620 (
            .O(N__44494),
            .I(cmd_rdadctmp_18_adj_1094));
    LocalMux I__10619 (
            .O(N__44491),
            .I(cmd_rdadctmp_18_adj_1094));
    InMux I__10618 (
            .O(N__44486),
            .I(N__44482));
    InMux I__10617 (
            .O(N__44485),
            .I(N__44479));
    LocalMux I__10616 (
            .O(N__44482),
            .I(N__44476));
    LocalMux I__10615 (
            .O(N__44479),
            .I(buf_adcdata2_13));
    Odrv4 I__10614 (
            .O(N__44476),
            .I(buf_adcdata2_13));
    CascadeMux I__10613 (
            .O(N__44471),
            .I(N__44468));
    InMux I__10612 (
            .O(N__44468),
            .I(N__44465));
    LocalMux I__10611 (
            .O(N__44465),
            .I(N__44461));
    InMux I__10610 (
            .O(N__44464),
            .I(N__44458));
    Span4Mux_v I__10609 (
            .O(N__44461),
            .I(N__44455));
    LocalMux I__10608 (
            .O(N__44458),
            .I(N__44452));
    Span4Mux_h I__10607 (
            .O(N__44455),
            .I(N__44448));
    Span4Mux_v I__10606 (
            .O(N__44452),
            .I(N__44445));
    CascadeMux I__10605 (
            .O(N__44451),
            .I(N__44442));
    Sp12to4 I__10604 (
            .O(N__44448),
            .I(N__44439));
    Span4Mux_h I__10603 (
            .O(N__44445),
            .I(N__44436));
    InMux I__10602 (
            .O(N__44442),
            .I(N__44433));
    Odrv12 I__10601 (
            .O(N__44439),
            .I(cmd_rdadctmp_10));
    Odrv4 I__10600 (
            .O(N__44436),
            .I(cmd_rdadctmp_10));
    LocalMux I__10599 (
            .O(N__44433),
            .I(cmd_rdadctmp_10));
    InMux I__10598 (
            .O(N__44426),
            .I(N__44423));
    LocalMux I__10597 (
            .O(N__44423),
            .I(N__44420));
    Span4Mux_h I__10596 (
            .O(N__44420),
            .I(N__44416));
    InMux I__10595 (
            .O(N__44419),
            .I(N__44413));
    Span4Mux_v I__10594 (
            .O(N__44416),
            .I(N__44410));
    LocalMux I__10593 (
            .O(N__44413),
            .I(buf_adcdata1_2));
    Odrv4 I__10592 (
            .O(N__44410),
            .I(buf_adcdata1_2));
    InMux I__10591 (
            .O(N__44405),
            .I(N__44395));
    InMux I__10590 (
            .O(N__44404),
            .I(N__44390));
    InMux I__10589 (
            .O(N__44403),
            .I(N__44390));
    InMux I__10588 (
            .O(N__44402),
            .I(N__44383));
    InMux I__10587 (
            .O(N__44401),
            .I(N__44383));
    InMux I__10586 (
            .O(N__44400),
            .I(N__44383));
    InMux I__10585 (
            .O(N__44399),
            .I(N__44379));
    InMux I__10584 (
            .O(N__44398),
            .I(N__44376));
    LocalMux I__10583 (
            .O(N__44395),
            .I(N__44373));
    LocalMux I__10582 (
            .O(N__44390),
            .I(N__44370));
    LocalMux I__10581 (
            .O(N__44383),
            .I(N__44364));
    InMux I__10580 (
            .O(N__44382),
            .I(N__44361));
    LocalMux I__10579 (
            .O(N__44379),
            .I(N__44348));
    LocalMux I__10578 (
            .O(N__44376),
            .I(N__44345));
    Span4Mux_h I__10577 (
            .O(N__44373),
            .I(N__44340));
    Span4Mux_v I__10576 (
            .O(N__44370),
            .I(N__44340));
    InMux I__10575 (
            .O(N__44369),
            .I(N__44337));
    InMux I__10574 (
            .O(N__44368),
            .I(N__44332));
    InMux I__10573 (
            .O(N__44367),
            .I(N__44332));
    Span4Mux_v I__10572 (
            .O(N__44364),
            .I(N__44326));
    LocalMux I__10571 (
            .O(N__44361),
            .I(N__44326));
    InMux I__10570 (
            .O(N__44360),
            .I(N__44321));
    InMux I__10569 (
            .O(N__44359),
            .I(N__44321));
    InMux I__10568 (
            .O(N__44358),
            .I(N__44314));
    InMux I__10567 (
            .O(N__44357),
            .I(N__44314));
    InMux I__10566 (
            .O(N__44356),
            .I(N__44314));
    InMux I__10565 (
            .O(N__44355),
            .I(N__44311));
    InMux I__10564 (
            .O(N__44354),
            .I(N__44308));
    InMux I__10563 (
            .O(N__44353),
            .I(N__44303));
    InMux I__10562 (
            .O(N__44352),
            .I(N__44303));
    InMux I__10561 (
            .O(N__44351),
            .I(N__44299));
    Span4Mux_h I__10560 (
            .O(N__44348),
            .I(N__44294));
    Span4Mux_v I__10559 (
            .O(N__44345),
            .I(N__44294));
    Span4Mux_h I__10558 (
            .O(N__44340),
            .I(N__44289));
    LocalMux I__10557 (
            .O(N__44337),
            .I(N__44289));
    LocalMux I__10556 (
            .O(N__44332),
            .I(N__44286));
    InMux I__10555 (
            .O(N__44331),
            .I(N__44283));
    Span4Mux_v I__10554 (
            .O(N__44326),
            .I(N__44280));
    LocalMux I__10553 (
            .O(N__44321),
            .I(N__44277));
    LocalMux I__10552 (
            .O(N__44314),
            .I(N__44274));
    LocalMux I__10551 (
            .O(N__44311),
            .I(N__44269));
    LocalMux I__10550 (
            .O(N__44308),
            .I(N__44269));
    LocalMux I__10549 (
            .O(N__44303),
            .I(N__44266));
    InMux I__10548 (
            .O(N__44302),
            .I(N__44263));
    LocalMux I__10547 (
            .O(N__44299),
            .I(N__44260));
    Span4Mux_h I__10546 (
            .O(N__44294),
            .I(N__44255));
    Span4Mux_v I__10545 (
            .O(N__44289),
            .I(N__44255));
    Span4Mux_v I__10544 (
            .O(N__44286),
            .I(N__44250));
    LocalMux I__10543 (
            .O(N__44283),
            .I(N__44250));
    Span4Mux_h I__10542 (
            .O(N__44280),
            .I(N__44247));
    Span4Mux_v I__10541 (
            .O(N__44277),
            .I(N__44244));
    Span4Mux_v I__10540 (
            .O(N__44274),
            .I(N__44241));
    Span4Mux_v I__10539 (
            .O(N__44269),
            .I(N__44236));
    Span4Mux_h I__10538 (
            .O(N__44266),
            .I(N__44236));
    LocalMux I__10537 (
            .O(N__44263),
            .I(N__44233));
    Span4Mux_v I__10536 (
            .O(N__44260),
            .I(N__44230));
    Span4Mux_h I__10535 (
            .O(N__44255),
            .I(N__44225));
    Span4Mux_h I__10534 (
            .O(N__44250),
            .I(N__44225));
    Span4Mux_h I__10533 (
            .O(N__44247),
            .I(N__44214));
    Span4Mux_v I__10532 (
            .O(N__44244),
            .I(N__44214));
    Span4Mux_v I__10531 (
            .O(N__44241),
            .I(N__44214));
    Span4Mux_v I__10530 (
            .O(N__44236),
            .I(N__44214));
    Span4Mux_h I__10529 (
            .O(N__44233),
            .I(N__44214));
    Odrv4 I__10528 (
            .O(N__44230),
            .I(n15147));
    Odrv4 I__10527 (
            .O(N__44225),
            .I(n15147));
    Odrv4 I__10526 (
            .O(N__44214),
            .I(n15147));
    InMux I__10525 (
            .O(N__44207),
            .I(N__44203));
    CascadeMux I__10524 (
            .O(N__44206),
            .I(N__44200));
    LocalMux I__10523 (
            .O(N__44203),
            .I(N__44196));
    InMux I__10522 (
            .O(N__44200),
            .I(N__44193));
    InMux I__10521 (
            .O(N__44199),
            .I(N__44190));
    Span12Mux_v I__10520 (
            .O(N__44196),
            .I(N__44187));
    LocalMux I__10519 (
            .O(N__44193),
            .I(buf_adcdata3_10));
    LocalMux I__10518 (
            .O(N__44190),
            .I(buf_adcdata3_10));
    Odrv12 I__10517 (
            .O(N__44187),
            .I(buf_adcdata3_10));
    InMux I__10516 (
            .O(N__44180),
            .I(N__44175));
    InMux I__10515 (
            .O(N__44179),
            .I(N__44172));
    InMux I__10514 (
            .O(N__44178),
            .I(N__44168));
    LocalMux I__10513 (
            .O(N__44175),
            .I(N__44163));
    LocalMux I__10512 (
            .O(N__44172),
            .I(N__44163));
    InMux I__10511 (
            .O(N__44171),
            .I(N__44160));
    LocalMux I__10510 (
            .O(N__44168),
            .I(N__44152));
    Span4Mux_v I__10509 (
            .O(N__44163),
            .I(N__44146));
    LocalMux I__10508 (
            .O(N__44160),
            .I(N__44146));
    InMux I__10507 (
            .O(N__44159),
            .I(N__44143));
    InMux I__10506 (
            .O(N__44158),
            .I(N__44140));
    InMux I__10505 (
            .O(N__44157),
            .I(N__44136));
    InMux I__10504 (
            .O(N__44156),
            .I(N__44133));
    InMux I__10503 (
            .O(N__44155),
            .I(N__44130));
    Span4Mux_v I__10502 (
            .O(N__44152),
            .I(N__44127));
    InMux I__10501 (
            .O(N__44151),
            .I(N__44124));
    Span4Mux_h I__10500 (
            .O(N__44146),
            .I(N__44119));
    LocalMux I__10499 (
            .O(N__44143),
            .I(N__44119));
    LocalMux I__10498 (
            .O(N__44140),
            .I(N__44116));
    InMux I__10497 (
            .O(N__44139),
            .I(N__44113));
    LocalMux I__10496 (
            .O(N__44136),
            .I(N__44108));
    LocalMux I__10495 (
            .O(N__44133),
            .I(N__44108));
    LocalMux I__10494 (
            .O(N__44130),
            .I(N__44105));
    Span4Mux_h I__10493 (
            .O(N__44127),
            .I(N__44100));
    LocalMux I__10492 (
            .O(N__44124),
            .I(N__44100));
    Span4Mux_h I__10491 (
            .O(N__44119),
            .I(N__44095));
    Span4Mux_h I__10490 (
            .O(N__44116),
            .I(N__44092));
    LocalMux I__10489 (
            .O(N__44113),
            .I(N__44089));
    Span4Mux_v I__10488 (
            .O(N__44108),
            .I(N__44086));
    Span4Mux_h I__10487 (
            .O(N__44105),
            .I(N__44081));
    Span4Mux_v I__10486 (
            .O(N__44100),
            .I(N__44081));
    InMux I__10485 (
            .O(N__44099),
            .I(N__44078));
    InMux I__10484 (
            .O(N__44098),
            .I(N__44075));
    Span4Mux_h I__10483 (
            .O(N__44095),
            .I(N__44071));
    Sp12to4 I__10482 (
            .O(N__44092),
            .I(N__44068));
    Span4Mux_v I__10481 (
            .O(N__44089),
            .I(N__44065));
    Sp12to4 I__10480 (
            .O(N__44086),
            .I(N__44056));
    Sp12to4 I__10479 (
            .O(N__44081),
            .I(N__44056));
    LocalMux I__10478 (
            .O(N__44078),
            .I(N__44056));
    LocalMux I__10477 (
            .O(N__44075),
            .I(N__44056));
    InMux I__10476 (
            .O(N__44074),
            .I(N__44053));
    Odrv4 I__10475 (
            .O(N__44071),
            .I(comm_rx_buf_1));
    Odrv12 I__10474 (
            .O(N__44068),
            .I(comm_rx_buf_1));
    Odrv4 I__10473 (
            .O(N__44065),
            .I(comm_rx_buf_1));
    Odrv12 I__10472 (
            .O(N__44056),
            .I(comm_rx_buf_1));
    LocalMux I__10471 (
            .O(N__44053),
            .I(comm_rx_buf_1));
    CascadeMux I__10470 (
            .O(N__44042),
            .I(N__44036));
    InMux I__10469 (
            .O(N__44041),
            .I(N__44029));
    InMux I__10468 (
            .O(N__44040),
            .I(N__44024));
    InMux I__10467 (
            .O(N__44039),
            .I(N__44024));
    InMux I__10466 (
            .O(N__44036),
            .I(N__44021));
    InMux I__10465 (
            .O(N__44035),
            .I(N__44012));
    InMux I__10464 (
            .O(N__44034),
            .I(N__44012));
    InMux I__10463 (
            .O(N__44033),
            .I(N__44012));
    InMux I__10462 (
            .O(N__44032),
            .I(N__44012));
    LocalMux I__10461 (
            .O(N__44029),
            .I(n8618));
    LocalMux I__10460 (
            .O(N__44024),
            .I(n8618));
    LocalMux I__10459 (
            .O(N__44021),
            .I(n8618));
    LocalMux I__10458 (
            .O(N__44012),
            .I(n8618));
    CascadeMux I__10457 (
            .O(N__44003),
            .I(N__43998));
    CascadeMux I__10456 (
            .O(N__44002),
            .I(N__43991));
    InMux I__10455 (
            .O(N__44001),
            .I(N__43988));
    InMux I__10454 (
            .O(N__43998),
            .I(N__43981));
    InMux I__10453 (
            .O(N__43997),
            .I(N__43981));
    InMux I__10452 (
            .O(N__43996),
            .I(N__43981));
    InMux I__10451 (
            .O(N__43995),
            .I(N__43974));
    InMux I__10450 (
            .O(N__43994),
            .I(N__43974));
    InMux I__10449 (
            .O(N__43991),
            .I(N__43974));
    LocalMux I__10448 (
            .O(N__43988),
            .I(n10363));
    LocalMux I__10447 (
            .O(N__43981),
            .I(n10363));
    LocalMux I__10446 (
            .O(N__43974),
            .I(n10363));
    InMux I__10445 (
            .O(N__43967),
            .I(N__43963));
    CascadeMux I__10444 (
            .O(N__43966),
            .I(N__43959));
    LocalMux I__10443 (
            .O(N__43963),
            .I(N__43956));
    CascadeMux I__10442 (
            .O(N__43962),
            .I(N__43953));
    InMux I__10441 (
            .O(N__43959),
            .I(N__43950));
    Span12Mux_v I__10440 (
            .O(N__43956),
            .I(N__43947));
    InMux I__10439 (
            .O(N__43953),
            .I(N__43944));
    LocalMux I__10438 (
            .O(N__43950),
            .I(cmd_rdadctmp_25_adj_1051));
    Odrv12 I__10437 (
            .O(N__43947),
            .I(cmd_rdadctmp_25_adj_1051));
    LocalMux I__10436 (
            .O(N__43944),
            .I(cmd_rdadctmp_25_adj_1051));
    InMux I__10435 (
            .O(N__43937),
            .I(N__43933));
    CascadeMux I__10434 (
            .O(N__43936),
            .I(N__43930));
    LocalMux I__10433 (
            .O(N__43933),
            .I(N__43927));
    InMux I__10432 (
            .O(N__43930),
            .I(N__43924));
    Span4Mux_h I__10431 (
            .O(N__43927),
            .I(N__43921));
    LocalMux I__10430 (
            .O(N__43924),
            .I(buf_adcdata2_18));
    Odrv4 I__10429 (
            .O(N__43921),
            .I(buf_adcdata2_18));
    CascadeMux I__10428 (
            .O(N__43916),
            .I(N__43913));
    InMux I__10427 (
            .O(N__43913),
            .I(N__43910));
    LocalMux I__10426 (
            .O(N__43910),
            .I(N__43906));
    InMux I__10425 (
            .O(N__43909),
            .I(N__43903));
    Span4Mux_h I__10424 (
            .O(N__43906),
            .I(N__43900));
    LocalMux I__10423 (
            .O(N__43903),
            .I(N__43897));
    Odrv4 I__10422 (
            .O(N__43900),
            .I(n14_adj_1215));
    Odrv12 I__10421 (
            .O(N__43897),
            .I(n14_adj_1215));
    CascadeMux I__10420 (
            .O(N__43892),
            .I(N__43887));
    InMux I__10419 (
            .O(N__43891),
            .I(N__43880));
    InMux I__10418 (
            .O(N__43890),
            .I(N__43880));
    InMux I__10417 (
            .O(N__43887),
            .I(N__43880));
    LocalMux I__10416 (
            .O(N__43880),
            .I(cmd_rdadctmp_26_adj_1050));
    CascadeMux I__10415 (
            .O(N__43877),
            .I(N__43874));
    InMux I__10414 (
            .O(N__43874),
            .I(N__43870));
    CascadeMux I__10413 (
            .O(N__43873),
            .I(N__43866));
    LocalMux I__10412 (
            .O(N__43870),
            .I(N__43863));
    InMux I__10411 (
            .O(N__43869),
            .I(N__43858));
    InMux I__10410 (
            .O(N__43866),
            .I(N__43858));
    Odrv4 I__10409 (
            .O(N__43863),
            .I(cmd_rdadctmp_27_adj_1049));
    LocalMux I__10408 (
            .O(N__43858),
            .I(cmd_rdadctmp_27_adj_1049));
    CascadeMux I__10407 (
            .O(N__43853),
            .I(N__43850));
    InMux I__10406 (
            .O(N__43850),
            .I(N__43847));
    LocalMux I__10405 (
            .O(N__43847),
            .I(N__43844));
    Span4Mux_v I__10404 (
            .O(N__43844),
            .I(N__43841));
    Span4Mux_h I__10403 (
            .O(N__43841),
            .I(N__43837));
    CascadeMux I__10402 (
            .O(N__43840),
            .I(N__43834));
    Span4Mux_h I__10401 (
            .O(N__43837),
            .I(N__43831));
    InMux I__10400 (
            .O(N__43834),
            .I(N__43828));
    Span4Mux_h I__10399 (
            .O(N__43831),
            .I(N__43822));
    LocalMux I__10398 (
            .O(N__43828),
            .I(N__43822));
    InMux I__10397 (
            .O(N__43827),
            .I(N__43819));
    Odrv4 I__10396 (
            .O(N__43822),
            .I(cmd_rdadctmp_8_adj_1104));
    LocalMux I__10395 (
            .O(N__43819),
            .I(cmd_rdadctmp_8_adj_1104));
    InMux I__10394 (
            .O(N__43814),
            .I(N__43811));
    LocalMux I__10393 (
            .O(N__43811),
            .I(N__43807));
    InMux I__10392 (
            .O(N__43810),
            .I(N__43804));
    Sp12to4 I__10391 (
            .O(N__43807),
            .I(N__43801));
    LocalMux I__10390 (
            .O(N__43804),
            .I(N__43797));
    Span12Mux_v I__10389 (
            .O(N__43801),
            .I(N__43794));
    InMux I__10388 (
            .O(N__43800),
            .I(N__43791));
    Span4Mux_h I__10387 (
            .O(N__43797),
            .I(N__43788));
    Span12Mux_h I__10386 (
            .O(N__43794),
            .I(N__43785));
    LocalMux I__10385 (
            .O(N__43791),
            .I(buf_adcdata3_0));
    Odrv4 I__10384 (
            .O(N__43788),
            .I(buf_adcdata3_0));
    Odrv12 I__10383 (
            .O(N__43785),
            .I(buf_adcdata3_0));
    InMux I__10382 (
            .O(N__43778),
            .I(N__43775));
    LocalMux I__10381 (
            .O(N__43775),
            .I(N__43771));
    InMux I__10380 (
            .O(N__43774),
            .I(N__43768));
    Span4Mux_h I__10379 (
            .O(N__43771),
            .I(N__43764));
    LocalMux I__10378 (
            .O(N__43768),
            .I(N__43761));
    InMux I__10377 (
            .O(N__43767),
            .I(N__43758));
    Span4Mux_v I__10376 (
            .O(N__43764),
            .I(N__43753));
    Span4Mux_h I__10375 (
            .O(N__43761),
            .I(N__43753));
    LocalMux I__10374 (
            .O(N__43758),
            .I(buf_adcdata3_11));
    Odrv4 I__10373 (
            .O(N__43753),
            .I(buf_adcdata3_11));
    CascadeMux I__10372 (
            .O(N__43748),
            .I(N__43745));
    InMux I__10371 (
            .O(N__43745),
            .I(N__43742));
    LocalMux I__10370 (
            .O(N__43742),
            .I(N__43739));
    Span4Mux_v I__10369 (
            .O(N__43739),
            .I(N__43735));
    CascadeMux I__10368 (
            .O(N__43738),
            .I(N__43731));
    Span4Mux_h I__10367 (
            .O(N__43735),
            .I(N__43728));
    InMux I__10366 (
            .O(N__43734),
            .I(N__43723));
    InMux I__10365 (
            .O(N__43731),
            .I(N__43723));
    Odrv4 I__10364 (
            .O(N__43728),
            .I(cmd_rdadctmp_30_adj_1082));
    LocalMux I__10363 (
            .O(N__43723),
            .I(cmd_rdadctmp_30_adj_1082));
    InMux I__10362 (
            .O(N__43718),
            .I(N__43715));
    LocalMux I__10361 (
            .O(N__43715),
            .I(N__43712));
    Span4Mux_h I__10360 (
            .O(N__43712),
            .I(N__43709));
    Span4Mux_v I__10359 (
            .O(N__43709),
            .I(N__43704));
    InMux I__10358 (
            .O(N__43708),
            .I(N__43699));
    InMux I__10357 (
            .O(N__43707),
            .I(N__43699));
    Odrv4 I__10356 (
            .O(N__43704),
            .I(buf_adcdata3_22));
    LocalMux I__10355 (
            .O(N__43699),
            .I(buf_adcdata3_22));
    InMux I__10354 (
            .O(N__43694),
            .I(N__43691));
    LocalMux I__10353 (
            .O(N__43691),
            .I(N__43688));
    Odrv4 I__10352 (
            .O(N__43688),
            .I(n7_adj_1190));
    InMux I__10351 (
            .O(N__43685),
            .I(N__43682));
    LocalMux I__10350 (
            .O(N__43682),
            .I(N__43678));
    InMux I__10349 (
            .O(N__43681),
            .I(N__43674));
    Span4Mux_h I__10348 (
            .O(N__43678),
            .I(N__43671));
    InMux I__10347 (
            .O(N__43677),
            .I(N__43668));
    LocalMux I__10346 (
            .O(N__43674),
            .I(buf_dds_2));
    Odrv4 I__10345 (
            .O(N__43671),
            .I(buf_dds_2));
    LocalMux I__10344 (
            .O(N__43668),
            .I(buf_dds_2));
    CascadeMux I__10343 (
            .O(N__43661),
            .I(N__43658));
    InMux I__10342 (
            .O(N__43658),
            .I(N__43655));
    LocalMux I__10341 (
            .O(N__43655),
            .I(N__43652));
    Span4Mux_v I__10340 (
            .O(N__43652),
            .I(N__43649));
    Span4Mux_h I__10339 (
            .O(N__43649),
            .I(N__43646));
    Odrv4 I__10338 (
            .O(N__43646),
            .I(n4207));
    InMux I__10337 (
            .O(N__43643),
            .I(N__43640));
    LocalMux I__10336 (
            .O(N__43640),
            .I(N__43637));
    Span4Mux_v I__10335 (
            .O(N__43637),
            .I(N__43632));
    InMux I__10334 (
            .O(N__43636),
            .I(N__43629));
    InMux I__10333 (
            .O(N__43635),
            .I(N__43626));
    Span4Mux_h I__10332 (
            .O(N__43632),
            .I(N__43621));
    LocalMux I__10331 (
            .O(N__43629),
            .I(N__43621));
    LocalMux I__10330 (
            .O(N__43626),
            .I(n8094));
    Odrv4 I__10329 (
            .O(N__43621),
            .I(n8094));
    InMux I__10328 (
            .O(N__43616),
            .I(N__43611));
    InMux I__10327 (
            .O(N__43615),
            .I(N__43608));
    InMux I__10326 (
            .O(N__43614),
            .I(N__43605));
    LocalMux I__10325 (
            .O(N__43611),
            .I(N__43602));
    LocalMux I__10324 (
            .O(N__43608),
            .I(N__43599));
    LocalMux I__10323 (
            .O(N__43605),
            .I(N__43596));
    Span4Mux_v I__10322 (
            .O(N__43602),
            .I(N__43593));
    Span4Mux_h I__10321 (
            .O(N__43599),
            .I(N__43590));
    Span4Mux_v I__10320 (
            .O(N__43596),
            .I(N__43585));
    Span4Mux_h I__10319 (
            .O(N__43593),
            .I(N__43585));
    Odrv4 I__10318 (
            .O(N__43590),
            .I(n729));
    Odrv4 I__10317 (
            .O(N__43585),
            .I(n729));
    InMux I__10316 (
            .O(N__43580),
            .I(N__43577));
    LocalMux I__10315 (
            .O(N__43577),
            .I(N__43573));
    InMux I__10314 (
            .O(N__43576),
            .I(N__43570));
    Span4Mux_h I__10313 (
            .O(N__43573),
            .I(N__43567));
    LocalMux I__10312 (
            .O(N__43570),
            .I(buf_adcdata2_19));
    Odrv4 I__10311 (
            .O(N__43567),
            .I(buf_adcdata2_19));
    InMux I__10310 (
            .O(N__43562),
            .I(N__43555));
    CascadeMux I__10309 (
            .O(N__43561),
            .I(N__43552));
    InMux I__10308 (
            .O(N__43560),
            .I(N__43549));
    InMux I__10307 (
            .O(N__43559),
            .I(N__43546));
    InMux I__10306 (
            .O(N__43558),
            .I(N__43543));
    LocalMux I__10305 (
            .O(N__43555),
            .I(N__43540));
    InMux I__10304 (
            .O(N__43552),
            .I(N__43537));
    LocalMux I__10303 (
            .O(N__43549),
            .I(N__43534));
    LocalMux I__10302 (
            .O(N__43546),
            .I(N__43529));
    LocalMux I__10301 (
            .O(N__43543),
            .I(N__43526));
    Span4Mux_h I__10300 (
            .O(N__43540),
            .I(N__43523));
    LocalMux I__10299 (
            .O(N__43537),
            .I(N__43518));
    Span4Mux_v I__10298 (
            .O(N__43534),
            .I(N__43518));
    InMux I__10297 (
            .O(N__43533),
            .I(N__43515));
    InMux I__10296 (
            .O(N__43532),
            .I(N__43512));
    Span12Mux_v I__10295 (
            .O(N__43529),
            .I(N__43509));
    Span4Mux_h I__10294 (
            .O(N__43526),
            .I(N__43502));
    Span4Mux_h I__10293 (
            .O(N__43523),
            .I(N__43502));
    Span4Mux_h I__10292 (
            .O(N__43518),
            .I(N__43502));
    LocalMux I__10291 (
            .O(N__43515),
            .I(comm_buf_0_3));
    LocalMux I__10290 (
            .O(N__43512),
            .I(comm_buf_0_3));
    Odrv12 I__10289 (
            .O(N__43509),
            .I(comm_buf_0_3));
    Odrv4 I__10288 (
            .O(N__43502),
            .I(comm_buf_0_3));
    InMux I__10287 (
            .O(N__43493),
            .I(N__43489));
    InMux I__10286 (
            .O(N__43492),
            .I(N__43486));
    LocalMux I__10285 (
            .O(N__43489),
            .I(N__43481));
    LocalMux I__10284 (
            .O(N__43486),
            .I(N__43481));
    Span4Mux_v I__10283 (
            .O(N__43481),
            .I(N__43478));
    Span4Mux_h I__10282 (
            .O(N__43478),
            .I(N__43475));
    Odrv4 I__10281 (
            .O(N__43475),
            .I(n14_adj_1208));
    CascadeMux I__10280 (
            .O(N__43472),
            .I(n26_adj_1192_cascade_));
    CEMux I__10279 (
            .O(N__43469),
            .I(N__43466));
    LocalMux I__10278 (
            .O(N__43466),
            .I(N__43463));
    Odrv4 I__10277 (
            .O(N__43463),
            .I(n18_adj_1191));
    InMux I__10276 (
            .O(N__43460),
            .I(N__43457));
    LocalMux I__10275 (
            .O(N__43457),
            .I(n15245));
    InMux I__10274 (
            .O(N__43454),
            .I(N__43451));
    LocalMux I__10273 (
            .O(N__43451),
            .I(N__43442));
    InMux I__10272 (
            .O(N__43450),
            .I(N__43433));
    InMux I__10271 (
            .O(N__43449),
            .I(N__43430));
    InMux I__10270 (
            .O(N__43448),
            .I(N__43421));
    InMux I__10269 (
            .O(N__43447),
            .I(N__43421));
    InMux I__10268 (
            .O(N__43446),
            .I(N__43421));
    InMux I__10267 (
            .O(N__43445),
            .I(N__43421));
    Span4Mux_v I__10266 (
            .O(N__43442),
            .I(N__43418));
    InMux I__10265 (
            .O(N__43441),
            .I(N__43413));
    InMux I__10264 (
            .O(N__43440),
            .I(N__43413));
    CascadeMux I__10263 (
            .O(N__43439),
            .I(N__43410));
    CascadeMux I__10262 (
            .O(N__43438),
            .I(N__43407));
    CascadeMux I__10261 (
            .O(N__43437),
            .I(N__43403));
    CascadeMux I__10260 (
            .O(N__43436),
            .I(N__43399));
    LocalMux I__10259 (
            .O(N__43433),
            .I(N__43395));
    LocalMux I__10258 (
            .O(N__43430),
            .I(N__43388));
    LocalMux I__10257 (
            .O(N__43421),
            .I(N__43385));
    Span4Mux_v I__10256 (
            .O(N__43418),
            .I(N__43380));
    LocalMux I__10255 (
            .O(N__43413),
            .I(N__43380));
    InMux I__10254 (
            .O(N__43410),
            .I(N__43376));
    InMux I__10253 (
            .O(N__43407),
            .I(N__43371));
    InMux I__10252 (
            .O(N__43406),
            .I(N__43371));
    InMux I__10251 (
            .O(N__43403),
            .I(N__43362));
    InMux I__10250 (
            .O(N__43402),
            .I(N__43362));
    InMux I__10249 (
            .O(N__43399),
            .I(N__43362));
    InMux I__10248 (
            .O(N__43398),
            .I(N__43362));
    Sp12to4 I__10247 (
            .O(N__43395),
            .I(N__43359));
    InMux I__10246 (
            .O(N__43394),
            .I(N__43350));
    InMux I__10245 (
            .O(N__43393),
            .I(N__43350));
    InMux I__10244 (
            .O(N__43392),
            .I(N__43350));
    InMux I__10243 (
            .O(N__43391),
            .I(N__43350));
    Span4Mux_v I__10242 (
            .O(N__43388),
            .I(N__43343));
    Span4Mux_v I__10241 (
            .O(N__43385),
            .I(N__43343));
    Span4Mux_h I__10240 (
            .O(N__43380),
            .I(N__43343));
    InMux I__10239 (
            .O(N__43379),
            .I(N__43340));
    LocalMux I__10238 (
            .O(N__43376),
            .I(N__43333));
    LocalMux I__10237 (
            .O(N__43371),
            .I(N__43333));
    LocalMux I__10236 (
            .O(N__43362),
            .I(N__43333));
    Span12Mux_h I__10235 (
            .O(N__43359),
            .I(N__43330));
    LocalMux I__10234 (
            .O(N__43350),
            .I(N__43323));
    Sp12to4 I__10233 (
            .O(N__43343),
            .I(N__43323));
    LocalMux I__10232 (
            .O(N__43340),
            .I(N__43323));
    Span12Mux_h I__10231 (
            .O(N__43333),
            .I(N__43320));
    Span12Mux_v I__10230 (
            .O(N__43330),
            .I(N__43317));
    Span12Mux_v I__10229 (
            .O(N__43323),
            .I(N__43314));
    Span12Mux_v I__10228 (
            .O(N__43320),
            .I(N__43311));
    Odrv12 I__10227 (
            .O(N__43317),
            .I(ICE_SPI_CE0));
    Odrv12 I__10226 (
            .O(N__43314),
            .I(ICE_SPI_CE0));
    Odrv12 I__10225 (
            .O(N__43311),
            .I(ICE_SPI_CE0));
    CascadeMux I__10224 (
            .O(N__43304),
            .I(n15245_cascade_));
    InMux I__10223 (
            .O(N__43301),
            .I(N__43290));
    InMux I__10222 (
            .O(N__43300),
            .I(N__43290));
    InMux I__10221 (
            .O(N__43299),
            .I(N__43290));
    InMux I__10220 (
            .O(N__43298),
            .I(N__43282));
    InMux I__10219 (
            .O(N__43297),
            .I(N__43282));
    LocalMux I__10218 (
            .O(N__43290),
            .I(N__43278));
    InMux I__10217 (
            .O(N__43289),
            .I(N__43275));
    InMux I__10216 (
            .O(N__43288),
            .I(N__43272));
    InMux I__10215 (
            .O(N__43287),
            .I(N__43269));
    LocalMux I__10214 (
            .O(N__43282),
            .I(N__43262));
    InMux I__10213 (
            .O(N__43281),
            .I(N__43259));
    Span4Mux_h I__10212 (
            .O(N__43278),
            .I(N__43256));
    LocalMux I__10211 (
            .O(N__43275),
            .I(N__43248));
    LocalMux I__10210 (
            .O(N__43272),
            .I(N__43248));
    LocalMux I__10209 (
            .O(N__43269),
            .I(N__43248));
    InMux I__10208 (
            .O(N__43268),
            .I(N__43239));
    InMux I__10207 (
            .O(N__43267),
            .I(N__43239));
    InMux I__10206 (
            .O(N__43266),
            .I(N__43239));
    InMux I__10205 (
            .O(N__43265),
            .I(N__43239));
    Span4Mux_v I__10204 (
            .O(N__43262),
            .I(N__43235));
    LocalMux I__10203 (
            .O(N__43259),
            .I(N__43232));
    Span4Mux_h I__10202 (
            .O(N__43256),
            .I(N__43229));
    InMux I__10201 (
            .O(N__43255),
            .I(N__43226));
    Span4Mux_v I__10200 (
            .O(N__43248),
            .I(N__43221));
    LocalMux I__10199 (
            .O(N__43239),
            .I(N__43221));
    InMux I__10198 (
            .O(N__43238),
            .I(N__43218));
    Odrv4 I__10197 (
            .O(N__43235),
            .I(comm_data_vld));
    Odrv4 I__10196 (
            .O(N__43232),
            .I(comm_data_vld));
    Odrv4 I__10195 (
            .O(N__43229),
            .I(comm_data_vld));
    LocalMux I__10194 (
            .O(N__43226),
            .I(comm_data_vld));
    Odrv4 I__10193 (
            .O(N__43221),
            .I(comm_data_vld));
    LocalMux I__10192 (
            .O(N__43218),
            .I(comm_data_vld));
    InMux I__10191 (
            .O(N__43205),
            .I(N__43202));
    LocalMux I__10190 (
            .O(N__43202),
            .I(n8544));
    InMux I__10189 (
            .O(N__43199),
            .I(N__43194));
    InMux I__10188 (
            .O(N__43198),
            .I(N__43189));
    InMux I__10187 (
            .O(N__43197),
            .I(N__43189));
    LocalMux I__10186 (
            .O(N__43194),
            .I(N__43185));
    LocalMux I__10185 (
            .O(N__43189),
            .I(N__43182));
    InMux I__10184 (
            .O(N__43188),
            .I(N__43179));
    Span4Mux_v I__10183 (
            .O(N__43185),
            .I(N__43174));
    Span4Mux_v I__10182 (
            .O(N__43182),
            .I(N__43174));
    LocalMux I__10181 (
            .O(N__43179),
            .I(N__43171));
    Odrv4 I__10180 (
            .O(N__43174),
            .I(n9_adj_1028));
    Odrv12 I__10179 (
            .O(N__43171),
            .I(n9_adj_1028));
    CascadeMux I__10178 (
            .O(N__43166),
            .I(N__43162));
    InMux I__10177 (
            .O(N__43165),
            .I(N__43159));
    InMux I__10176 (
            .O(N__43162),
            .I(N__43156));
    LocalMux I__10175 (
            .O(N__43159),
            .I(N__43153));
    LocalMux I__10174 (
            .O(N__43156),
            .I(N__43150));
    Span4Mux_h I__10173 (
            .O(N__43153),
            .I(N__43145));
    Span4Mux_v I__10172 (
            .O(N__43150),
            .I(N__43145));
    Odrv4 I__10171 (
            .O(N__43145),
            .I(n9011));
    CascadeMux I__10170 (
            .O(N__43142),
            .I(n9011_cascade_));
    CEMux I__10169 (
            .O(N__43139),
            .I(N__43135));
    CEMux I__10168 (
            .O(N__43138),
            .I(N__43131));
    LocalMux I__10167 (
            .O(N__43135),
            .I(N__43128));
    CEMux I__10166 (
            .O(N__43134),
            .I(N__43123));
    LocalMux I__10165 (
            .O(N__43131),
            .I(N__43117));
    Span4Mux_v I__10164 (
            .O(N__43128),
            .I(N__43117));
    CEMux I__10163 (
            .O(N__43127),
            .I(N__43114));
    CEMux I__10162 (
            .O(N__43126),
            .I(N__43111));
    LocalMux I__10161 (
            .O(N__43123),
            .I(N__43106));
    CEMux I__10160 (
            .O(N__43122),
            .I(N__43103));
    Span4Mux_h I__10159 (
            .O(N__43117),
            .I(N__43096));
    LocalMux I__10158 (
            .O(N__43114),
            .I(N__43096));
    LocalMux I__10157 (
            .O(N__43111),
            .I(N__43096));
    CEMux I__10156 (
            .O(N__43110),
            .I(N__43093));
    CEMux I__10155 (
            .O(N__43109),
            .I(N__43090));
    Span4Mux_v I__10154 (
            .O(N__43106),
            .I(N__43085));
    LocalMux I__10153 (
            .O(N__43103),
            .I(N__43085));
    Span4Mux_v I__10152 (
            .O(N__43096),
            .I(N__43082));
    LocalMux I__10151 (
            .O(N__43093),
            .I(N__43079));
    LocalMux I__10150 (
            .O(N__43090),
            .I(N__43075));
    Span4Mux_v I__10149 (
            .O(N__43085),
            .I(N__43072));
    Sp12to4 I__10148 (
            .O(N__43082),
            .I(N__43069));
    Sp12to4 I__10147 (
            .O(N__43079),
            .I(N__43066));
    InMux I__10146 (
            .O(N__43078),
            .I(N__43063));
    Sp12to4 I__10145 (
            .O(N__43075),
            .I(N__43058));
    Sp12to4 I__10144 (
            .O(N__43072),
            .I(N__43058));
    Span12Mux_v I__10143 (
            .O(N__43069),
            .I(N__43051));
    Span12Mux_v I__10142 (
            .O(N__43066),
            .I(N__43051));
    LocalMux I__10141 (
            .O(N__43063),
            .I(N__43051));
    Span12Mux_h I__10140 (
            .O(N__43058),
            .I(N__43048));
    Span12Mux_h I__10139 (
            .O(N__43051),
            .I(N__43045));
    Odrv12 I__10138 (
            .O(N__43048),
            .I(n9215));
    Odrv12 I__10137 (
            .O(N__43045),
            .I(n9215));
    InMux I__10136 (
            .O(N__43040),
            .I(N__43037));
    LocalMux I__10135 (
            .O(N__43037),
            .I(N__43034));
    Odrv4 I__10134 (
            .O(N__43034),
            .I(buf_data2_19));
    InMux I__10133 (
            .O(N__43031),
            .I(N__43028));
    LocalMux I__10132 (
            .O(N__43028),
            .I(N__43025));
    Span4Mux_h I__10131 (
            .O(N__43025),
            .I(N__43021));
    InMux I__10130 (
            .O(N__43024),
            .I(N__43018));
    Sp12to4 I__10129 (
            .O(N__43021),
            .I(N__43012));
    LocalMux I__10128 (
            .O(N__43018),
            .I(N__43012));
    InMux I__10127 (
            .O(N__43017),
            .I(N__43009));
    Span12Mux_v I__10126 (
            .O(N__43012),
            .I(N__43006));
    LocalMux I__10125 (
            .O(N__43009),
            .I(buf_adcdata4_19));
    Odrv12 I__10124 (
            .O(N__43006),
            .I(buf_adcdata4_19));
    InMux I__10123 (
            .O(N__43001),
            .I(N__42998));
    LocalMux I__10122 (
            .O(N__42998),
            .I(N__42995));
    Sp12to4 I__10121 (
            .O(N__42995),
            .I(N__42992));
    Span12Mux_v I__10120 (
            .O(N__42992),
            .I(N__42989));
    Odrv12 I__10119 (
            .O(N__42989),
            .I(comm_buf_3_7_N_501_3));
    CascadeMux I__10118 (
            .O(N__42986),
            .I(N__42982));
    CascadeMux I__10117 (
            .O(N__42985),
            .I(N__42979));
    InMux I__10116 (
            .O(N__42982),
            .I(N__42976));
    InMux I__10115 (
            .O(N__42979),
            .I(N__42973));
    LocalMux I__10114 (
            .O(N__42976),
            .I(buf_control_6));
    LocalMux I__10113 (
            .O(N__42973),
            .I(buf_control_6));
    InMux I__10112 (
            .O(N__42968),
            .I(N__42965));
    LocalMux I__10111 (
            .O(N__42965),
            .I(N__42962));
    Span4Mux_h I__10110 (
            .O(N__42962),
            .I(N__42959));
    Span4Mux_h I__10109 (
            .O(N__42959),
            .I(N__42956));
    Odrv4 I__10108 (
            .O(N__42956),
            .I(n60));
    SRMux I__10107 (
            .O(N__42953),
            .I(N__42950));
    LocalMux I__10106 (
            .O(N__42950),
            .I(N__42947));
    Odrv12 I__10105 (
            .O(N__42947),
            .I(\comm_spi.imosi_N_791 ));
    CascadeMux I__10104 (
            .O(N__42944),
            .I(N__42941));
    InMux I__10103 (
            .O(N__42941),
            .I(N__42938));
    LocalMux I__10102 (
            .O(N__42938),
            .I(N__42935));
    Span4Mux_v I__10101 (
            .O(N__42935),
            .I(N__42932));
    Sp12to4 I__10100 (
            .O(N__42932),
            .I(N__42928));
    CascadeMux I__10099 (
            .O(N__42931),
            .I(N__42924));
    Span12Mux_h I__10098 (
            .O(N__42928),
            .I(N__42921));
    InMux I__10097 (
            .O(N__42927),
            .I(N__42916));
    InMux I__10096 (
            .O(N__42924),
            .I(N__42916));
    Span12Mux_h I__10095 (
            .O(N__42921),
            .I(N__42913));
    LocalMux I__10094 (
            .O(N__42916),
            .I(cmd_rdadctmp_9_adj_1067));
    Odrv12 I__10093 (
            .O(N__42913),
            .I(cmd_rdadctmp_9_adj_1067));
    InMux I__10092 (
            .O(N__42908),
            .I(N__42905));
    LocalMux I__10091 (
            .O(N__42905),
            .I(N__42901));
    InMux I__10090 (
            .O(N__42904),
            .I(N__42898));
    Span4Mux_v I__10089 (
            .O(N__42901),
            .I(N__42895));
    LocalMux I__10088 (
            .O(N__42898),
            .I(buf_adcdata2_1));
    Odrv4 I__10087 (
            .O(N__42895),
            .I(buf_adcdata2_1));
    InMux I__10086 (
            .O(N__42890),
            .I(N__42886));
    InMux I__10085 (
            .O(N__42889),
            .I(N__42883));
    LocalMux I__10084 (
            .O(N__42886),
            .I(\comm_spi.imosi ));
    LocalMux I__10083 (
            .O(N__42883),
            .I(\comm_spi.imosi ));
    SRMux I__10082 (
            .O(N__42878),
            .I(N__42875));
    LocalMux I__10081 (
            .O(N__42875),
            .I(N__42872));
    Span4Mux_h I__10080 (
            .O(N__42872),
            .I(N__42869));
    Span4Mux_h I__10079 (
            .O(N__42869),
            .I(N__42866));
    Odrv4 I__10078 (
            .O(N__42866),
            .I(\comm_spi.DOUT_7__N_786 ));
    InMux I__10077 (
            .O(N__42863),
            .I(N__42857));
    InMux I__10076 (
            .O(N__42862),
            .I(N__42857));
    LocalMux I__10075 (
            .O(N__42857),
            .I(N__42853));
    InMux I__10074 (
            .O(N__42856),
            .I(N__42850));
    Span4Mux_v I__10073 (
            .O(N__42853),
            .I(N__42846));
    LocalMux I__10072 (
            .O(N__42850),
            .I(N__42843));
    InMux I__10071 (
            .O(N__42849),
            .I(N__42840));
    Span4Mux_h I__10070 (
            .O(N__42846),
            .I(N__42833));
    Span4Mux_v I__10069 (
            .O(N__42843),
            .I(N__42833));
    LocalMux I__10068 (
            .O(N__42840),
            .I(N__42830));
    InMux I__10067 (
            .O(N__42839),
            .I(N__42825));
    InMux I__10066 (
            .O(N__42838),
            .I(N__42825));
    Sp12to4 I__10065 (
            .O(N__42833),
            .I(N__42820));
    Span12Mux_h I__10064 (
            .O(N__42830),
            .I(N__42820));
    LocalMux I__10063 (
            .O(N__42825),
            .I(n15131));
    Odrv12 I__10062 (
            .O(N__42820),
            .I(n15131));
    CascadeMux I__10061 (
            .O(N__42815),
            .I(N__42812));
    InMux I__10060 (
            .O(N__42812),
            .I(N__42808));
    InMux I__10059 (
            .O(N__42811),
            .I(N__42805));
    LocalMux I__10058 (
            .O(N__42808),
            .I(n15241));
    LocalMux I__10057 (
            .O(N__42805),
            .I(n15241));
    InMux I__10056 (
            .O(N__42800),
            .I(N__42788));
    InMux I__10055 (
            .O(N__42799),
            .I(N__42788));
    InMux I__10054 (
            .O(N__42798),
            .I(N__42788));
    InMux I__10053 (
            .O(N__42797),
            .I(N__42785));
    InMux I__10052 (
            .O(N__42796),
            .I(N__42780));
    InMux I__10051 (
            .O(N__42795),
            .I(N__42780));
    LocalMux I__10050 (
            .O(N__42788),
            .I(N__42775));
    LocalMux I__10049 (
            .O(N__42785),
            .I(N__42775));
    LocalMux I__10048 (
            .O(N__42780),
            .I(N__42772));
    Span4Mux_h I__10047 (
            .O(N__42775),
            .I(N__42769));
    Span4Mux_h I__10046 (
            .O(N__42772),
            .I(N__42766));
    Span4Mux_h I__10045 (
            .O(N__42769),
            .I(N__42763));
    Span4Mux_h I__10044 (
            .O(N__42766),
            .I(N__42760));
    Odrv4 I__10043 (
            .O(N__42763),
            .I(n15191));
    Odrv4 I__10042 (
            .O(N__42760),
            .I(n15191));
    CascadeMux I__10041 (
            .O(N__42755),
            .I(N__42752));
    InMux I__10040 (
            .O(N__42752),
            .I(N__42749));
    LocalMux I__10039 (
            .O(N__42749),
            .I(N__42745));
    CascadeMux I__10038 (
            .O(N__42748),
            .I(N__42742));
    Span4Mux_v I__10037 (
            .O(N__42745),
            .I(N__42739));
    InMux I__10036 (
            .O(N__42742),
            .I(N__42736));
    Odrv4 I__10035 (
            .O(N__42739),
            .I(n10148));
    LocalMux I__10034 (
            .O(N__42736),
            .I(n10148));
    CascadeMux I__10033 (
            .O(N__42731),
            .I(N__42728));
    InMux I__10032 (
            .O(N__42728),
            .I(N__42723));
    InMux I__10031 (
            .O(N__42727),
            .I(N__42718));
    InMux I__10030 (
            .O(N__42726),
            .I(N__42718));
    LocalMux I__10029 (
            .O(N__42723),
            .I(N__42713));
    LocalMux I__10028 (
            .O(N__42718),
            .I(N__42713));
    Span4Mux_h I__10027 (
            .O(N__42713),
            .I(N__42710));
    Odrv4 I__10026 (
            .O(N__42710),
            .I(n7));
    InMux I__10025 (
            .O(N__42707),
            .I(N__42703));
    InMux I__10024 (
            .O(N__42706),
            .I(N__42700));
    LocalMux I__10023 (
            .O(N__42703),
            .I(comm_state_3_N_418_1));
    LocalMux I__10022 (
            .O(N__42700),
            .I(comm_state_3_N_418_1));
    CascadeMux I__10021 (
            .O(N__42695),
            .I(n15711_cascade_));
    InMux I__10020 (
            .O(N__42692),
            .I(N__42689));
    LocalMux I__10019 (
            .O(N__42689),
            .I(n8_adj_1193));
    InMux I__10018 (
            .O(N__42686),
            .I(N__42683));
    LocalMux I__10017 (
            .O(N__42683),
            .I(N__42680));
    Span4Mux_h I__10016 (
            .O(N__42680),
            .I(N__42677));
    Odrv4 I__10015 (
            .O(N__42677),
            .I(buf_data2_9));
    CascadeMux I__10014 (
            .O(N__42674),
            .I(N__42671));
    InMux I__10013 (
            .O(N__42671),
            .I(N__42667));
    InMux I__10012 (
            .O(N__42670),
            .I(N__42664));
    LocalMux I__10011 (
            .O(N__42667),
            .I(N__42661));
    LocalMux I__10010 (
            .O(N__42664),
            .I(N__42658));
    Span4Mux_v I__10009 (
            .O(N__42661),
            .I(N__42653));
    Span4Mux_h I__10008 (
            .O(N__42658),
            .I(N__42653));
    Span4Mux_v I__10007 (
            .O(N__42653),
            .I(N__42649));
    CascadeMux I__10006 (
            .O(N__42652),
            .I(N__42646));
    Sp12to4 I__10005 (
            .O(N__42649),
            .I(N__42643));
    InMux I__10004 (
            .O(N__42646),
            .I(N__42640));
    Span12Mux_h I__10003 (
            .O(N__42643),
            .I(N__42637));
    LocalMux I__10002 (
            .O(N__42640),
            .I(buf_adcdata4_9));
    Odrv12 I__10001 (
            .O(N__42637),
            .I(buf_adcdata4_9));
    InMux I__10000 (
            .O(N__42632),
            .I(N__42629));
    LocalMux I__9999 (
            .O(N__42629),
            .I(N__42626));
    Span12Mux_h I__9998 (
            .O(N__42626),
            .I(N__42623));
    Odrv12 I__9997 (
            .O(N__42623),
            .I(n4063));
    InMux I__9996 (
            .O(N__42620),
            .I(N__42617));
    LocalMux I__9995 (
            .O(N__42617),
            .I(N__42613));
    InMux I__9994 (
            .O(N__42616),
            .I(N__42610));
    Span4Mux_h I__9993 (
            .O(N__42613),
            .I(N__42607));
    LocalMux I__9992 (
            .O(N__42610),
            .I(buf_adcdata2_11));
    Odrv4 I__9991 (
            .O(N__42607),
            .I(buf_adcdata2_11));
    InMux I__9990 (
            .O(N__42602),
            .I(N__42598));
    InMux I__9989 (
            .O(N__42601),
            .I(N__42595));
    LocalMux I__9988 (
            .O(N__42598),
            .I(N__42592));
    LocalMux I__9987 (
            .O(N__42595),
            .I(N__42589));
    Span4Mux_v I__9986 (
            .O(N__42592),
            .I(N__42586));
    Odrv4 I__9985 (
            .O(N__42589),
            .I(n8_adj_1219));
    Odrv4 I__9984 (
            .O(N__42586),
            .I(n8_adj_1219));
    InMux I__9983 (
            .O(N__42581),
            .I(N__42577));
    InMux I__9982 (
            .O(N__42580),
            .I(N__42574));
    LocalMux I__9981 (
            .O(N__42577),
            .I(N__42571));
    LocalMux I__9980 (
            .O(N__42574),
            .I(N__42566));
    Span4Mux_h I__9979 (
            .O(N__42571),
            .I(N__42566));
    Odrv4 I__9978 (
            .O(N__42566),
            .I(n7_adj_1218));
    CascadeMux I__9977 (
            .O(N__42563),
            .I(N__42560));
    CascadeBuf I__9976 (
            .O(N__42560),
            .I(N__42557));
    CascadeMux I__9975 (
            .O(N__42557),
            .I(N__42554));
    CascadeBuf I__9974 (
            .O(N__42554),
            .I(N__42551));
    CascadeMux I__9973 (
            .O(N__42551),
            .I(N__42548));
    CascadeBuf I__9972 (
            .O(N__42548),
            .I(N__42545));
    CascadeMux I__9971 (
            .O(N__42545),
            .I(N__42542));
    CascadeBuf I__9970 (
            .O(N__42542),
            .I(N__42539));
    CascadeMux I__9969 (
            .O(N__42539),
            .I(N__42536));
    CascadeBuf I__9968 (
            .O(N__42536),
            .I(N__42533));
    CascadeMux I__9967 (
            .O(N__42533),
            .I(N__42530));
    CascadeBuf I__9966 (
            .O(N__42530),
            .I(N__42527));
    CascadeMux I__9965 (
            .O(N__42527),
            .I(N__42524));
    CascadeBuf I__9964 (
            .O(N__42524),
            .I(N__42520));
    CascadeMux I__9963 (
            .O(N__42523),
            .I(N__42517));
    CascadeMux I__9962 (
            .O(N__42520),
            .I(N__42514));
    CascadeBuf I__9961 (
            .O(N__42517),
            .I(N__42511));
    CascadeBuf I__9960 (
            .O(N__42514),
            .I(N__42508));
    CascadeMux I__9959 (
            .O(N__42511),
            .I(N__42505));
    CascadeMux I__9958 (
            .O(N__42508),
            .I(N__42502));
    InMux I__9957 (
            .O(N__42505),
            .I(N__42499));
    CascadeBuf I__9956 (
            .O(N__42502),
            .I(N__42496));
    LocalMux I__9955 (
            .O(N__42499),
            .I(N__42493));
    CascadeMux I__9954 (
            .O(N__42496),
            .I(N__42490));
    Span12Mux_h I__9953 (
            .O(N__42493),
            .I(N__42487));
    InMux I__9952 (
            .O(N__42490),
            .I(N__42484));
    Span12Mux_v I__9951 (
            .O(N__42487),
            .I(N__42481));
    LocalMux I__9950 (
            .O(N__42484),
            .I(N__42478));
    Odrv12 I__9949 (
            .O(N__42481),
            .I(data_index_9_N_258_8));
    Odrv4 I__9948 (
            .O(N__42478),
            .I(data_index_9_N_258_8));
    InMux I__9947 (
            .O(N__42473),
            .I(N__42470));
    LocalMux I__9946 (
            .O(N__42470),
            .I(\comm_spi.n10456 ));
    ClkMux I__9945 (
            .O(N__42467),
            .I(N__42456));
    ClkMux I__9944 (
            .O(N__42466),
            .I(N__42452));
    ClkMux I__9943 (
            .O(N__42465),
            .I(N__42449));
    ClkMux I__9942 (
            .O(N__42464),
            .I(N__42444));
    ClkMux I__9941 (
            .O(N__42463),
            .I(N__42441));
    ClkMux I__9940 (
            .O(N__42462),
            .I(N__42435));
    ClkMux I__9939 (
            .O(N__42461),
            .I(N__42432));
    ClkMux I__9938 (
            .O(N__42460),
            .I(N__42428));
    ClkMux I__9937 (
            .O(N__42459),
            .I(N__42425));
    LocalMux I__9936 (
            .O(N__42456),
            .I(N__42421));
    ClkMux I__9935 (
            .O(N__42455),
            .I(N__42417));
    LocalMux I__9934 (
            .O(N__42452),
            .I(N__42414));
    LocalMux I__9933 (
            .O(N__42449),
            .I(N__42411));
    ClkMux I__9932 (
            .O(N__42448),
            .I(N__42408));
    ClkMux I__9931 (
            .O(N__42447),
            .I(N__42405));
    LocalMux I__9930 (
            .O(N__42444),
            .I(N__42399));
    LocalMux I__9929 (
            .O(N__42441),
            .I(N__42399));
    ClkMux I__9928 (
            .O(N__42440),
            .I(N__42396));
    ClkMux I__9927 (
            .O(N__42439),
            .I(N__42393));
    ClkMux I__9926 (
            .O(N__42438),
            .I(N__42390));
    LocalMux I__9925 (
            .O(N__42435),
            .I(N__42385));
    LocalMux I__9924 (
            .O(N__42432),
            .I(N__42385));
    ClkMux I__9923 (
            .O(N__42431),
            .I(N__42382));
    LocalMux I__9922 (
            .O(N__42428),
            .I(N__42376));
    LocalMux I__9921 (
            .O(N__42425),
            .I(N__42376));
    ClkMux I__9920 (
            .O(N__42424),
            .I(N__42372));
    Span4Mux_h I__9919 (
            .O(N__42421),
            .I(N__42368));
    ClkMux I__9918 (
            .O(N__42420),
            .I(N__42365));
    LocalMux I__9917 (
            .O(N__42417),
            .I(N__42362));
    Span4Mux_h I__9916 (
            .O(N__42414),
            .I(N__42353));
    Span4Mux_h I__9915 (
            .O(N__42411),
            .I(N__42353));
    LocalMux I__9914 (
            .O(N__42408),
            .I(N__42353));
    LocalMux I__9913 (
            .O(N__42405),
            .I(N__42353));
    ClkMux I__9912 (
            .O(N__42404),
            .I(N__42350));
    Span4Mux_v I__9911 (
            .O(N__42399),
            .I(N__42345));
    LocalMux I__9910 (
            .O(N__42396),
            .I(N__42345));
    LocalMux I__9909 (
            .O(N__42393),
            .I(N__42342));
    LocalMux I__9908 (
            .O(N__42390),
            .I(N__42339));
    Span4Mux_v I__9907 (
            .O(N__42385),
            .I(N__42334));
    LocalMux I__9906 (
            .O(N__42382),
            .I(N__42334));
    ClkMux I__9905 (
            .O(N__42381),
            .I(N__42331));
    Span4Mux_v I__9904 (
            .O(N__42376),
            .I(N__42328));
    ClkMux I__9903 (
            .O(N__42375),
            .I(N__42325));
    LocalMux I__9902 (
            .O(N__42372),
            .I(N__42322));
    ClkMux I__9901 (
            .O(N__42371),
            .I(N__42319));
    Span4Mux_h I__9900 (
            .O(N__42368),
            .I(N__42314));
    LocalMux I__9899 (
            .O(N__42365),
            .I(N__42314));
    Span4Mux_h I__9898 (
            .O(N__42362),
            .I(N__42307));
    Span4Mux_h I__9897 (
            .O(N__42353),
            .I(N__42307));
    LocalMux I__9896 (
            .O(N__42350),
            .I(N__42307));
    Span4Mux_v I__9895 (
            .O(N__42345),
            .I(N__42302));
    Span4Mux_v I__9894 (
            .O(N__42342),
            .I(N__42302));
    Span4Mux_h I__9893 (
            .O(N__42339),
            .I(N__42299));
    Span4Mux_h I__9892 (
            .O(N__42334),
            .I(N__42294));
    LocalMux I__9891 (
            .O(N__42331),
            .I(N__42294));
    Span4Mux_h I__9890 (
            .O(N__42328),
            .I(N__42285));
    LocalMux I__9889 (
            .O(N__42325),
            .I(N__42285));
    Span4Mux_v I__9888 (
            .O(N__42322),
            .I(N__42285));
    LocalMux I__9887 (
            .O(N__42319),
            .I(N__42285));
    Span4Mux_h I__9886 (
            .O(N__42314),
            .I(N__42280));
    Span4Mux_h I__9885 (
            .O(N__42307),
            .I(N__42280));
    Span4Mux_h I__9884 (
            .O(N__42302),
            .I(N__42277));
    Span4Mux_v I__9883 (
            .O(N__42299),
            .I(N__42272));
    Span4Mux_h I__9882 (
            .O(N__42294),
            .I(N__42272));
    Span4Mux_h I__9881 (
            .O(N__42285),
            .I(N__42269));
    Odrv4 I__9880 (
            .O(N__42280),
            .I(\comm_spi.iclk ));
    Odrv4 I__9879 (
            .O(N__42277),
            .I(\comm_spi.iclk ));
    Odrv4 I__9878 (
            .O(N__42272),
            .I(\comm_spi.iclk ));
    Odrv4 I__9877 (
            .O(N__42269),
            .I(\comm_spi.iclk ));
    InMux I__9876 (
            .O(N__42260),
            .I(N__42257));
    LocalMux I__9875 (
            .O(N__42257),
            .I(N__42254));
    Span4Mux_v I__9874 (
            .O(N__42254),
            .I(N__42249));
    InMux I__9873 (
            .O(N__42253),
            .I(N__42246));
    InMux I__9872 (
            .O(N__42252),
            .I(N__42243));
    Odrv4 I__9871 (
            .O(N__42249),
            .I(\comm_spi.n16893 ));
    LocalMux I__9870 (
            .O(N__42246),
            .I(\comm_spi.n16893 ));
    LocalMux I__9869 (
            .O(N__42243),
            .I(\comm_spi.n16893 ));
    InMux I__9868 (
            .O(N__42236),
            .I(N__42233));
    LocalMux I__9867 (
            .O(N__42233),
            .I(N__42229));
    InMux I__9866 (
            .O(N__42232),
            .I(N__42225));
    Span4Mux_v I__9865 (
            .O(N__42229),
            .I(N__42222));
    InMux I__9864 (
            .O(N__42228),
            .I(N__42219));
    LocalMux I__9863 (
            .O(N__42225),
            .I(N__42216));
    Odrv4 I__9862 (
            .O(N__42222),
            .I(\comm_spi.n10441 ));
    LocalMux I__9861 (
            .O(N__42219),
            .I(\comm_spi.n10441 ));
    Odrv4 I__9860 (
            .O(N__42216),
            .I(\comm_spi.n10441 ));
    CascadeMux I__9859 (
            .O(N__42209),
            .I(\comm_spi.n16893_cascade_ ));
    CascadeMux I__9858 (
            .O(N__42206),
            .I(\comm_spi.imosi_cascade_ ));
    SRMux I__9857 (
            .O(N__42203),
            .I(N__42200));
    LocalMux I__9856 (
            .O(N__42200),
            .I(N__42197));
    Span4Mux_h I__9855 (
            .O(N__42197),
            .I(N__42194));
    Odrv4 I__9854 (
            .O(N__42194),
            .I(\comm_spi.DOUT_7__N_785 ));
    InMux I__9853 (
            .O(N__42191),
            .I(N__42188));
    LocalMux I__9852 (
            .O(N__42188),
            .I(N__42184));
    CascadeMux I__9851 (
            .O(N__42187),
            .I(N__42181));
    Span4Mux_v I__9850 (
            .O(N__42184),
            .I(N__42178));
    InMux I__9849 (
            .O(N__42181),
            .I(N__42174));
    Span4Mux_h I__9848 (
            .O(N__42178),
            .I(N__42171));
    InMux I__9847 (
            .O(N__42177),
            .I(N__42168));
    LocalMux I__9846 (
            .O(N__42174),
            .I(acadc_skipCount_1));
    Odrv4 I__9845 (
            .O(N__42171),
            .I(acadc_skipCount_1));
    LocalMux I__9844 (
            .O(N__42168),
            .I(acadc_skipCount_1));
    InMux I__9843 (
            .O(N__42161),
            .I(N__42156));
    InMux I__9842 (
            .O(N__42160),
            .I(N__42153));
    InMux I__9841 (
            .O(N__42159),
            .I(N__42150));
    LocalMux I__9840 (
            .O(N__42156),
            .I(req_data_cnt_1));
    LocalMux I__9839 (
            .O(N__42153),
            .I(req_data_cnt_1));
    LocalMux I__9838 (
            .O(N__42150),
            .I(req_data_cnt_1));
    CascadeMux I__9837 (
            .O(N__42143),
            .I(n4220_cascade_));
    CascadeMux I__9836 (
            .O(N__42140),
            .I(n4253_cascade_));
    InMux I__9835 (
            .O(N__42137),
            .I(N__42134));
    LocalMux I__9834 (
            .O(N__42134),
            .I(N__42131));
    Span12Mux_v I__9833 (
            .O(N__42131),
            .I(N__42128));
    Odrv12 I__9832 (
            .O(N__42128),
            .I(n4263));
    InMux I__9831 (
            .O(N__42125),
            .I(N__42121));
    CascadeMux I__9830 (
            .O(N__42124),
            .I(N__42117));
    LocalMux I__9829 (
            .O(N__42121),
            .I(N__42114));
    InMux I__9828 (
            .O(N__42120),
            .I(N__42111));
    InMux I__9827 (
            .O(N__42117),
            .I(N__42108));
    Span4Mux_v I__9826 (
            .O(N__42114),
            .I(N__42105));
    LocalMux I__9825 (
            .O(N__42111),
            .I(N__42102));
    LocalMux I__9824 (
            .O(N__42108),
            .I(buf_dds_1));
    Odrv4 I__9823 (
            .O(N__42105),
            .I(buf_dds_1));
    Odrv12 I__9822 (
            .O(N__42102),
            .I(buf_dds_1));
    InMux I__9821 (
            .O(N__42095),
            .I(N__42092));
    LocalMux I__9820 (
            .O(N__42092),
            .I(N__42089));
    Span4Mux_v I__9819 (
            .O(N__42089),
            .I(N__42084));
    InMux I__9818 (
            .O(N__42088),
            .I(N__42081));
    InMux I__9817 (
            .O(N__42087),
            .I(N__42078));
    Sp12to4 I__9816 (
            .O(N__42084),
            .I(N__42073));
    LocalMux I__9815 (
            .O(N__42081),
            .I(N__42073));
    LocalMux I__9814 (
            .O(N__42078),
            .I(buf_adcdata3_9));
    Odrv12 I__9813 (
            .O(N__42073),
            .I(buf_adcdata3_9));
    InMux I__9812 (
            .O(N__42068),
            .I(N__42065));
    LocalMux I__9811 (
            .O(N__42065),
            .I(n4208));
    CascadeMux I__9810 (
            .O(N__42062),
            .I(N__42059));
    InMux I__9809 (
            .O(N__42059),
            .I(N__42056));
    LocalMux I__9808 (
            .O(N__42056),
            .I(N__42053));
    Span4Mux_h I__9807 (
            .O(N__42053),
            .I(N__42050));
    Odrv4 I__9806 (
            .O(N__42050),
            .I(buf_data1_9));
    InMux I__9805 (
            .O(N__42047),
            .I(N__42044));
    LocalMux I__9804 (
            .O(N__42044),
            .I(n4196));
    InMux I__9803 (
            .O(N__42041),
            .I(N__42038));
    LocalMux I__9802 (
            .O(N__42038),
            .I(n4233));
    InMux I__9801 (
            .O(N__42035),
            .I(N__42032));
    LocalMux I__9800 (
            .O(N__42032),
            .I(N__42028));
    InMux I__9799 (
            .O(N__42031),
            .I(N__42025));
    Span4Mux_v I__9798 (
            .O(N__42028),
            .I(N__42022));
    LocalMux I__9797 (
            .O(N__42025),
            .I(data_idxvec_3));
    Odrv4 I__9796 (
            .O(N__42022),
            .I(data_idxvec_3));
    InMux I__9795 (
            .O(N__42017),
            .I(N__42012));
    InMux I__9794 (
            .O(N__42016),
            .I(N__42009));
    InMux I__9793 (
            .O(N__42015),
            .I(N__42006));
    LocalMux I__9792 (
            .O(N__42012),
            .I(N__42003));
    LocalMux I__9791 (
            .O(N__42009),
            .I(data_cntvec_3));
    LocalMux I__9790 (
            .O(N__42006),
            .I(data_cntvec_3));
    Odrv4 I__9789 (
            .O(N__42003),
            .I(data_cntvec_3));
    InMux I__9788 (
            .O(N__41996),
            .I(N__41993));
    LocalMux I__9787 (
            .O(N__41993),
            .I(N__41990));
    Span4Mux_v I__9786 (
            .O(N__41990),
            .I(N__41987));
    Span4Mux_h I__9785 (
            .O(N__41987),
            .I(N__41984));
    Odrv4 I__9784 (
            .O(N__41984),
            .I(buf_data1_11));
    CascadeMux I__9783 (
            .O(N__41981),
            .I(n4194_cascade_));
    InMux I__9782 (
            .O(N__41978),
            .I(N__41975));
    LocalMux I__9781 (
            .O(N__41975),
            .I(n4218));
    CascadeMux I__9780 (
            .O(N__41972),
            .I(n4231_cascade_));
    InMux I__9779 (
            .O(N__41969),
            .I(N__41966));
    LocalMux I__9778 (
            .O(N__41966),
            .I(N__41963));
    Odrv4 I__9777 (
            .O(N__41963),
            .I(n4206));
    CascadeMux I__9776 (
            .O(N__41960),
            .I(n4251_cascade_));
    CascadeMux I__9775 (
            .O(N__41957),
            .I(N__41953));
    CascadeMux I__9774 (
            .O(N__41956),
            .I(N__41950));
    InMux I__9773 (
            .O(N__41953),
            .I(N__41944));
    InMux I__9772 (
            .O(N__41950),
            .I(N__41944));
    InMux I__9771 (
            .O(N__41949),
            .I(N__41941));
    LocalMux I__9770 (
            .O(N__41944),
            .I(cmd_rdadctmp_21_adj_1091));
    LocalMux I__9769 (
            .O(N__41941),
            .I(cmd_rdadctmp_21_adj_1091));
    InMux I__9768 (
            .O(N__41936),
            .I(N__41932));
    InMux I__9767 (
            .O(N__41935),
            .I(N__41928));
    LocalMux I__9766 (
            .O(N__41932),
            .I(N__41925));
    InMux I__9765 (
            .O(N__41931),
            .I(N__41922));
    LocalMux I__9764 (
            .O(N__41928),
            .I(N__41919));
    Span4Mux_v I__9763 (
            .O(N__41925),
            .I(N__41914));
    LocalMux I__9762 (
            .O(N__41922),
            .I(N__41914));
    Span4Mux_v I__9761 (
            .O(N__41919),
            .I(N__41910));
    Span4Mux_h I__9760 (
            .O(N__41914),
            .I(N__41907));
    InMux I__9759 (
            .O(N__41913),
            .I(N__41904));
    Odrv4 I__9758 (
            .O(N__41910),
            .I(n4_adj_1041));
    Odrv4 I__9757 (
            .O(N__41907),
            .I(n4_adj_1041));
    LocalMux I__9756 (
            .O(N__41904),
            .I(n4_adj_1041));
    CascadeMux I__9755 (
            .O(N__41897),
            .I(N__41891));
    InMux I__9754 (
            .O(N__41896),
            .I(N__41888));
    InMux I__9753 (
            .O(N__41895),
            .I(N__41883));
    InMux I__9752 (
            .O(N__41894),
            .I(N__41880));
    InMux I__9751 (
            .O(N__41891),
            .I(N__41877));
    LocalMux I__9750 (
            .O(N__41888),
            .I(N__41874));
    InMux I__9749 (
            .O(N__41887),
            .I(N__41869));
    InMux I__9748 (
            .O(N__41886),
            .I(N__41869));
    LocalMux I__9747 (
            .O(N__41883),
            .I(N__41864));
    LocalMux I__9746 (
            .O(N__41880),
            .I(N__41864));
    LocalMux I__9745 (
            .O(N__41877),
            .I(N__41860));
    Span4Mux_v I__9744 (
            .O(N__41874),
            .I(N__41855));
    LocalMux I__9743 (
            .O(N__41869),
            .I(N__41855));
    Span4Mux_v I__9742 (
            .O(N__41864),
            .I(N__41852));
    InMux I__9741 (
            .O(N__41863),
            .I(N__41849));
    Span4Mux_h I__9740 (
            .O(N__41860),
            .I(N__41846));
    Span4Mux_h I__9739 (
            .O(N__41855),
            .I(N__41843));
    Sp12to4 I__9738 (
            .O(N__41852),
            .I(N__41838));
    LocalMux I__9737 (
            .O(N__41849),
            .I(N__41838));
    Span4Mux_v I__9736 (
            .O(N__41846),
            .I(N__41835));
    Odrv4 I__9735 (
            .O(N__41843),
            .I(comm_buf_0_6));
    Odrv12 I__9734 (
            .O(N__41838),
            .I(comm_buf_0_6));
    Odrv4 I__9733 (
            .O(N__41835),
            .I(comm_buf_0_6));
    CascadeMux I__9732 (
            .O(N__41828),
            .I(N__41815));
    InMux I__9731 (
            .O(N__41827),
            .I(N__41812));
    InMux I__9730 (
            .O(N__41826),
            .I(N__41807));
    InMux I__9729 (
            .O(N__41825),
            .I(N__41807));
    InMux I__9728 (
            .O(N__41824),
            .I(N__41804));
    InMux I__9727 (
            .O(N__41823),
            .I(N__41801));
    InMux I__9726 (
            .O(N__41822),
            .I(N__41798));
    InMux I__9725 (
            .O(N__41821),
            .I(N__41791));
    InMux I__9724 (
            .O(N__41820),
            .I(N__41791));
    InMux I__9723 (
            .O(N__41819),
            .I(N__41791));
    InMux I__9722 (
            .O(N__41818),
            .I(N__41786));
    InMux I__9721 (
            .O(N__41815),
            .I(N__41782));
    LocalMux I__9720 (
            .O(N__41812),
            .I(N__41779));
    LocalMux I__9719 (
            .O(N__41807),
            .I(N__41776));
    LocalMux I__9718 (
            .O(N__41804),
            .I(N__41773));
    LocalMux I__9717 (
            .O(N__41801),
            .I(N__41766));
    LocalMux I__9716 (
            .O(N__41798),
            .I(N__41766));
    LocalMux I__9715 (
            .O(N__41791),
            .I(N__41766));
    InMux I__9714 (
            .O(N__41790),
            .I(N__41761));
    InMux I__9713 (
            .O(N__41789),
            .I(N__41761));
    LocalMux I__9712 (
            .O(N__41786),
            .I(N__41758));
    InMux I__9711 (
            .O(N__41785),
            .I(N__41753));
    LocalMux I__9710 (
            .O(N__41782),
            .I(N__41746));
    Span4Mux_v I__9709 (
            .O(N__41779),
            .I(N__41746));
    Span4Mux_h I__9708 (
            .O(N__41776),
            .I(N__41746));
    Span4Mux_h I__9707 (
            .O(N__41773),
            .I(N__41739));
    Span4Mux_v I__9706 (
            .O(N__41766),
            .I(N__41739));
    LocalMux I__9705 (
            .O(N__41761),
            .I(N__41739));
    Span4Mux_h I__9704 (
            .O(N__41758),
            .I(N__41736));
    InMux I__9703 (
            .O(N__41757),
            .I(N__41733));
    InMux I__9702 (
            .O(N__41756),
            .I(N__41730));
    LocalMux I__9701 (
            .O(N__41753),
            .I(N__41727));
    Span4Mux_h I__9700 (
            .O(N__41746),
            .I(N__41724));
    Span4Mux_h I__9699 (
            .O(N__41739),
            .I(N__41719));
    Span4Mux_h I__9698 (
            .O(N__41736),
            .I(N__41719));
    LocalMux I__9697 (
            .O(N__41733),
            .I(n8250));
    LocalMux I__9696 (
            .O(N__41730),
            .I(n8250));
    Odrv12 I__9695 (
            .O(N__41727),
            .I(n8250));
    Odrv4 I__9694 (
            .O(N__41724),
            .I(n8250));
    Odrv4 I__9693 (
            .O(N__41719),
            .I(n8250));
    InMux I__9692 (
            .O(N__41708),
            .I(N__41705));
    LocalMux I__9691 (
            .O(N__41705),
            .I(N__41701));
    InMux I__9690 (
            .O(N__41704),
            .I(N__41698));
    Span4Mux_h I__9689 (
            .O(N__41701),
            .I(N__41694));
    LocalMux I__9688 (
            .O(N__41698),
            .I(N__41691));
    InMux I__9687 (
            .O(N__41697),
            .I(N__41688));
    Span4Mux_h I__9686 (
            .O(N__41694),
            .I(N__41685));
    Span4Mux_v I__9685 (
            .O(N__41691),
            .I(N__41682));
    LocalMux I__9684 (
            .O(N__41688),
            .I(acadc_skipCount_14));
    Odrv4 I__9683 (
            .O(N__41685),
            .I(acadc_skipCount_14));
    Odrv4 I__9682 (
            .O(N__41682),
            .I(acadc_skipCount_14));
    CascadeMux I__9681 (
            .O(N__41675),
            .I(N__41671));
    CascadeMux I__9680 (
            .O(N__41674),
            .I(N__41668));
    InMux I__9679 (
            .O(N__41671),
            .I(N__41665));
    InMux I__9678 (
            .O(N__41668),
            .I(N__41662));
    LocalMux I__9677 (
            .O(N__41665),
            .I(data_idxvec_15));
    LocalMux I__9676 (
            .O(N__41662),
            .I(data_idxvec_15));
    CascadeMux I__9675 (
            .O(N__41657),
            .I(N__41653));
    InMux I__9674 (
            .O(N__41656),
            .I(N__41649));
    InMux I__9673 (
            .O(N__41653),
            .I(N__41646));
    InMux I__9672 (
            .O(N__41652),
            .I(N__41643));
    LocalMux I__9671 (
            .O(N__41649),
            .I(N__41640));
    LocalMux I__9670 (
            .O(N__41646),
            .I(acadc_skipCount_15));
    LocalMux I__9669 (
            .O(N__41643),
            .I(acadc_skipCount_15));
    Odrv4 I__9668 (
            .O(N__41640),
            .I(acadc_skipCount_15));
    CascadeMux I__9667 (
            .O(N__41633),
            .I(N__41630));
    InMux I__9666 (
            .O(N__41630),
            .I(N__41627));
    LocalMux I__9665 (
            .O(N__41627),
            .I(N__41624));
    Span4Mux_v I__9664 (
            .O(N__41624),
            .I(N__41621));
    Span4Mux_h I__9663 (
            .O(N__41621),
            .I(N__41618));
    Odrv4 I__9662 (
            .O(N__41618),
            .I(n15468));
    InMux I__9661 (
            .O(N__41615),
            .I(N__41612));
    LocalMux I__9660 (
            .O(N__41612),
            .I(N__41609));
    Odrv4 I__9659 (
            .O(N__41609),
            .I(n4217));
    InMux I__9658 (
            .O(N__41606),
            .I(N__41603));
    LocalMux I__9657 (
            .O(N__41603),
            .I(n4230));
    InMux I__9656 (
            .O(N__41600),
            .I(N__41597));
    LocalMux I__9655 (
            .O(N__41597),
            .I(N__41594));
    Span4Mux_h I__9654 (
            .O(N__41594),
            .I(N__41591));
    Span4Mux_v I__9653 (
            .O(N__41591),
            .I(N__41588));
    Odrv4 I__9652 (
            .O(N__41588),
            .I(n4250));
    InMux I__9651 (
            .O(N__41585),
            .I(N__41582));
    LocalMux I__9650 (
            .O(N__41582),
            .I(N__41579));
    Span4Mux_v I__9649 (
            .O(N__41579),
            .I(N__41575));
    InMux I__9648 (
            .O(N__41578),
            .I(N__41571));
    Span4Mux_h I__9647 (
            .O(N__41575),
            .I(N__41568));
    InMux I__9646 (
            .O(N__41574),
            .I(N__41565));
    LocalMux I__9645 (
            .O(N__41571),
            .I(cmd_rdadctmp_22_adj_1090));
    Odrv4 I__9644 (
            .O(N__41568),
            .I(cmd_rdadctmp_22_adj_1090));
    LocalMux I__9643 (
            .O(N__41565),
            .I(cmd_rdadctmp_22_adj_1090));
    InMux I__9642 (
            .O(N__41558),
            .I(N__41554));
    InMux I__9641 (
            .O(N__41557),
            .I(N__41551));
    LocalMux I__9640 (
            .O(N__41554),
            .I(N__41547));
    LocalMux I__9639 (
            .O(N__41551),
            .I(N__41544));
    InMux I__9638 (
            .O(N__41550),
            .I(N__41541));
    Span4Mux_v I__9637 (
            .O(N__41547),
            .I(N__41538));
    Span4Mux_v I__9636 (
            .O(N__41544),
            .I(N__41535));
    LocalMux I__9635 (
            .O(N__41541),
            .I(buf_adcdata3_14));
    Odrv4 I__9634 (
            .O(N__41538),
            .I(buf_adcdata3_14));
    Odrv4 I__9633 (
            .O(N__41535),
            .I(buf_adcdata3_14));
    CascadeMux I__9632 (
            .O(N__41528),
            .I(N__41521));
    CascadeMux I__9631 (
            .O(N__41527),
            .I(N__41515));
    CascadeMux I__9630 (
            .O(N__41526),
            .I(N__41512));
    InMux I__9629 (
            .O(N__41525),
            .I(N__41507));
    InMux I__9628 (
            .O(N__41524),
            .I(N__41502));
    InMux I__9627 (
            .O(N__41521),
            .I(N__41499));
    CascadeMux I__9626 (
            .O(N__41520),
            .I(N__41494));
    CascadeMux I__9625 (
            .O(N__41519),
            .I(N__41491));
    CascadeMux I__9624 (
            .O(N__41518),
            .I(N__41488));
    InMux I__9623 (
            .O(N__41515),
            .I(N__41485));
    InMux I__9622 (
            .O(N__41512),
            .I(N__41482));
    CascadeMux I__9621 (
            .O(N__41511),
            .I(N__41479));
    InMux I__9620 (
            .O(N__41510),
            .I(N__41476));
    LocalMux I__9619 (
            .O(N__41507),
            .I(N__41473));
    CascadeMux I__9618 (
            .O(N__41506),
            .I(N__41470));
    CascadeMux I__9617 (
            .O(N__41505),
            .I(N__41467));
    LocalMux I__9616 (
            .O(N__41502),
            .I(N__41464));
    LocalMux I__9615 (
            .O(N__41499),
            .I(N__41461));
    InMux I__9614 (
            .O(N__41498),
            .I(N__41454));
    InMux I__9613 (
            .O(N__41497),
            .I(N__41454));
    InMux I__9612 (
            .O(N__41494),
            .I(N__41454));
    InMux I__9611 (
            .O(N__41491),
            .I(N__41451));
    InMux I__9610 (
            .O(N__41488),
            .I(N__41448));
    LocalMux I__9609 (
            .O(N__41485),
            .I(N__41443));
    LocalMux I__9608 (
            .O(N__41482),
            .I(N__41443));
    InMux I__9607 (
            .O(N__41479),
            .I(N__41440));
    LocalMux I__9606 (
            .O(N__41476),
            .I(N__41437));
    Span4Mux_h I__9605 (
            .O(N__41473),
            .I(N__41434));
    InMux I__9604 (
            .O(N__41470),
            .I(N__41429));
    InMux I__9603 (
            .O(N__41467),
            .I(N__41429));
    Span4Mux_v I__9602 (
            .O(N__41464),
            .I(N__41426));
    Span4Mux_v I__9601 (
            .O(N__41461),
            .I(N__41423));
    LocalMux I__9600 (
            .O(N__41454),
            .I(N__41420));
    LocalMux I__9599 (
            .O(N__41451),
            .I(N__41417));
    LocalMux I__9598 (
            .O(N__41448),
            .I(N__41404));
    Span4Mux_h I__9597 (
            .O(N__41443),
            .I(N__41404));
    LocalMux I__9596 (
            .O(N__41440),
            .I(N__41404));
    Span4Mux_v I__9595 (
            .O(N__41437),
            .I(N__41404));
    Span4Mux_h I__9594 (
            .O(N__41434),
            .I(N__41404));
    LocalMux I__9593 (
            .O(N__41429),
            .I(N__41404));
    Span4Mux_h I__9592 (
            .O(N__41426),
            .I(N__41399));
    Span4Mux_h I__9591 (
            .O(N__41423),
            .I(N__41399));
    Span4Mux_v I__9590 (
            .O(N__41420),
            .I(N__41396));
    Span4Mux_h I__9589 (
            .O(N__41417),
            .I(N__41391));
    Span4Mux_v I__9588 (
            .O(N__41404),
            .I(N__41391));
    Span4Mux_v I__9587 (
            .O(N__41399),
            .I(N__41388));
    Odrv4 I__9586 (
            .O(N__41396),
            .I(n1));
    Odrv4 I__9585 (
            .O(N__41391),
            .I(n1));
    Odrv4 I__9584 (
            .O(N__41388),
            .I(n1));
    CascadeMux I__9583 (
            .O(N__41381),
            .I(N__41375));
    InMux I__9582 (
            .O(N__41380),
            .I(N__41370));
    InMux I__9581 (
            .O(N__41379),
            .I(N__41365));
    InMux I__9580 (
            .O(N__41378),
            .I(N__41362));
    InMux I__9579 (
            .O(N__41375),
            .I(N__41357));
    InMux I__9578 (
            .O(N__41374),
            .I(N__41353));
    InMux I__9577 (
            .O(N__41373),
            .I(N__41350));
    LocalMux I__9576 (
            .O(N__41370),
            .I(N__41347));
    InMux I__9575 (
            .O(N__41369),
            .I(N__41343));
    InMux I__9574 (
            .O(N__41368),
            .I(N__41340));
    LocalMux I__9573 (
            .O(N__41365),
            .I(N__41337));
    LocalMux I__9572 (
            .O(N__41362),
            .I(N__41334));
    InMux I__9571 (
            .O(N__41361),
            .I(N__41329));
    InMux I__9570 (
            .O(N__41360),
            .I(N__41329));
    LocalMux I__9569 (
            .O(N__41357),
            .I(N__41326));
    InMux I__9568 (
            .O(N__41356),
            .I(N__41323));
    LocalMux I__9567 (
            .O(N__41353),
            .I(N__41320));
    LocalMux I__9566 (
            .O(N__41350),
            .I(N__41315));
    Span4Mux_h I__9565 (
            .O(N__41347),
            .I(N__41315));
    InMux I__9564 (
            .O(N__41346),
            .I(N__41309));
    LocalMux I__9563 (
            .O(N__41343),
            .I(N__41306));
    LocalMux I__9562 (
            .O(N__41340),
            .I(N__41301));
    Span4Mux_v I__9561 (
            .O(N__41337),
            .I(N__41301));
    Span4Mux_h I__9560 (
            .O(N__41334),
            .I(N__41288));
    LocalMux I__9559 (
            .O(N__41329),
            .I(N__41288));
    Span4Mux_h I__9558 (
            .O(N__41326),
            .I(N__41288));
    LocalMux I__9557 (
            .O(N__41323),
            .I(N__41288));
    Span4Mux_v I__9556 (
            .O(N__41320),
            .I(N__41288));
    Span4Mux_h I__9555 (
            .O(N__41315),
            .I(N__41288));
    InMux I__9554 (
            .O(N__41314),
            .I(N__41285));
    InMux I__9553 (
            .O(N__41313),
            .I(N__41280));
    InMux I__9552 (
            .O(N__41312),
            .I(N__41280));
    LocalMux I__9551 (
            .O(N__41309),
            .I(N__41277));
    Span4Mux_v I__9550 (
            .O(N__41306),
            .I(N__41272));
    Span4Mux_v I__9549 (
            .O(N__41301),
            .I(N__41272));
    Span4Mux_v I__9548 (
            .O(N__41288),
            .I(N__41269));
    LocalMux I__9547 (
            .O(N__41285),
            .I(n8525));
    LocalMux I__9546 (
            .O(N__41280),
            .I(n8525));
    Odrv4 I__9545 (
            .O(N__41277),
            .I(n8525));
    Odrv4 I__9544 (
            .O(N__41272),
            .I(n8525));
    Odrv4 I__9543 (
            .O(N__41269),
            .I(n8525));
    InMux I__9542 (
            .O(N__41258),
            .I(N__41254));
    InMux I__9541 (
            .O(N__41257),
            .I(N__41251));
    LocalMux I__9540 (
            .O(N__41254),
            .I(N__41248));
    LocalMux I__9539 (
            .O(N__41251),
            .I(N__41245));
    Span4Mux_v I__9538 (
            .O(N__41248),
            .I(N__41242));
    Span4Mux_h I__9537 (
            .O(N__41245),
            .I(N__41238));
    Span4Mux_h I__9536 (
            .O(N__41242),
            .I(N__41235));
    InMux I__9535 (
            .O(N__41241),
            .I(N__41232));
    Span4Mux_v I__9534 (
            .O(N__41238),
            .I(N__41227));
    Span4Mux_h I__9533 (
            .O(N__41235),
            .I(N__41227));
    LocalMux I__9532 (
            .O(N__41232),
            .I(buf_dds_11));
    Odrv4 I__9531 (
            .O(N__41227),
            .I(buf_dds_11));
    CascadeMux I__9530 (
            .O(N__41222),
            .I(N__41218));
    InMux I__9529 (
            .O(N__41221),
            .I(N__41215));
    InMux I__9528 (
            .O(N__41218),
            .I(N__41212));
    LocalMux I__9527 (
            .O(N__41215),
            .I(N__41207));
    LocalMux I__9526 (
            .O(N__41212),
            .I(N__41204));
    InMux I__9525 (
            .O(N__41211),
            .I(N__41201));
    InMux I__9524 (
            .O(N__41210),
            .I(N__41197));
    Span4Mux_h I__9523 (
            .O(N__41207),
            .I(N__41190));
    Span4Mux_v I__9522 (
            .O(N__41204),
            .I(N__41190));
    LocalMux I__9521 (
            .O(N__41201),
            .I(N__41190));
    InMux I__9520 (
            .O(N__41200),
            .I(N__41187));
    LocalMux I__9519 (
            .O(N__41197),
            .I(n12));
    Odrv4 I__9518 (
            .O(N__41190),
            .I(n12));
    LocalMux I__9517 (
            .O(N__41187),
            .I(n12));
    InMux I__9516 (
            .O(N__41180),
            .I(N__41177));
    LocalMux I__9515 (
            .O(N__41177),
            .I(N__41174));
    Odrv4 I__9514 (
            .O(N__41174),
            .I(n13_adj_1025));
    InMux I__9513 (
            .O(N__41171),
            .I(N__41161));
    InMux I__9512 (
            .O(N__41170),
            .I(N__41161));
    InMux I__9511 (
            .O(N__41169),
            .I(N__41158));
    InMux I__9510 (
            .O(N__41168),
            .I(N__41155));
    InMux I__9509 (
            .O(N__41167),
            .I(N__41152));
    InMux I__9508 (
            .O(N__41166),
            .I(N__41148));
    LocalMux I__9507 (
            .O(N__41161),
            .I(N__41139));
    LocalMux I__9506 (
            .O(N__41158),
            .I(N__41139));
    LocalMux I__9505 (
            .O(N__41155),
            .I(N__41139));
    LocalMux I__9504 (
            .O(N__41152),
            .I(N__41139));
    InMux I__9503 (
            .O(N__41151),
            .I(N__41136));
    LocalMux I__9502 (
            .O(N__41148),
            .I(N__41133));
    Span4Mux_v I__9501 (
            .O(N__41139),
            .I(N__41130));
    LocalMux I__9500 (
            .O(N__41136),
            .I(N__41127));
    Span12Mux_v I__9499 (
            .O(N__41133),
            .I(N__41123));
    Span4Mux_h I__9498 (
            .O(N__41130),
            .I(N__41120));
    Span4Mux_v I__9497 (
            .O(N__41127),
            .I(N__41117));
    InMux I__9496 (
            .O(N__41126),
            .I(N__41114));
    Odrv12 I__9495 (
            .O(N__41123),
            .I(n7511));
    Odrv4 I__9494 (
            .O(N__41120),
            .I(n7511));
    Odrv4 I__9493 (
            .O(N__41117),
            .I(n7511));
    LocalMux I__9492 (
            .O(N__41114),
            .I(n7511));
    InMux I__9491 (
            .O(N__41105),
            .I(N__41102));
    LocalMux I__9490 (
            .O(N__41102),
            .I(N__41098));
    InMux I__9489 (
            .O(N__41101),
            .I(N__41093));
    Span4Mux_v I__9488 (
            .O(N__41098),
            .I(N__41089));
    InMux I__9487 (
            .O(N__41097),
            .I(N__41086));
    InMux I__9486 (
            .O(N__41096),
            .I(N__41083));
    LocalMux I__9485 (
            .O(N__41093),
            .I(N__41080));
    InMux I__9484 (
            .O(N__41092),
            .I(N__41077));
    Span4Mux_h I__9483 (
            .O(N__41089),
            .I(N__41074));
    LocalMux I__9482 (
            .O(N__41086),
            .I(N__41071));
    LocalMux I__9481 (
            .O(N__41083),
            .I(N__41068));
    Span4Mux_v I__9480 (
            .O(N__41080),
            .I(N__41063));
    LocalMux I__9479 (
            .O(N__41077),
            .I(N__41063));
    Span4Mux_h I__9478 (
            .O(N__41074),
            .I(N__41060));
    Span4Mux_h I__9477 (
            .O(N__41071),
            .I(N__41055));
    Span4Mux_h I__9476 (
            .O(N__41068),
            .I(N__41055));
    Span4Mux_h I__9475 (
            .O(N__41063),
            .I(N__41052));
    Odrv4 I__9474 (
            .O(N__41060),
            .I(comm_buf_1_1));
    Odrv4 I__9473 (
            .O(N__41055),
            .I(comm_buf_1_1));
    Odrv4 I__9472 (
            .O(N__41052),
            .I(comm_buf_1_1));
    InMux I__9471 (
            .O(N__41045),
            .I(N__41041));
    InMux I__9470 (
            .O(N__41044),
            .I(N__41034));
    LocalMux I__9469 (
            .O(N__41041),
            .I(N__41031));
    InMux I__9468 (
            .O(N__41040),
            .I(N__41028));
    InMux I__9467 (
            .O(N__41039),
            .I(N__41021));
    InMux I__9466 (
            .O(N__41038),
            .I(N__41021));
    InMux I__9465 (
            .O(N__41037),
            .I(N__41021));
    LocalMux I__9464 (
            .O(N__41034),
            .I(N__41016));
    Span4Mux_v I__9463 (
            .O(N__41031),
            .I(N__41016));
    LocalMux I__9462 (
            .O(N__41028),
            .I(N__41013));
    LocalMux I__9461 (
            .O(N__41021),
            .I(N__41010));
    Odrv4 I__9460 (
            .O(N__41016),
            .I(eis_start));
    Odrv12 I__9459 (
            .O(N__41013),
            .I(eis_start));
    Odrv4 I__9458 (
            .O(N__41010),
            .I(eis_start));
    CascadeMux I__9457 (
            .O(N__41003),
            .I(N__40999));
    CascadeMux I__9456 (
            .O(N__41002),
            .I(N__40996));
    InMux I__9455 (
            .O(N__40999),
            .I(N__40993));
    InMux I__9454 (
            .O(N__40996),
            .I(N__40990));
    LocalMux I__9453 (
            .O(N__40993),
            .I(N__40985));
    LocalMux I__9452 (
            .O(N__40990),
            .I(N__40985));
    Odrv4 I__9451 (
            .O(N__40985),
            .I(data_idxvec_8));
    InMux I__9450 (
            .O(N__40982),
            .I(N__40979));
    LocalMux I__9449 (
            .O(N__40979),
            .I(N__40976));
    Span4Mux_h I__9448 (
            .O(N__40976),
            .I(N__40973));
    Odrv4 I__9447 (
            .O(N__40973),
            .I(n78_adj_1022));
    InMux I__9446 (
            .O(N__40970),
            .I(N__40966));
    InMux I__9445 (
            .O(N__40969),
            .I(N__40962));
    LocalMux I__9444 (
            .O(N__40966),
            .I(N__40959));
    InMux I__9443 (
            .O(N__40965),
            .I(N__40956));
    LocalMux I__9442 (
            .O(N__40962),
            .I(N__40951));
    Span4Mux_v I__9441 (
            .O(N__40959),
            .I(N__40951));
    LocalMux I__9440 (
            .O(N__40956),
            .I(buf_dds_3));
    Odrv4 I__9439 (
            .O(N__40951),
            .I(buf_dds_3));
    InMux I__9438 (
            .O(N__40946),
            .I(N__40941));
    InMux I__9437 (
            .O(N__40945),
            .I(N__40938));
    InMux I__9436 (
            .O(N__40944),
            .I(N__40935));
    LocalMux I__9435 (
            .O(N__40941),
            .I(N__40930));
    LocalMux I__9434 (
            .O(N__40938),
            .I(N__40930));
    LocalMux I__9433 (
            .O(N__40935),
            .I(n8));
    Odrv4 I__9432 (
            .O(N__40930),
            .I(n8));
    InMux I__9431 (
            .O(N__40925),
            .I(N__40922));
    LocalMux I__9430 (
            .O(N__40922),
            .I(N__40919));
    Span4Mux_h I__9429 (
            .O(N__40919),
            .I(N__40916));
    Span4Mux_v I__9428 (
            .O(N__40916),
            .I(N__40913));
    Odrv4 I__9427 (
            .O(N__40913),
            .I(n15188));
    InMux I__9426 (
            .O(N__40910),
            .I(N__40907));
    LocalMux I__9425 (
            .O(N__40907),
            .I(N__40903));
    InMux I__9424 (
            .O(N__40906),
            .I(N__40900));
    Span4Mux_h I__9423 (
            .O(N__40903),
            .I(N__40897));
    LocalMux I__9422 (
            .O(N__40900),
            .I(N__40894));
    Odrv4 I__9421 (
            .O(N__40897),
            .I(n12702));
    Odrv4 I__9420 (
            .O(N__40894),
            .I(n12702));
    CascadeMux I__9419 (
            .O(N__40889),
            .I(n15188_cascade_));
    InMux I__9418 (
            .O(N__40886),
            .I(N__40881));
    InMux I__9417 (
            .O(N__40885),
            .I(N__40876));
    InMux I__9416 (
            .O(N__40884),
            .I(N__40872));
    LocalMux I__9415 (
            .O(N__40881),
            .I(N__40869));
    InMux I__9414 (
            .O(N__40880),
            .I(N__40864));
    InMux I__9413 (
            .O(N__40879),
            .I(N__40864));
    LocalMux I__9412 (
            .O(N__40876),
            .I(N__40856));
    InMux I__9411 (
            .O(N__40875),
            .I(N__40853));
    LocalMux I__9410 (
            .O(N__40872),
            .I(N__40850));
    Span4Mux_h I__9409 (
            .O(N__40869),
            .I(N__40847));
    LocalMux I__9408 (
            .O(N__40864),
            .I(N__40844));
    InMux I__9407 (
            .O(N__40863),
            .I(N__40837));
    InMux I__9406 (
            .O(N__40862),
            .I(N__40837));
    InMux I__9405 (
            .O(N__40861),
            .I(N__40837));
    InMux I__9404 (
            .O(N__40860),
            .I(N__40834));
    InMux I__9403 (
            .O(N__40859),
            .I(N__40831));
    Span4Mux_v I__9402 (
            .O(N__40856),
            .I(N__40827));
    LocalMux I__9401 (
            .O(N__40853),
            .I(N__40822));
    Span12Mux_h I__9400 (
            .O(N__40850),
            .I(N__40822));
    Span4Mux_h I__9399 (
            .O(N__40847),
            .I(N__40813));
    Span4Mux_h I__9398 (
            .O(N__40844),
            .I(N__40813));
    LocalMux I__9397 (
            .O(N__40837),
            .I(N__40813));
    LocalMux I__9396 (
            .O(N__40834),
            .I(N__40813));
    LocalMux I__9395 (
            .O(N__40831),
            .I(N__40810));
    InMux I__9394 (
            .O(N__40830),
            .I(N__40807));
    Odrv4 I__9393 (
            .O(N__40827),
            .I(n8085));
    Odrv12 I__9392 (
            .O(N__40822),
            .I(n8085));
    Odrv4 I__9391 (
            .O(N__40813),
            .I(n8085));
    Odrv4 I__9390 (
            .O(N__40810),
            .I(n8085));
    LocalMux I__9389 (
            .O(N__40807),
            .I(n8085));
    CascadeMux I__9388 (
            .O(N__40796),
            .I(n6_adj_1171_cascade_));
    InMux I__9387 (
            .O(N__40793),
            .I(N__40790));
    LocalMux I__9386 (
            .O(N__40790),
            .I(N__40787));
    Odrv12 I__9385 (
            .O(N__40787),
            .I(n15190));
    InMux I__9384 (
            .O(N__40784),
            .I(N__40779));
    InMux I__9383 (
            .O(N__40783),
            .I(N__40776));
    CascadeMux I__9382 (
            .O(N__40782),
            .I(N__40773));
    LocalMux I__9381 (
            .O(N__40779),
            .I(N__40770));
    LocalMux I__9380 (
            .O(N__40776),
            .I(N__40767));
    InMux I__9379 (
            .O(N__40773),
            .I(N__40764));
    Span4Mux_h I__9378 (
            .O(N__40770),
            .I(N__40759));
    Span4Mux_h I__9377 (
            .O(N__40767),
            .I(N__40759));
    LocalMux I__9376 (
            .O(N__40764),
            .I(buf_adcdata3_12));
    Odrv4 I__9375 (
            .O(N__40759),
            .I(buf_adcdata3_12));
    InMux I__9374 (
            .O(N__40754),
            .I(N__40750));
    InMux I__9373 (
            .O(N__40753),
            .I(N__40747));
    LocalMux I__9372 (
            .O(N__40750),
            .I(N__40744));
    LocalMux I__9371 (
            .O(N__40747),
            .I(n24));
    Odrv4 I__9370 (
            .O(N__40744),
            .I(n24));
    InMux I__9369 (
            .O(N__40739),
            .I(N__40736));
    LocalMux I__9368 (
            .O(N__40736),
            .I(N__40733));
    Span4Mux_v I__9367 (
            .O(N__40733),
            .I(N__40727));
    InMux I__9366 (
            .O(N__40732),
            .I(N__40724));
    InMux I__9365 (
            .O(N__40731),
            .I(N__40719));
    InMux I__9364 (
            .O(N__40730),
            .I(N__40716));
    Span4Mux_h I__9363 (
            .O(N__40727),
            .I(N__40710));
    LocalMux I__9362 (
            .O(N__40724),
            .I(N__40710));
    InMux I__9361 (
            .O(N__40723),
            .I(N__40707));
    CascadeMux I__9360 (
            .O(N__40722),
            .I(N__40703));
    LocalMux I__9359 (
            .O(N__40719),
            .I(N__40700));
    LocalMux I__9358 (
            .O(N__40716),
            .I(N__40697));
    InMux I__9357 (
            .O(N__40715),
            .I(N__40694));
    Span4Mux_v I__9356 (
            .O(N__40710),
            .I(N__40687));
    LocalMux I__9355 (
            .O(N__40707),
            .I(N__40684));
    InMux I__9354 (
            .O(N__40706),
            .I(N__40681));
    InMux I__9353 (
            .O(N__40703),
            .I(N__40678));
    Span4Mux_v I__9352 (
            .O(N__40700),
            .I(N__40673));
    Span4Mux_h I__9351 (
            .O(N__40697),
            .I(N__40673));
    LocalMux I__9350 (
            .O(N__40694),
            .I(N__40670));
    InMux I__9349 (
            .O(N__40693),
            .I(N__40667));
    InMux I__9348 (
            .O(N__40692),
            .I(N__40664));
    InMux I__9347 (
            .O(N__40691),
            .I(N__40661));
    InMux I__9346 (
            .O(N__40690),
            .I(N__40658));
    Span4Mux_h I__9345 (
            .O(N__40687),
            .I(N__40652));
    Span4Mux_v I__9344 (
            .O(N__40684),
            .I(N__40652));
    LocalMux I__9343 (
            .O(N__40681),
            .I(N__40647));
    LocalMux I__9342 (
            .O(N__40678),
            .I(N__40647));
    Span4Mux_h I__9341 (
            .O(N__40673),
            .I(N__40644));
    Span4Mux_h I__9340 (
            .O(N__40670),
            .I(N__40641));
    LocalMux I__9339 (
            .O(N__40667),
            .I(N__40632));
    LocalMux I__9338 (
            .O(N__40664),
            .I(N__40632));
    LocalMux I__9337 (
            .O(N__40661),
            .I(N__40632));
    LocalMux I__9336 (
            .O(N__40658),
            .I(N__40632));
    InMux I__9335 (
            .O(N__40657),
            .I(N__40629));
    Span4Mux_h I__9334 (
            .O(N__40652),
            .I(N__40625));
    Span12Mux_h I__9333 (
            .O(N__40647),
            .I(N__40622));
    Span4Mux_h I__9332 (
            .O(N__40644),
            .I(N__40617));
    Span4Mux_v I__9331 (
            .O(N__40641),
            .I(N__40617));
    Span12Mux_h I__9330 (
            .O(N__40632),
            .I(N__40614));
    LocalMux I__9329 (
            .O(N__40629),
            .I(N__40611));
    InMux I__9328 (
            .O(N__40628),
            .I(N__40608));
    Odrv4 I__9327 (
            .O(N__40625),
            .I(comm_rx_buf_6));
    Odrv12 I__9326 (
            .O(N__40622),
            .I(comm_rx_buf_6));
    Odrv4 I__9325 (
            .O(N__40617),
            .I(comm_rx_buf_6));
    Odrv12 I__9324 (
            .O(N__40614),
            .I(comm_rx_buf_6));
    Odrv12 I__9323 (
            .O(N__40611),
            .I(comm_rx_buf_6));
    LocalMux I__9322 (
            .O(N__40608),
            .I(comm_rx_buf_6));
    InMux I__9321 (
            .O(N__40595),
            .I(N__40592));
    LocalMux I__9320 (
            .O(N__40592),
            .I(N__40589));
    Span4Mux_h I__9319 (
            .O(N__40589),
            .I(N__40586));
    Odrv4 I__9318 (
            .O(N__40586),
            .I(buf_data1_19));
    CascadeMux I__9317 (
            .O(N__40583),
            .I(N__40580));
    InMux I__9316 (
            .O(N__40580),
            .I(N__40576));
    InMux I__9315 (
            .O(N__40579),
            .I(N__40573));
    LocalMux I__9314 (
            .O(N__40576),
            .I(N__40570));
    LocalMux I__9313 (
            .O(N__40573),
            .I(data_idxvec_11));
    Odrv4 I__9312 (
            .O(N__40570),
            .I(data_idxvec_11));
    InMux I__9311 (
            .O(N__40565),
            .I(N__40562));
    LocalMux I__9310 (
            .O(N__40562),
            .I(N__40559));
    Span4Mux_h I__9309 (
            .O(N__40559),
            .I(N__40556));
    Span4Mux_h I__9308 (
            .O(N__40556),
            .I(N__40553));
    Odrv4 I__9307 (
            .O(N__40553),
            .I(n75));
    CascadeMux I__9306 (
            .O(N__40550),
            .I(n12_cascade_));
    InMux I__9305 (
            .O(N__40547),
            .I(N__40540));
    InMux I__9304 (
            .O(N__40546),
            .I(N__40535));
    InMux I__9303 (
            .O(N__40545),
            .I(N__40535));
    InMux I__9302 (
            .O(N__40544),
            .I(N__40529));
    InMux I__9301 (
            .O(N__40543),
            .I(N__40525));
    LocalMux I__9300 (
            .O(N__40540),
            .I(N__40520));
    LocalMux I__9299 (
            .O(N__40535),
            .I(N__40520));
    InMux I__9298 (
            .O(N__40534),
            .I(N__40517));
    InMux I__9297 (
            .O(N__40533),
            .I(N__40512));
    InMux I__9296 (
            .O(N__40532),
            .I(N__40512));
    LocalMux I__9295 (
            .O(N__40529),
            .I(N__40509));
    InMux I__9294 (
            .O(N__40528),
            .I(N__40506));
    LocalMux I__9293 (
            .O(N__40525),
            .I(N__40496));
    Span4Mux_v I__9292 (
            .O(N__40520),
            .I(N__40496));
    LocalMux I__9291 (
            .O(N__40517),
            .I(N__40496));
    LocalMux I__9290 (
            .O(N__40512),
            .I(N__40496));
    Span4Mux_v I__9289 (
            .O(N__40509),
            .I(N__40493));
    LocalMux I__9288 (
            .O(N__40506),
            .I(N__40490));
    InMux I__9287 (
            .O(N__40505),
            .I(N__40487));
    Span4Mux_v I__9286 (
            .O(N__40496),
            .I(N__40484));
    Sp12to4 I__9285 (
            .O(N__40493),
            .I(N__40477));
    Span12Mux_v I__9284 (
            .O(N__40490),
            .I(N__40477));
    LocalMux I__9283 (
            .O(N__40487),
            .I(N__40477));
    Odrv4 I__9282 (
            .O(N__40484),
            .I(n6301));
    Odrv12 I__9281 (
            .O(N__40477),
            .I(n6301));
    InMux I__9280 (
            .O(N__40472),
            .I(N__40465));
    InMux I__9279 (
            .O(N__40471),
            .I(N__40465));
    InMux I__9278 (
            .O(N__40470),
            .I(N__40451));
    LocalMux I__9277 (
            .O(N__40465),
            .I(N__40448));
    InMux I__9276 (
            .O(N__40464),
            .I(N__40445));
    InMux I__9275 (
            .O(N__40463),
            .I(N__40438));
    InMux I__9274 (
            .O(N__40462),
            .I(N__40438));
    InMux I__9273 (
            .O(N__40461),
            .I(N__40438));
    CascadeMux I__9272 (
            .O(N__40460),
            .I(N__40435));
    InMux I__9271 (
            .O(N__40459),
            .I(N__40428));
    InMux I__9270 (
            .O(N__40458),
            .I(N__40428));
    InMux I__9269 (
            .O(N__40457),
            .I(N__40425));
    InMux I__9268 (
            .O(N__40456),
            .I(N__40422));
    InMux I__9267 (
            .O(N__40455),
            .I(N__40419));
    InMux I__9266 (
            .O(N__40454),
            .I(N__40416));
    LocalMux I__9265 (
            .O(N__40451),
            .I(N__40413));
    Span4Mux_v I__9264 (
            .O(N__40448),
            .I(N__40408));
    LocalMux I__9263 (
            .O(N__40445),
            .I(N__40408));
    LocalMux I__9262 (
            .O(N__40438),
            .I(N__40405));
    InMux I__9261 (
            .O(N__40435),
            .I(N__40400));
    InMux I__9260 (
            .O(N__40434),
            .I(N__40400));
    InMux I__9259 (
            .O(N__40433),
            .I(N__40397));
    LocalMux I__9258 (
            .O(N__40428),
            .I(N__40394));
    LocalMux I__9257 (
            .O(N__40425),
            .I(N__40391));
    LocalMux I__9256 (
            .O(N__40422),
            .I(N__40388));
    LocalMux I__9255 (
            .O(N__40419),
            .I(N__40381));
    LocalMux I__9254 (
            .O(N__40416),
            .I(N__40381));
    Span4Mux_v I__9253 (
            .O(N__40413),
            .I(N__40381));
    Span4Mux_v I__9252 (
            .O(N__40408),
            .I(N__40378));
    Span4Mux_v I__9251 (
            .O(N__40405),
            .I(N__40375));
    LocalMux I__9250 (
            .O(N__40400),
            .I(N__40368));
    LocalMux I__9249 (
            .O(N__40397),
            .I(N__40368));
    Span4Mux_v I__9248 (
            .O(N__40394),
            .I(N__40368));
    Span12Mux_v I__9247 (
            .O(N__40391),
            .I(N__40365));
    Span4Mux_v I__9246 (
            .O(N__40388),
            .I(N__40358));
    Span4Mux_v I__9245 (
            .O(N__40381),
            .I(N__40358));
    Span4Mux_h I__9244 (
            .O(N__40378),
            .I(N__40358));
    Odrv4 I__9243 (
            .O(N__40375),
            .I(n8253));
    Odrv4 I__9242 (
            .O(N__40368),
            .I(n8253));
    Odrv12 I__9241 (
            .O(N__40365),
            .I(n8253));
    Odrv4 I__9240 (
            .O(N__40358),
            .I(n8253));
    InMux I__9239 (
            .O(N__40349),
            .I(N__40346));
    LocalMux I__9238 (
            .O(N__40346),
            .I(N__40342));
    InMux I__9237 (
            .O(N__40345),
            .I(N__40339));
    Span4Mux_v I__9236 (
            .O(N__40342),
            .I(N__40336));
    LocalMux I__9235 (
            .O(N__40339),
            .I(N__40333));
    Sp12to4 I__9234 (
            .O(N__40336),
            .I(N__40330));
    Odrv4 I__9233 (
            .O(N__40333),
            .I(n14_adj_1197));
    Odrv12 I__9232 (
            .O(N__40330),
            .I(n14_adj_1197));
    InMux I__9231 (
            .O(N__40325),
            .I(N__40320));
    InMux I__9230 (
            .O(N__40324),
            .I(N__40317));
    InMux I__9229 (
            .O(N__40323),
            .I(N__40314));
    LocalMux I__9228 (
            .O(N__40320),
            .I(N__40309));
    LocalMux I__9227 (
            .O(N__40317),
            .I(N__40309));
    LocalMux I__9226 (
            .O(N__40314),
            .I(req_data_cnt_2));
    Odrv12 I__9225 (
            .O(N__40309),
            .I(req_data_cnt_2));
    InMux I__9224 (
            .O(N__40304),
            .I(N__40299));
    InMux I__9223 (
            .O(N__40303),
            .I(N__40294));
    InMux I__9222 (
            .O(N__40302),
            .I(N__40294));
    LocalMux I__9221 (
            .O(N__40299),
            .I(comm_cmd_5));
    LocalMux I__9220 (
            .O(N__40294),
            .I(comm_cmd_5));
    InMux I__9219 (
            .O(N__40289),
            .I(N__40285));
    InMux I__9218 (
            .O(N__40288),
            .I(N__40281));
    LocalMux I__9217 (
            .O(N__40285),
            .I(N__40278));
    InMux I__9216 (
            .O(N__40284),
            .I(N__40275));
    LocalMux I__9215 (
            .O(N__40281),
            .I(comm_cmd_4));
    Odrv4 I__9214 (
            .O(N__40278),
            .I(comm_cmd_4));
    LocalMux I__9213 (
            .O(N__40275),
            .I(comm_cmd_4));
    InMux I__9212 (
            .O(N__40268),
            .I(N__40263));
    InMux I__9211 (
            .O(N__40267),
            .I(N__40258));
    InMux I__9210 (
            .O(N__40266),
            .I(N__40258));
    LocalMux I__9209 (
            .O(N__40263),
            .I(comm_cmd_6));
    LocalMux I__9208 (
            .O(N__40258),
            .I(comm_cmd_6));
    InMux I__9207 (
            .O(N__40253),
            .I(N__40248));
    InMux I__9206 (
            .O(N__40252),
            .I(N__40245));
    InMux I__9205 (
            .O(N__40251),
            .I(N__40242));
    LocalMux I__9204 (
            .O(N__40248),
            .I(N__40234));
    LocalMux I__9203 (
            .O(N__40245),
            .I(N__40229));
    LocalMux I__9202 (
            .O(N__40242),
            .I(N__40229));
    InMux I__9201 (
            .O(N__40241),
            .I(N__40226));
    InMux I__9200 (
            .O(N__40240),
            .I(N__40221));
    InMux I__9199 (
            .O(N__40239),
            .I(N__40218));
    InMux I__9198 (
            .O(N__40238),
            .I(N__40213));
    InMux I__9197 (
            .O(N__40237),
            .I(N__40213));
    Span4Mux_v I__9196 (
            .O(N__40234),
            .I(N__40203));
    Span4Mux_h I__9195 (
            .O(N__40229),
            .I(N__40203));
    LocalMux I__9194 (
            .O(N__40226),
            .I(N__40203));
    CascadeMux I__9193 (
            .O(N__40225),
            .I(N__40200));
    CascadeMux I__9192 (
            .O(N__40224),
            .I(N__40197));
    LocalMux I__9191 (
            .O(N__40221),
            .I(N__40190));
    LocalMux I__9190 (
            .O(N__40218),
            .I(N__40190));
    LocalMux I__9189 (
            .O(N__40213),
            .I(N__40187));
    InMux I__9188 (
            .O(N__40212),
            .I(N__40184));
    InMux I__9187 (
            .O(N__40211),
            .I(N__40181));
    InMux I__9186 (
            .O(N__40210),
            .I(N__40178));
    Span4Mux_h I__9185 (
            .O(N__40203),
            .I(N__40175));
    InMux I__9184 (
            .O(N__40200),
            .I(N__40172));
    InMux I__9183 (
            .O(N__40197),
            .I(N__40165));
    InMux I__9182 (
            .O(N__40196),
            .I(N__40165));
    InMux I__9181 (
            .O(N__40195),
            .I(N__40165));
    Span4Mux_v I__9180 (
            .O(N__40190),
            .I(N__40161));
    Span4Mux_v I__9179 (
            .O(N__40187),
            .I(N__40156));
    LocalMux I__9178 (
            .O(N__40184),
            .I(N__40156));
    LocalMux I__9177 (
            .O(N__40181),
            .I(N__40151));
    LocalMux I__9176 (
            .O(N__40178),
            .I(N__40151));
    Span4Mux_h I__9175 (
            .O(N__40175),
            .I(N__40148));
    LocalMux I__9174 (
            .O(N__40172),
            .I(N__40143));
    LocalMux I__9173 (
            .O(N__40165),
            .I(N__40143));
    InMux I__9172 (
            .O(N__40164),
            .I(N__40140));
    Span4Mux_h I__9171 (
            .O(N__40161),
            .I(N__40135));
    Span4Mux_v I__9170 (
            .O(N__40156),
            .I(N__40135));
    Odrv12 I__9169 (
            .O(N__40151),
            .I(n8043));
    Odrv4 I__9168 (
            .O(N__40148),
            .I(n8043));
    Odrv4 I__9167 (
            .O(N__40143),
            .I(n8043));
    LocalMux I__9166 (
            .O(N__40140),
            .I(n8043));
    Odrv4 I__9165 (
            .O(N__40135),
            .I(n8043));
    InMux I__9164 (
            .O(N__40124),
            .I(N__40113));
    InMux I__9163 (
            .O(N__40123),
            .I(N__40110));
    InMux I__9162 (
            .O(N__40122),
            .I(N__40107));
    InMux I__9161 (
            .O(N__40121),
            .I(N__40104));
    InMux I__9160 (
            .O(N__40120),
            .I(N__40101));
    InMux I__9159 (
            .O(N__40119),
            .I(N__40098));
    InMux I__9158 (
            .O(N__40118),
            .I(N__40095));
    InMux I__9157 (
            .O(N__40117),
            .I(N__40092));
    InMux I__9156 (
            .O(N__40116),
            .I(N__40089));
    LocalMux I__9155 (
            .O(N__40113),
            .I(N__40082));
    LocalMux I__9154 (
            .O(N__40110),
            .I(N__40082));
    LocalMux I__9153 (
            .O(N__40107),
            .I(N__40082));
    LocalMux I__9152 (
            .O(N__40104),
            .I(N__40077));
    LocalMux I__9151 (
            .O(N__40101),
            .I(N__40077));
    LocalMux I__9150 (
            .O(N__40098),
            .I(N__40068));
    LocalMux I__9149 (
            .O(N__40095),
            .I(N__40068));
    LocalMux I__9148 (
            .O(N__40092),
            .I(N__40068));
    LocalMux I__9147 (
            .O(N__40089),
            .I(N__40065));
    Span4Mux_v I__9146 (
            .O(N__40082),
            .I(N__40060));
    Span4Mux_v I__9145 (
            .O(N__40077),
            .I(N__40060));
    InMux I__9144 (
            .O(N__40076),
            .I(N__40057));
    InMux I__9143 (
            .O(N__40075),
            .I(N__40054));
    Span4Mux_v I__9142 (
            .O(N__40068),
            .I(N__40050));
    Span4Mux_h I__9141 (
            .O(N__40065),
            .I(N__40047));
    Span4Mux_h I__9140 (
            .O(N__40060),
            .I(N__40040));
    LocalMux I__9139 (
            .O(N__40057),
            .I(N__40040));
    LocalMux I__9138 (
            .O(N__40054),
            .I(N__40040));
    InMux I__9137 (
            .O(N__40053),
            .I(N__40037));
    Span4Mux_h I__9136 (
            .O(N__40050),
            .I(N__40033));
    Span4Mux_v I__9135 (
            .O(N__40047),
            .I(N__40028));
    Span4Mux_h I__9134 (
            .O(N__40040),
            .I(N__40028));
    LocalMux I__9133 (
            .O(N__40037),
            .I(N__40025));
    InMux I__9132 (
            .O(N__40036),
            .I(N__40022));
    Span4Mux_h I__9131 (
            .O(N__40033),
            .I(N__40018));
    Span4Mux_h I__9130 (
            .O(N__40028),
            .I(N__40015));
    Span12Mux_h I__9129 (
            .O(N__40025),
            .I(N__40010));
    LocalMux I__9128 (
            .O(N__40022),
            .I(N__40010));
    InMux I__9127 (
            .O(N__40021),
            .I(N__40007));
    Odrv4 I__9126 (
            .O(N__40018),
            .I(comm_rx_buf_2));
    Odrv4 I__9125 (
            .O(N__40015),
            .I(comm_rx_buf_2));
    Odrv12 I__9124 (
            .O(N__40010),
            .I(comm_rx_buf_2));
    LocalMux I__9123 (
            .O(N__40007),
            .I(comm_rx_buf_2));
    InMux I__9122 (
            .O(N__39998),
            .I(N__39992));
    InMux I__9121 (
            .O(N__39997),
            .I(N__39989));
    InMux I__9120 (
            .O(N__39996),
            .I(N__39986));
    InMux I__9119 (
            .O(N__39995),
            .I(N__39983));
    LocalMux I__9118 (
            .O(N__39992),
            .I(N__39980));
    LocalMux I__9117 (
            .O(N__39989),
            .I(N__39977));
    LocalMux I__9116 (
            .O(N__39986),
            .I(N__39974));
    LocalMux I__9115 (
            .O(N__39983),
            .I(N__39971));
    Span4Mux_h I__9114 (
            .O(N__39980),
            .I(N__39965));
    Span4Mux_h I__9113 (
            .O(N__39977),
            .I(N__39965));
    Span4Mux_v I__9112 (
            .O(N__39974),
            .I(N__39960));
    Span4Mux_h I__9111 (
            .O(N__39971),
            .I(N__39960));
    InMux I__9110 (
            .O(N__39970),
            .I(N__39957));
    Sp12to4 I__9109 (
            .O(N__39965),
            .I(N__39952));
    Sp12to4 I__9108 (
            .O(N__39960),
            .I(N__39952));
    LocalMux I__9107 (
            .O(N__39957),
            .I(comm_buf_1_2));
    Odrv12 I__9106 (
            .O(N__39952),
            .I(comm_buf_1_2));
    InMux I__9105 (
            .O(N__39947),
            .I(N__39944));
    LocalMux I__9104 (
            .O(N__39944),
            .I(N__39941));
    Span4Mux_v I__9103 (
            .O(N__39941),
            .I(N__39936));
    InMux I__9102 (
            .O(N__39940),
            .I(N__39933));
    InMux I__9101 (
            .O(N__39939),
            .I(N__39929));
    Span4Mux_h I__9100 (
            .O(N__39936),
            .I(N__39923));
    LocalMux I__9099 (
            .O(N__39933),
            .I(N__39923));
    InMux I__9098 (
            .O(N__39932),
            .I(N__39919));
    LocalMux I__9097 (
            .O(N__39929),
            .I(N__39916));
    InMux I__9096 (
            .O(N__39928),
            .I(N__39911));
    Span4Mux_v I__9095 (
            .O(N__39923),
            .I(N__39908));
    InMux I__9094 (
            .O(N__39922),
            .I(N__39905));
    LocalMux I__9093 (
            .O(N__39919),
            .I(N__39900));
    Span4Mux_h I__9092 (
            .O(N__39916),
            .I(N__39897));
    InMux I__9091 (
            .O(N__39915),
            .I(N__39894));
    InMux I__9090 (
            .O(N__39914),
            .I(N__39891));
    LocalMux I__9089 (
            .O(N__39911),
            .I(N__39888));
    Span4Mux_v I__9088 (
            .O(N__39908),
            .I(N__39882));
    LocalMux I__9087 (
            .O(N__39905),
            .I(N__39882));
    InMux I__9086 (
            .O(N__39904),
            .I(N__39879));
    InMux I__9085 (
            .O(N__39903),
            .I(N__39875));
    Span4Mux_h I__9084 (
            .O(N__39900),
            .I(N__39872));
    Span4Mux_v I__9083 (
            .O(N__39897),
            .I(N__39863));
    LocalMux I__9082 (
            .O(N__39894),
            .I(N__39863));
    LocalMux I__9081 (
            .O(N__39891),
            .I(N__39863));
    Span4Mux_v I__9080 (
            .O(N__39888),
            .I(N__39863));
    InMux I__9079 (
            .O(N__39887),
            .I(N__39860));
    Span4Mux_h I__9078 (
            .O(N__39882),
            .I(N__39854));
    LocalMux I__9077 (
            .O(N__39879),
            .I(N__39854));
    InMux I__9076 (
            .O(N__39878),
            .I(N__39851));
    LocalMux I__9075 (
            .O(N__39875),
            .I(N__39848));
    Sp12to4 I__9074 (
            .O(N__39872),
            .I(N__39841));
    Sp12to4 I__9073 (
            .O(N__39863),
            .I(N__39841));
    LocalMux I__9072 (
            .O(N__39860),
            .I(N__39841));
    InMux I__9071 (
            .O(N__39859),
            .I(N__39838));
    Span4Mux_h I__9070 (
            .O(N__39854),
            .I(N__39833));
    LocalMux I__9069 (
            .O(N__39851),
            .I(N__39833));
    Span12Mux_h I__9068 (
            .O(N__39848),
            .I(N__39825));
    Span12Mux_v I__9067 (
            .O(N__39841),
            .I(N__39825));
    LocalMux I__9066 (
            .O(N__39838),
            .I(N__39825));
    Span4Mux_v I__9065 (
            .O(N__39833),
            .I(N__39822));
    InMux I__9064 (
            .O(N__39832),
            .I(N__39819));
    Odrv12 I__9063 (
            .O(N__39825),
            .I(comm_rx_buf_4));
    Odrv4 I__9062 (
            .O(N__39822),
            .I(comm_rx_buf_4));
    LocalMux I__9061 (
            .O(N__39819),
            .I(comm_rx_buf_4));
    CascadeMux I__9060 (
            .O(N__39812),
            .I(n10363_cascade_));
    InMux I__9059 (
            .O(N__39809),
            .I(N__39805));
    InMux I__9058 (
            .O(N__39808),
            .I(N__39799));
    LocalMux I__9057 (
            .O(N__39805),
            .I(N__39792));
    InMux I__9056 (
            .O(N__39804),
            .I(N__39789));
    InMux I__9055 (
            .O(N__39803),
            .I(N__39786));
    CascadeMux I__9054 (
            .O(N__39802),
            .I(N__39782));
    LocalMux I__9053 (
            .O(N__39799),
            .I(N__39779));
    InMux I__9052 (
            .O(N__39798),
            .I(N__39776));
    InMux I__9051 (
            .O(N__39797),
            .I(N__39773));
    InMux I__9050 (
            .O(N__39796),
            .I(N__39770));
    CascadeMux I__9049 (
            .O(N__39795),
            .I(N__39767));
    Span4Mux_v I__9048 (
            .O(N__39792),
            .I(N__39760));
    LocalMux I__9047 (
            .O(N__39789),
            .I(N__39760));
    LocalMux I__9046 (
            .O(N__39786),
            .I(N__39757));
    InMux I__9045 (
            .O(N__39785),
            .I(N__39754));
    InMux I__9044 (
            .O(N__39782),
            .I(N__39751));
    Span4Mux_v I__9043 (
            .O(N__39779),
            .I(N__39746));
    LocalMux I__9042 (
            .O(N__39776),
            .I(N__39746));
    LocalMux I__9041 (
            .O(N__39773),
            .I(N__39741));
    LocalMux I__9040 (
            .O(N__39770),
            .I(N__39741));
    InMux I__9039 (
            .O(N__39767),
            .I(N__39738));
    InMux I__9038 (
            .O(N__39766),
            .I(N__39735));
    InMux I__9037 (
            .O(N__39765),
            .I(N__39732));
    Span4Mux_h I__9036 (
            .O(N__39760),
            .I(N__39728));
    Span4Mux_v I__9035 (
            .O(N__39757),
            .I(N__39723));
    LocalMux I__9034 (
            .O(N__39754),
            .I(N__39723));
    LocalMux I__9033 (
            .O(N__39751),
            .I(N__39720));
    Span4Mux_v I__9032 (
            .O(N__39746),
            .I(N__39711));
    Span4Mux_h I__9031 (
            .O(N__39741),
            .I(N__39711));
    LocalMux I__9030 (
            .O(N__39738),
            .I(N__39711));
    LocalMux I__9029 (
            .O(N__39735),
            .I(N__39711));
    LocalMux I__9028 (
            .O(N__39732),
            .I(N__39708));
    CascadeMux I__9027 (
            .O(N__39731),
            .I(N__39705));
    Span4Mux_h I__9026 (
            .O(N__39728),
            .I(N__39700));
    Span4Mux_h I__9025 (
            .O(N__39723),
            .I(N__39700));
    Span4Mux_v I__9024 (
            .O(N__39720),
            .I(N__39695));
    Span4Mux_h I__9023 (
            .O(N__39711),
            .I(N__39695));
    Span4Mux_v I__9022 (
            .O(N__39708),
            .I(N__39692));
    InMux I__9021 (
            .O(N__39705),
            .I(N__39689));
    Span4Mux_h I__9020 (
            .O(N__39700),
            .I(N__39685));
    Span4Mux_h I__9019 (
            .O(N__39695),
            .I(N__39682));
    Sp12to4 I__9018 (
            .O(N__39692),
            .I(N__39677));
    LocalMux I__9017 (
            .O(N__39689),
            .I(N__39677));
    InMux I__9016 (
            .O(N__39688),
            .I(N__39674));
    Odrv4 I__9015 (
            .O(N__39685),
            .I(comm_rx_buf_5));
    Odrv4 I__9014 (
            .O(N__39682),
            .I(comm_rx_buf_5));
    Odrv12 I__9013 (
            .O(N__39677),
            .I(comm_rx_buf_5));
    LocalMux I__9012 (
            .O(N__39674),
            .I(comm_rx_buf_5));
    InMux I__9011 (
            .O(N__39665),
            .I(N__39659));
    CascadeMux I__9010 (
            .O(N__39664),
            .I(N__39656));
    CascadeMux I__9009 (
            .O(N__39663),
            .I(N__39651));
    InMux I__9008 (
            .O(N__39662),
            .I(N__39647));
    LocalMux I__9007 (
            .O(N__39659),
            .I(N__39644));
    InMux I__9006 (
            .O(N__39656),
            .I(N__39641));
    InMux I__9005 (
            .O(N__39655),
            .I(N__39635));
    InMux I__9004 (
            .O(N__39654),
            .I(N__39635));
    InMux I__9003 (
            .O(N__39651),
            .I(N__39632));
    InMux I__9002 (
            .O(N__39650),
            .I(N__39629));
    LocalMux I__9001 (
            .O(N__39647),
            .I(N__39622));
    Span4Mux_v I__9000 (
            .O(N__39644),
            .I(N__39622));
    LocalMux I__8999 (
            .O(N__39641),
            .I(N__39622));
    InMux I__8998 (
            .O(N__39640),
            .I(N__39619));
    LocalMux I__8997 (
            .O(N__39635),
            .I(N__39614));
    LocalMux I__8996 (
            .O(N__39632),
            .I(N__39614));
    LocalMux I__8995 (
            .O(N__39629),
            .I(N__39609));
    Span4Mux_h I__8994 (
            .O(N__39622),
            .I(N__39609));
    LocalMux I__8993 (
            .O(N__39619),
            .I(N__39606));
    Span4Mux_h I__8992 (
            .O(N__39614),
            .I(N__39603));
    Span4Mux_h I__8991 (
            .O(N__39609),
            .I(N__39600));
    Odrv4 I__8990 (
            .O(N__39606),
            .I(n8062));
    Odrv4 I__8989 (
            .O(N__39603),
            .I(n8062));
    Odrv4 I__8988 (
            .O(N__39600),
            .I(n8062));
    CascadeMux I__8987 (
            .O(N__39593),
            .I(n8085_cascade_));
    InMux I__8986 (
            .O(N__39590),
            .I(N__39587));
    LocalMux I__8985 (
            .O(N__39587),
            .I(N__39584));
    Odrv4 I__8984 (
            .O(N__39584),
            .I(n14_adj_1152));
    CascadeMux I__8983 (
            .O(N__39581),
            .I(N__39577));
    CascadeMux I__8982 (
            .O(N__39580),
            .I(N__39574));
    InMux I__8981 (
            .O(N__39577),
            .I(N__39571));
    InMux I__8980 (
            .O(N__39574),
            .I(N__39565));
    LocalMux I__8979 (
            .O(N__39571),
            .I(N__39562));
    InMux I__8978 (
            .O(N__39570),
            .I(N__39557));
    InMux I__8977 (
            .O(N__39569),
            .I(N__39557));
    InMux I__8976 (
            .O(N__39568),
            .I(N__39553));
    LocalMux I__8975 (
            .O(N__39565),
            .I(N__39549));
    Span4Mux_v I__8974 (
            .O(N__39562),
            .I(N__39544));
    LocalMux I__8973 (
            .O(N__39557),
            .I(N__39544));
    CascadeMux I__8972 (
            .O(N__39556),
            .I(N__39538));
    LocalMux I__8971 (
            .O(N__39553),
            .I(N__39535));
    InMux I__8970 (
            .O(N__39552),
            .I(N__39532));
    Span4Mux_h I__8969 (
            .O(N__39549),
            .I(N__39527));
    Span4Mux_h I__8968 (
            .O(N__39544),
            .I(N__39527));
    InMux I__8967 (
            .O(N__39543),
            .I(N__39524));
    InMux I__8966 (
            .O(N__39542),
            .I(N__39521));
    InMux I__8965 (
            .O(N__39541),
            .I(N__39518));
    InMux I__8964 (
            .O(N__39538),
            .I(N__39515));
    Span4Mux_h I__8963 (
            .O(N__39535),
            .I(N__39512));
    LocalMux I__8962 (
            .O(N__39532),
            .I(N__39509));
    Span4Mux_h I__8961 (
            .O(N__39527),
            .I(N__39506));
    LocalMux I__8960 (
            .O(N__39524),
            .I(N__39497));
    LocalMux I__8959 (
            .O(N__39521),
            .I(N__39497));
    LocalMux I__8958 (
            .O(N__39518),
            .I(N__39497));
    LocalMux I__8957 (
            .O(N__39515),
            .I(N__39497));
    Span4Mux_h I__8956 (
            .O(N__39512),
            .I(N__39494));
    Span4Mux_h I__8955 (
            .O(N__39509),
            .I(N__39491));
    Span4Mux_h I__8954 (
            .O(N__39506),
            .I(N__39488));
    Span12Mux_h I__8953 (
            .O(N__39497),
            .I(N__39485));
    Odrv4 I__8952 (
            .O(N__39494),
            .I(n93));
    Odrv4 I__8951 (
            .O(N__39491),
            .I(n93));
    Odrv4 I__8950 (
            .O(N__39488),
            .I(n93));
    Odrv12 I__8949 (
            .O(N__39485),
            .I(n93));
    CascadeMux I__8948 (
            .O(N__39476),
            .I(N__39472));
    CascadeMux I__8947 (
            .O(N__39475),
            .I(N__39469));
    InMux I__8946 (
            .O(N__39472),
            .I(N__39466));
    InMux I__8945 (
            .O(N__39469),
            .I(N__39463));
    LocalMux I__8944 (
            .O(N__39466),
            .I(N__39458));
    LocalMux I__8943 (
            .O(N__39463),
            .I(N__39458));
    Span4Mux_h I__8942 (
            .O(N__39458),
            .I(N__39455));
    Odrv4 I__8941 (
            .O(N__39455),
            .I(n27));
    InMux I__8940 (
            .O(N__39452),
            .I(N__39449));
    LocalMux I__8939 (
            .O(N__39449),
            .I(n4));
    CascadeMux I__8938 (
            .O(N__39446),
            .I(n15309_cascade_));
    CascadeMux I__8937 (
            .O(N__39443),
            .I(N__39440));
    InMux I__8936 (
            .O(N__39440),
            .I(N__39437));
    LocalMux I__8935 (
            .O(N__39437),
            .I(N__39433));
    InMux I__8934 (
            .O(N__39436),
            .I(N__39430));
    Odrv4 I__8933 (
            .O(N__39433),
            .I(comm_state_3_N_402_3));
    LocalMux I__8932 (
            .O(N__39430),
            .I(comm_state_3_N_402_3));
    InMux I__8931 (
            .O(N__39425),
            .I(N__39422));
    LocalMux I__8930 (
            .O(N__39422),
            .I(N__39419));
    Odrv4 I__8929 (
            .O(N__39419),
            .I(n15637));
    InMux I__8928 (
            .O(N__39416),
            .I(N__39413));
    LocalMux I__8927 (
            .O(N__39413),
            .I(n13_adj_1040));
    InMux I__8926 (
            .O(N__39410),
            .I(N__39407));
    LocalMux I__8925 (
            .O(N__39407),
            .I(N__39404));
    Odrv4 I__8924 (
            .O(N__39404),
            .I(n22_adj_1078));
    CascadeMux I__8923 (
            .O(N__39401),
            .I(N__39398));
    InMux I__8922 (
            .O(N__39398),
            .I(N__39391));
    InMux I__8921 (
            .O(N__39397),
            .I(N__39387));
    InMux I__8920 (
            .O(N__39396),
            .I(N__39384));
    InMux I__8919 (
            .O(N__39395),
            .I(N__39380));
    InMux I__8918 (
            .O(N__39394),
            .I(N__39377));
    LocalMux I__8917 (
            .O(N__39391),
            .I(N__39374));
    InMux I__8916 (
            .O(N__39390),
            .I(N__39371));
    LocalMux I__8915 (
            .O(N__39387),
            .I(N__39368));
    LocalMux I__8914 (
            .O(N__39384),
            .I(N__39365));
    InMux I__8913 (
            .O(N__39383),
            .I(N__39362));
    LocalMux I__8912 (
            .O(N__39380),
            .I(N__39355));
    LocalMux I__8911 (
            .O(N__39377),
            .I(N__39355));
    Span4Mux_v I__8910 (
            .O(N__39374),
            .I(N__39350));
    LocalMux I__8909 (
            .O(N__39371),
            .I(N__39350));
    Span4Mux_v I__8908 (
            .O(N__39368),
            .I(N__39347));
    Span4Mux_v I__8907 (
            .O(N__39365),
            .I(N__39342));
    LocalMux I__8906 (
            .O(N__39362),
            .I(N__39342));
    InMux I__8905 (
            .O(N__39361),
            .I(N__39339));
    InMux I__8904 (
            .O(N__39360),
            .I(N__39335));
    Span4Mux_v I__8903 (
            .O(N__39355),
            .I(N__39328));
    Span4Mux_v I__8902 (
            .O(N__39350),
            .I(N__39328));
    Span4Mux_h I__8901 (
            .O(N__39347),
            .I(N__39323));
    Span4Mux_v I__8900 (
            .O(N__39342),
            .I(N__39323));
    LocalMux I__8899 (
            .O(N__39339),
            .I(N__39320));
    InMux I__8898 (
            .O(N__39338),
            .I(N__39317));
    LocalMux I__8897 (
            .O(N__39335),
            .I(N__39314));
    InMux I__8896 (
            .O(N__39334),
            .I(N__39311));
    InMux I__8895 (
            .O(N__39333),
            .I(N__39308));
    Span4Mux_h I__8894 (
            .O(N__39328),
            .I(N__39304));
    Span4Mux_h I__8893 (
            .O(N__39323),
            .I(N__39301));
    Span4Mux_v I__8892 (
            .O(N__39320),
            .I(N__39298));
    LocalMux I__8891 (
            .O(N__39317),
            .I(N__39289));
    Sp12to4 I__8890 (
            .O(N__39314),
            .I(N__39289));
    LocalMux I__8889 (
            .O(N__39311),
            .I(N__39289));
    LocalMux I__8888 (
            .O(N__39308),
            .I(N__39289));
    InMux I__8887 (
            .O(N__39307),
            .I(N__39286));
    Span4Mux_h I__8886 (
            .O(N__39304),
            .I(N__39283));
    Span4Mux_h I__8885 (
            .O(N__39301),
            .I(N__39278));
    Span4Mux_v I__8884 (
            .O(N__39298),
            .I(N__39278));
    Span12Mux_h I__8883 (
            .O(N__39289),
            .I(N__39275));
    LocalMux I__8882 (
            .O(N__39286),
            .I(N__39272));
    Odrv4 I__8881 (
            .O(N__39283),
            .I(comm_rx_buf_7));
    Odrv4 I__8880 (
            .O(N__39278),
            .I(comm_rx_buf_7));
    Odrv12 I__8879 (
            .O(N__39275),
            .I(comm_rx_buf_7));
    Odrv12 I__8878 (
            .O(N__39272),
            .I(comm_rx_buf_7));
    InMux I__8877 (
            .O(N__39263),
            .I(N__39260));
    LocalMux I__8876 (
            .O(N__39260),
            .I(N__39257));
    Span4Mux_v I__8875 (
            .O(N__39257),
            .I(N__39251));
    InMux I__8874 (
            .O(N__39256),
            .I(N__39248));
    CascadeMux I__8873 (
            .O(N__39255),
            .I(N__39245));
    InMux I__8872 (
            .O(N__39254),
            .I(N__39242));
    Span4Mux_h I__8871 (
            .O(N__39251),
            .I(N__39239));
    LocalMux I__8870 (
            .O(N__39248),
            .I(N__39236));
    InMux I__8869 (
            .O(N__39245),
            .I(N__39233));
    LocalMux I__8868 (
            .O(N__39242),
            .I(N__39230));
    Span4Mux_h I__8867 (
            .O(N__39239),
            .I(N__39227));
    Span12Mux_v I__8866 (
            .O(N__39236),
            .I(N__39224));
    LocalMux I__8865 (
            .O(N__39233),
            .I(comm_cmd_7));
    Odrv4 I__8864 (
            .O(N__39230),
            .I(comm_cmd_7));
    Odrv4 I__8863 (
            .O(N__39227),
            .I(comm_cmd_7));
    Odrv12 I__8862 (
            .O(N__39224),
            .I(comm_cmd_7));
    InMux I__8861 (
            .O(N__39215),
            .I(N__39210));
    InMux I__8860 (
            .O(N__39214),
            .I(N__39206));
    InMux I__8859 (
            .O(N__39213),
            .I(N__39202));
    LocalMux I__8858 (
            .O(N__39210),
            .I(N__39198));
    InMux I__8857 (
            .O(N__39209),
            .I(N__39195));
    LocalMux I__8856 (
            .O(N__39206),
            .I(N__39192));
    InMux I__8855 (
            .O(N__39205),
            .I(N__39189));
    LocalMux I__8854 (
            .O(N__39202),
            .I(N__39184));
    InMux I__8853 (
            .O(N__39201),
            .I(N__39181));
    Span4Mux_v I__8852 (
            .O(N__39198),
            .I(N__39170));
    LocalMux I__8851 (
            .O(N__39195),
            .I(N__39170));
    Span4Mux_v I__8850 (
            .O(N__39192),
            .I(N__39170));
    LocalMux I__8849 (
            .O(N__39189),
            .I(N__39167));
    InMux I__8848 (
            .O(N__39188),
            .I(N__39164));
    InMux I__8847 (
            .O(N__39187),
            .I(N__39161));
    Span4Mux_h I__8846 (
            .O(N__39184),
            .I(N__39158));
    LocalMux I__8845 (
            .O(N__39181),
            .I(N__39155));
    InMux I__8844 (
            .O(N__39180),
            .I(N__39152));
    InMux I__8843 (
            .O(N__39179),
            .I(N__39149));
    InMux I__8842 (
            .O(N__39178),
            .I(N__39146));
    InMux I__8841 (
            .O(N__39177),
            .I(N__39143));
    Span4Mux_h I__8840 (
            .O(N__39170),
            .I(N__39135));
    Span4Mux_v I__8839 (
            .O(N__39167),
            .I(N__39135));
    LocalMux I__8838 (
            .O(N__39164),
            .I(N__39135));
    LocalMux I__8837 (
            .O(N__39161),
            .I(N__39132));
    Span4Mux_h I__8836 (
            .O(N__39158),
            .I(N__39119));
    Span4Mux_v I__8835 (
            .O(N__39155),
            .I(N__39119));
    LocalMux I__8834 (
            .O(N__39152),
            .I(N__39119));
    LocalMux I__8833 (
            .O(N__39149),
            .I(N__39119));
    LocalMux I__8832 (
            .O(N__39146),
            .I(N__39119));
    LocalMux I__8831 (
            .O(N__39143),
            .I(N__39119));
    InMux I__8830 (
            .O(N__39142),
            .I(N__39115));
    Span4Mux_h I__8829 (
            .O(N__39135),
            .I(N__39112));
    Span4Mux_v I__8828 (
            .O(N__39132),
            .I(N__39109));
    Span4Mux_v I__8827 (
            .O(N__39119),
            .I(N__39106));
    InMux I__8826 (
            .O(N__39118),
            .I(N__39103));
    LocalMux I__8825 (
            .O(N__39115),
            .I(N__39100));
    Span4Mux_h I__8824 (
            .O(N__39112),
            .I(N__39097));
    Span4Mux_v I__8823 (
            .O(N__39109),
            .I(N__39092));
    Span4Mux_h I__8822 (
            .O(N__39106),
            .I(N__39092));
    LocalMux I__8821 (
            .O(N__39103),
            .I(comm_rx_buf_0));
    Odrv12 I__8820 (
            .O(N__39100),
            .I(comm_rx_buf_0));
    Odrv4 I__8819 (
            .O(N__39097),
            .I(comm_rx_buf_0));
    Odrv4 I__8818 (
            .O(N__39092),
            .I(comm_rx_buf_0));
    InMux I__8817 (
            .O(N__39083),
            .I(N__39077));
    InMux I__8816 (
            .O(N__39082),
            .I(N__39077));
    LocalMux I__8815 (
            .O(N__39077),
            .I(n8530));
    InMux I__8814 (
            .O(N__39074),
            .I(N__39068));
    InMux I__8813 (
            .O(N__39073),
            .I(N__39068));
    LocalMux I__8812 (
            .O(N__39068),
            .I(n15198));
    InMux I__8811 (
            .O(N__39065),
            .I(N__39062));
    LocalMux I__8810 (
            .O(N__39062),
            .I(n15266));
    CascadeMux I__8809 (
            .O(N__39059),
            .I(n15410_cascade_));
    CEMux I__8808 (
            .O(N__39056),
            .I(N__39053));
    LocalMux I__8807 (
            .O(N__39053),
            .I(n15130));
    CascadeMux I__8806 (
            .O(N__39050),
            .I(N__39047));
    InMux I__8805 (
            .O(N__39047),
            .I(N__39044));
    LocalMux I__8804 (
            .O(N__39044),
            .I(n15408));
    InMux I__8803 (
            .O(N__39041),
            .I(N__39037));
    InMux I__8802 (
            .O(N__39040),
            .I(N__39034));
    LocalMux I__8801 (
            .O(N__39037),
            .I(n10394));
    LocalMux I__8800 (
            .O(N__39034),
            .I(n10394));
    InMux I__8799 (
            .O(N__39029),
            .I(N__39026));
    LocalMux I__8798 (
            .O(N__39026),
            .I(n16190));
    InMux I__8797 (
            .O(N__39023),
            .I(N__39020));
    LocalMux I__8796 (
            .O(N__39020),
            .I(n15635));
    CascadeMux I__8795 (
            .O(N__39017),
            .I(N__39014));
    InMux I__8794 (
            .O(N__39014),
            .I(N__39010));
    CascadeMux I__8793 (
            .O(N__39013),
            .I(N__39007));
    LocalMux I__8792 (
            .O(N__39010),
            .I(N__39004));
    InMux I__8791 (
            .O(N__39007),
            .I(N__39001));
    Odrv4 I__8790 (
            .O(N__39004),
            .I(n12_adj_1027));
    LocalMux I__8789 (
            .O(N__39001),
            .I(n12_adj_1027));
    InMux I__8788 (
            .O(N__38996),
            .I(N__38992));
    InMux I__8787 (
            .O(N__38995),
            .I(N__38989));
    LocalMux I__8786 (
            .O(N__38992),
            .I(N__38984));
    LocalMux I__8785 (
            .O(N__38989),
            .I(N__38984));
    Span4Mux_v I__8784 (
            .O(N__38984),
            .I(N__38981));
    Odrv4 I__8783 (
            .O(N__38981),
            .I(n12622));
    InMux I__8782 (
            .O(N__38978),
            .I(N__38973));
    InMux I__8781 (
            .O(N__38977),
            .I(N__38968));
    InMux I__8780 (
            .O(N__38976),
            .I(N__38965));
    LocalMux I__8779 (
            .O(N__38973),
            .I(N__38962));
    InMux I__8778 (
            .O(N__38972),
            .I(N__38959));
    CascadeMux I__8777 (
            .O(N__38971),
            .I(N__38956));
    LocalMux I__8776 (
            .O(N__38968),
            .I(N__38953));
    LocalMux I__8775 (
            .O(N__38965),
            .I(N__38948));
    Span4Mux_h I__8774 (
            .O(N__38962),
            .I(N__38948));
    LocalMux I__8773 (
            .O(N__38959),
            .I(N__38945));
    InMux I__8772 (
            .O(N__38956),
            .I(N__38942));
    Span4Mux_h I__8771 (
            .O(N__38953),
            .I(N__38939));
    Sp12to4 I__8770 (
            .O(N__38948),
            .I(N__38936));
    Odrv4 I__8769 (
            .O(N__38945),
            .I(comm_buf_1_7));
    LocalMux I__8768 (
            .O(N__38942),
            .I(comm_buf_1_7));
    Odrv4 I__8767 (
            .O(N__38939),
            .I(comm_buf_1_7));
    Odrv12 I__8766 (
            .O(N__38936),
            .I(comm_buf_1_7));
    InMux I__8765 (
            .O(N__38927),
            .I(N__38920));
    InMux I__8764 (
            .O(N__38926),
            .I(N__38917));
    InMux I__8763 (
            .O(N__38925),
            .I(N__38914));
    InMux I__8762 (
            .O(N__38924),
            .I(N__38911));
    InMux I__8761 (
            .O(N__38923),
            .I(N__38908));
    LocalMux I__8760 (
            .O(N__38920),
            .I(N__38905));
    LocalMux I__8759 (
            .O(N__38917),
            .I(N__38899));
    LocalMux I__8758 (
            .O(N__38914),
            .I(N__38899));
    LocalMux I__8757 (
            .O(N__38911),
            .I(N__38896));
    LocalMux I__8756 (
            .O(N__38908),
            .I(N__38893));
    Span4Mux_h I__8755 (
            .O(N__38905),
            .I(N__38890));
    InMux I__8754 (
            .O(N__38904),
            .I(N__38887));
    Span4Mux_v I__8753 (
            .O(N__38899),
            .I(N__38884));
    Span4Mux_v I__8752 (
            .O(N__38896),
            .I(N__38881));
    Span4Mux_h I__8751 (
            .O(N__38893),
            .I(N__38878));
    Span4Mux_h I__8750 (
            .O(N__38890),
            .I(N__38875));
    LocalMux I__8749 (
            .O(N__38887),
            .I(N__38868));
    Span4Mux_h I__8748 (
            .O(N__38884),
            .I(N__38868));
    Span4Mux_h I__8747 (
            .O(N__38881),
            .I(N__38868));
    Span4Mux_h I__8746 (
            .O(N__38878),
            .I(N__38865));
    Span4Mux_v I__8745 (
            .O(N__38875),
            .I(N__38862));
    Sp12to4 I__8744 (
            .O(N__38868),
            .I(N__38859));
    Span4Mux_h I__8743 (
            .O(N__38865),
            .I(N__38854));
    Span4Mux_h I__8742 (
            .O(N__38862),
            .I(N__38854));
    Odrv12 I__8741 (
            .O(N__38859),
            .I(comm_buf_0_7));
    Odrv4 I__8740 (
            .O(N__38854),
            .I(comm_buf_0_7));
    InMux I__8739 (
            .O(N__38849),
            .I(N__38816));
    InMux I__8738 (
            .O(N__38848),
            .I(N__38816));
    InMux I__8737 (
            .O(N__38847),
            .I(N__38811));
    InMux I__8736 (
            .O(N__38846),
            .I(N__38811));
    InMux I__8735 (
            .O(N__38845),
            .I(N__38802));
    InMux I__8734 (
            .O(N__38844),
            .I(N__38802));
    InMux I__8733 (
            .O(N__38843),
            .I(N__38802));
    InMux I__8732 (
            .O(N__38842),
            .I(N__38795));
    InMux I__8731 (
            .O(N__38841),
            .I(N__38795));
    InMux I__8730 (
            .O(N__38840),
            .I(N__38795));
    InMux I__8729 (
            .O(N__38839),
            .I(N__38790));
    InMux I__8728 (
            .O(N__38838),
            .I(N__38790));
    InMux I__8727 (
            .O(N__38837),
            .I(N__38776));
    InMux I__8726 (
            .O(N__38836),
            .I(N__38767));
    InMux I__8725 (
            .O(N__38835),
            .I(N__38767));
    InMux I__8724 (
            .O(N__38834),
            .I(N__38767));
    InMux I__8723 (
            .O(N__38833),
            .I(N__38767));
    InMux I__8722 (
            .O(N__38832),
            .I(N__38760));
    InMux I__8721 (
            .O(N__38831),
            .I(N__38753));
    InMux I__8720 (
            .O(N__38830),
            .I(N__38753));
    InMux I__8719 (
            .O(N__38829),
            .I(N__38753));
    InMux I__8718 (
            .O(N__38828),
            .I(N__38746));
    InMux I__8717 (
            .O(N__38827),
            .I(N__38746));
    InMux I__8716 (
            .O(N__38826),
            .I(N__38746));
    InMux I__8715 (
            .O(N__38825),
            .I(N__38735));
    InMux I__8714 (
            .O(N__38824),
            .I(N__38735));
    InMux I__8713 (
            .O(N__38823),
            .I(N__38735));
    InMux I__8712 (
            .O(N__38822),
            .I(N__38735));
    InMux I__8711 (
            .O(N__38821),
            .I(N__38735));
    LocalMux I__8710 (
            .O(N__38816),
            .I(N__38730));
    LocalMux I__8709 (
            .O(N__38811),
            .I(N__38730));
    InMux I__8708 (
            .O(N__38810),
            .I(N__38725));
    InMux I__8707 (
            .O(N__38809),
            .I(N__38725));
    LocalMux I__8706 (
            .O(N__38802),
            .I(N__38718));
    LocalMux I__8705 (
            .O(N__38795),
            .I(N__38718));
    LocalMux I__8704 (
            .O(N__38790),
            .I(N__38718));
    InMux I__8703 (
            .O(N__38789),
            .I(N__38711));
    InMux I__8702 (
            .O(N__38788),
            .I(N__38711));
    InMux I__8701 (
            .O(N__38787),
            .I(N__38711));
    InMux I__8700 (
            .O(N__38786),
            .I(N__38704));
    InMux I__8699 (
            .O(N__38785),
            .I(N__38704));
    InMux I__8698 (
            .O(N__38784),
            .I(N__38704));
    InMux I__8697 (
            .O(N__38783),
            .I(N__38699));
    InMux I__8696 (
            .O(N__38782),
            .I(N__38699));
    InMux I__8695 (
            .O(N__38781),
            .I(N__38694));
    InMux I__8694 (
            .O(N__38780),
            .I(N__38694));
    InMux I__8693 (
            .O(N__38779),
            .I(N__38690));
    LocalMux I__8692 (
            .O(N__38776),
            .I(N__38686));
    LocalMux I__8691 (
            .O(N__38767),
            .I(N__38683));
    InMux I__8690 (
            .O(N__38766),
            .I(N__38680));
    InMux I__8689 (
            .O(N__38765),
            .I(N__38675));
    InMux I__8688 (
            .O(N__38764),
            .I(N__38675));
    InMux I__8687 (
            .O(N__38763),
            .I(N__38672));
    LocalMux I__8686 (
            .O(N__38760),
            .I(N__38669));
    LocalMux I__8685 (
            .O(N__38753),
            .I(N__38666));
    LocalMux I__8684 (
            .O(N__38746),
            .I(N__38655));
    LocalMux I__8683 (
            .O(N__38735),
            .I(N__38655));
    Span4Mux_v I__8682 (
            .O(N__38730),
            .I(N__38655));
    LocalMux I__8681 (
            .O(N__38725),
            .I(N__38655));
    Span4Mux_v I__8680 (
            .O(N__38718),
            .I(N__38655));
    LocalMux I__8679 (
            .O(N__38711),
            .I(N__38646));
    LocalMux I__8678 (
            .O(N__38704),
            .I(N__38646));
    LocalMux I__8677 (
            .O(N__38699),
            .I(N__38646));
    LocalMux I__8676 (
            .O(N__38694),
            .I(N__38646));
    CascadeMux I__8675 (
            .O(N__38693),
            .I(N__38643));
    LocalMux I__8674 (
            .O(N__38690),
            .I(N__38639));
    InMux I__8673 (
            .O(N__38689),
            .I(N__38636));
    Span4Mux_v I__8672 (
            .O(N__38686),
            .I(N__38631));
    Span4Mux_v I__8671 (
            .O(N__38683),
            .I(N__38631));
    LocalMux I__8670 (
            .O(N__38680),
            .I(N__38619));
    LocalMux I__8669 (
            .O(N__38675),
            .I(N__38619));
    LocalMux I__8668 (
            .O(N__38672),
            .I(N__38619));
    Span4Mux_v I__8667 (
            .O(N__38669),
            .I(N__38619));
    Span4Mux_v I__8666 (
            .O(N__38666),
            .I(N__38619));
    Span4Mux_h I__8665 (
            .O(N__38655),
            .I(N__38614));
    Span4Mux_v I__8664 (
            .O(N__38646),
            .I(N__38614));
    InMux I__8663 (
            .O(N__38643),
            .I(N__38609));
    InMux I__8662 (
            .O(N__38642),
            .I(N__38609));
    Span4Mux_v I__8661 (
            .O(N__38639),
            .I(N__38602));
    LocalMux I__8660 (
            .O(N__38636),
            .I(N__38602));
    Span4Mux_h I__8659 (
            .O(N__38631),
            .I(N__38602));
    InMux I__8658 (
            .O(N__38630),
            .I(N__38599));
    Span4Mux_h I__8657 (
            .O(N__38619),
            .I(N__38596));
    Span4Mux_h I__8656 (
            .O(N__38614),
            .I(N__38593));
    LocalMux I__8655 (
            .O(N__38609),
            .I(comm_index_0));
    Odrv4 I__8654 (
            .O(N__38602),
            .I(comm_index_0));
    LocalMux I__8653 (
            .O(N__38599),
            .I(comm_index_0));
    Odrv4 I__8652 (
            .O(N__38596),
            .I(comm_index_0));
    Odrv4 I__8651 (
            .O(N__38593),
            .I(comm_index_0));
    InMux I__8650 (
            .O(N__38582),
            .I(N__38579));
    LocalMux I__8649 (
            .O(N__38579),
            .I(N__38576));
    Span12Mux_h I__8648 (
            .O(N__38576),
            .I(N__38573));
    Odrv12 I__8647 (
            .O(N__38573),
            .I(n15381));
    CascadeMux I__8646 (
            .O(N__38570),
            .I(n12846_cascade_));
    InMux I__8645 (
            .O(N__38567),
            .I(N__38564));
    LocalMux I__8644 (
            .O(N__38564),
            .I(n4_adj_1179));
    CascadeMux I__8643 (
            .O(N__38561),
            .I(N__38555));
    CascadeMux I__8642 (
            .O(N__38560),
            .I(N__38552));
    CascadeMux I__8641 (
            .O(N__38559),
            .I(N__38549));
    InMux I__8640 (
            .O(N__38558),
            .I(N__38545));
    InMux I__8639 (
            .O(N__38555),
            .I(N__38538));
    InMux I__8638 (
            .O(N__38552),
            .I(N__38538));
    InMux I__8637 (
            .O(N__38549),
            .I(N__38538));
    CascadeMux I__8636 (
            .O(N__38548),
            .I(N__38535));
    LocalMux I__8635 (
            .O(N__38545),
            .I(N__38530));
    LocalMux I__8634 (
            .O(N__38538),
            .I(N__38527));
    InMux I__8633 (
            .O(N__38535),
            .I(N__38522));
    InMux I__8632 (
            .O(N__38534),
            .I(N__38522));
    InMux I__8631 (
            .O(N__38533),
            .I(N__38519));
    Span4Mux_h I__8630 (
            .O(N__38530),
            .I(N__38516));
    Span4Mux_v I__8629 (
            .O(N__38527),
            .I(N__38511));
    LocalMux I__8628 (
            .O(N__38522),
            .I(N__38511));
    LocalMux I__8627 (
            .O(N__38519),
            .I(N__38508));
    Odrv4 I__8626 (
            .O(N__38516),
            .I(n15204));
    Odrv4 I__8625 (
            .O(N__38511),
            .I(n15204));
    Odrv4 I__8624 (
            .O(N__38508),
            .I(n15204));
    CascadeMux I__8623 (
            .O(N__38501),
            .I(n4_adj_1184_cascade_));
    InMux I__8622 (
            .O(N__38498),
            .I(N__38495));
    LocalMux I__8621 (
            .O(N__38495),
            .I(N__38492));
    Odrv4 I__8620 (
            .O(N__38492),
            .I(n15290));
    CascadeMux I__8619 (
            .O(N__38489),
            .I(n15241_cascade_));
    InMux I__8618 (
            .O(N__38486),
            .I(N__38480));
    InMux I__8617 (
            .O(N__38485),
            .I(N__38480));
    LocalMux I__8616 (
            .O(N__38480),
            .I(n15108));
    CEMux I__8615 (
            .O(N__38477),
            .I(N__38474));
    LocalMux I__8614 (
            .O(N__38474),
            .I(N__38471));
    Span4Mux_v I__8613 (
            .O(N__38471),
            .I(N__38468));
    Odrv4 I__8612 (
            .O(N__38468),
            .I(n15128));
    InMux I__8611 (
            .O(N__38465),
            .I(N__38462));
    LocalMux I__8610 (
            .O(N__38462),
            .I(N__38459));
    Span4Mux_v I__8609 (
            .O(N__38459),
            .I(N__38456));
    Odrv4 I__8608 (
            .O(N__38456),
            .I(\comm_spi.n10438 ));
    SRMux I__8607 (
            .O(N__38453),
            .I(N__38450));
    LocalMux I__8606 (
            .O(N__38450),
            .I(N__38447));
    Span4Mux_h I__8605 (
            .O(N__38447),
            .I(N__38444));
    Span4Mux_h I__8604 (
            .O(N__38444),
            .I(N__38441));
    Odrv4 I__8603 (
            .O(N__38441),
            .I(\comm_spi.iclk_N_802 ));
    InMux I__8602 (
            .O(N__38438),
            .I(N__38435));
    LocalMux I__8601 (
            .O(N__38435),
            .I(\comm_spi.n16890 ));
    InMux I__8600 (
            .O(N__38432),
            .I(N__38429));
    LocalMux I__8599 (
            .O(N__38429),
            .I(\comm_spi.n10455 ));
    CascadeMux I__8598 (
            .O(N__38426),
            .I(\comm_spi.n16890_cascade_ ));
    InMux I__8597 (
            .O(N__38423),
            .I(N__38420));
    LocalMux I__8596 (
            .O(N__38420),
            .I(N__38409));
    InMux I__8595 (
            .O(N__38419),
            .I(N__38406));
    InMux I__8594 (
            .O(N__38418),
            .I(N__38391));
    InMux I__8593 (
            .O(N__38417),
            .I(N__38391));
    InMux I__8592 (
            .O(N__38416),
            .I(N__38391));
    InMux I__8591 (
            .O(N__38415),
            .I(N__38391));
    InMux I__8590 (
            .O(N__38414),
            .I(N__38391));
    InMux I__8589 (
            .O(N__38413),
            .I(N__38391));
    InMux I__8588 (
            .O(N__38412),
            .I(N__38391));
    Odrv12 I__8587 (
            .O(N__38409),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__8586 (
            .O(N__38406),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__8585 (
            .O(N__38391),
            .I(\comm_spi.bit_cnt_3 ));
    InMux I__8584 (
            .O(N__38384),
            .I(N__38381));
    LocalMux I__8583 (
            .O(N__38381),
            .I(N__38378));
    Span4Mux_v I__8582 (
            .O(N__38378),
            .I(N__38368));
    InMux I__8581 (
            .O(N__38377),
            .I(N__38353));
    InMux I__8580 (
            .O(N__38376),
            .I(N__38353));
    InMux I__8579 (
            .O(N__38375),
            .I(N__38353));
    InMux I__8578 (
            .O(N__38374),
            .I(N__38353));
    InMux I__8577 (
            .O(N__38373),
            .I(N__38353));
    InMux I__8576 (
            .O(N__38372),
            .I(N__38353));
    InMux I__8575 (
            .O(N__38371),
            .I(N__38353));
    Odrv4 I__8574 (
            .O(N__38368),
            .I(\comm_spi.n12175 ));
    LocalMux I__8573 (
            .O(N__38353),
            .I(\comm_spi.n12175 ));
    InMux I__8572 (
            .O(N__38348),
            .I(N__38344));
    InMux I__8571 (
            .O(N__38347),
            .I(N__38341));
    LocalMux I__8570 (
            .O(N__38344),
            .I(N__38338));
    LocalMux I__8569 (
            .O(N__38341),
            .I(data_idxvec_5));
    Odrv4 I__8568 (
            .O(N__38338),
            .I(data_idxvec_5));
    InMux I__8567 (
            .O(N__38333),
            .I(N__38328));
    InMux I__8566 (
            .O(N__38332),
            .I(N__38325));
    InMux I__8565 (
            .O(N__38331),
            .I(N__38322));
    LocalMux I__8564 (
            .O(N__38328),
            .I(data_cntvec_5));
    LocalMux I__8563 (
            .O(N__38325),
            .I(data_cntvec_5));
    LocalMux I__8562 (
            .O(N__38322),
            .I(data_cntvec_5));
    InMux I__8561 (
            .O(N__38315),
            .I(N__38312));
    LocalMux I__8560 (
            .O(N__38312),
            .I(N__38309));
    Span4Mux_h I__8559 (
            .O(N__38309),
            .I(N__38306));
    Odrv4 I__8558 (
            .O(N__38306),
            .I(buf_data1_13));
    CascadeMux I__8557 (
            .O(N__38303),
            .I(n4192_cascade_));
    InMux I__8556 (
            .O(N__38300),
            .I(N__38297));
    LocalMux I__8555 (
            .O(N__38297),
            .I(n4229));
    CascadeMux I__8554 (
            .O(N__38294),
            .I(N__38291));
    InMux I__8553 (
            .O(N__38291),
            .I(N__38288));
    LocalMux I__8552 (
            .O(N__38288),
            .I(N__38285));
    Sp12to4 I__8551 (
            .O(N__38285),
            .I(N__38280));
    InMux I__8550 (
            .O(N__38284),
            .I(N__38277));
    CascadeMux I__8549 (
            .O(N__38283),
            .I(N__38274));
    Span12Mux_s9_v I__8548 (
            .O(N__38280),
            .I(N__38269));
    LocalMux I__8547 (
            .O(N__38277),
            .I(N__38269));
    InMux I__8546 (
            .O(N__38274),
            .I(N__38266));
    Odrv12 I__8545 (
            .O(N__38269),
            .I(cmd_rdadctmp_18_adj_1058));
    LocalMux I__8544 (
            .O(N__38266),
            .I(cmd_rdadctmp_18_adj_1058));
    InMux I__8543 (
            .O(N__38261),
            .I(N__38258));
    LocalMux I__8542 (
            .O(N__38258),
            .I(N__38254));
    InMux I__8541 (
            .O(N__38257),
            .I(N__38251));
    Span4Mux_v I__8540 (
            .O(N__38254),
            .I(N__38248));
    LocalMux I__8539 (
            .O(N__38251),
            .I(buf_adcdata2_10));
    Odrv4 I__8538 (
            .O(N__38248),
            .I(buf_adcdata2_10));
    InMux I__8537 (
            .O(N__38243),
            .I(N__38239));
    InMux I__8536 (
            .O(N__38242),
            .I(N__38236));
    LocalMux I__8535 (
            .O(N__38239),
            .I(N__38233));
    LocalMux I__8534 (
            .O(N__38236),
            .I(data_idxvec_1));
    Odrv12 I__8533 (
            .O(N__38233),
            .I(data_idxvec_1));
    InMux I__8532 (
            .O(N__38228),
            .I(N__38224));
    InMux I__8531 (
            .O(N__38227),
            .I(N__38220));
    LocalMux I__8530 (
            .O(N__38224),
            .I(N__38217));
    InMux I__8529 (
            .O(N__38223),
            .I(N__38214));
    LocalMux I__8528 (
            .O(N__38220),
            .I(data_cntvec_1));
    Odrv4 I__8527 (
            .O(N__38217),
            .I(data_cntvec_1));
    LocalMux I__8526 (
            .O(N__38214),
            .I(data_cntvec_1));
    CascadeMux I__8525 (
            .O(N__38207),
            .I(N__38204));
    InMux I__8524 (
            .O(N__38204),
            .I(N__38201));
    LocalMux I__8523 (
            .O(N__38201),
            .I(N__38197));
    InMux I__8522 (
            .O(N__38200),
            .I(N__38194));
    Sp12to4 I__8521 (
            .O(N__38197),
            .I(N__38188));
    LocalMux I__8520 (
            .O(N__38194),
            .I(N__38188));
    CascadeMux I__8519 (
            .O(N__38193),
            .I(N__38185));
    Span12Mux_h I__8518 (
            .O(N__38188),
            .I(N__38182));
    InMux I__8517 (
            .O(N__38185),
            .I(N__38179));
    Odrv12 I__8516 (
            .O(N__38182),
            .I(cmd_rdadctmp_16_adj_1096));
    LocalMux I__8515 (
            .O(N__38179),
            .I(cmd_rdadctmp_16_adj_1096));
    InMux I__8514 (
            .O(N__38174),
            .I(N__38171));
    LocalMux I__8513 (
            .O(N__38171),
            .I(N__38167));
    InMux I__8512 (
            .O(N__38170),
            .I(N__38163));
    Span4Mux_v I__8511 (
            .O(N__38167),
            .I(N__38160));
    InMux I__8510 (
            .O(N__38166),
            .I(N__38157));
    LocalMux I__8509 (
            .O(N__38163),
            .I(req_data_cnt_3));
    Odrv4 I__8508 (
            .O(N__38160),
            .I(req_data_cnt_3));
    LocalMux I__8507 (
            .O(N__38157),
            .I(req_data_cnt_3));
    InMux I__8506 (
            .O(N__38150),
            .I(N__38147));
    LocalMux I__8505 (
            .O(N__38147),
            .I(N__38142));
    InMux I__8504 (
            .O(N__38146),
            .I(N__38137));
    InMux I__8503 (
            .O(N__38145),
            .I(N__38137));
    Odrv4 I__8502 (
            .O(N__38142),
            .I(acadc_skipCount_3));
    LocalMux I__8501 (
            .O(N__38137),
            .I(acadc_skipCount_3));
    InMux I__8500 (
            .O(N__38132),
            .I(N__38128));
    InMux I__8499 (
            .O(N__38131),
            .I(N__38124));
    LocalMux I__8498 (
            .O(N__38128),
            .I(N__38119));
    InMux I__8497 (
            .O(N__38127),
            .I(N__38116));
    LocalMux I__8496 (
            .O(N__38124),
            .I(N__38113));
    InMux I__8495 (
            .O(N__38123),
            .I(N__38108));
    InMux I__8494 (
            .O(N__38122),
            .I(N__38108));
    Span4Mux_v I__8493 (
            .O(N__38119),
            .I(N__38103));
    LocalMux I__8492 (
            .O(N__38116),
            .I(N__38103));
    Span4Mux_h I__8491 (
            .O(N__38113),
            .I(N__38098));
    LocalMux I__8490 (
            .O(N__38108),
            .I(N__38098));
    Span4Mux_v I__8489 (
            .O(N__38103),
            .I(N__38087));
    Span4Mux_v I__8488 (
            .O(N__38098),
            .I(N__38084));
    InMux I__8487 (
            .O(N__38097),
            .I(N__38081));
    InMux I__8486 (
            .O(N__38096),
            .I(N__38074));
    InMux I__8485 (
            .O(N__38095),
            .I(N__38074));
    InMux I__8484 (
            .O(N__38094),
            .I(N__38074));
    InMux I__8483 (
            .O(N__38093),
            .I(N__38071));
    InMux I__8482 (
            .O(N__38092),
            .I(N__38064));
    InMux I__8481 (
            .O(N__38091),
            .I(N__38064));
    InMux I__8480 (
            .O(N__38090),
            .I(N__38064));
    Span4Mux_h I__8479 (
            .O(N__38087),
            .I(N__38061));
    Odrv4 I__8478 (
            .O(N__38084),
            .I(eis_state_1));
    LocalMux I__8477 (
            .O(N__38081),
            .I(eis_state_1));
    LocalMux I__8476 (
            .O(N__38074),
            .I(eis_state_1));
    LocalMux I__8475 (
            .O(N__38071),
            .I(eis_state_1));
    LocalMux I__8474 (
            .O(N__38064),
            .I(eis_state_1));
    Odrv4 I__8473 (
            .O(N__38061),
            .I(eis_state_1));
    CEMux I__8472 (
            .O(N__38048),
            .I(N__38044));
    InMux I__8471 (
            .O(N__38047),
            .I(N__38038));
    LocalMux I__8470 (
            .O(N__38044),
            .I(N__38035));
    CEMux I__8469 (
            .O(N__38043),
            .I(N__38032));
    CEMux I__8468 (
            .O(N__38042),
            .I(N__38029));
    CEMux I__8467 (
            .O(N__38041),
            .I(N__38026));
    LocalMux I__8466 (
            .O(N__38038),
            .I(N__38023));
    Span4Mux_v I__8465 (
            .O(N__38035),
            .I(N__38016));
    LocalMux I__8464 (
            .O(N__38032),
            .I(N__38016));
    LocalMux I__8463 (
            .O(N__38029),
            .I(N__38016));
    LocalMux I__8462 (
            .O(N__38026),
            .I(N__38011));
    Span4Mux_v I__8461 (
            .O(N__38023),
            .I(N__38011));
    Odrv4 I__8460 (
            .O(N__38016),
            .I(n9790));
    Odrv4 I__8459 (
            .O(N__38011),
            .I(n9790));
    SRMux I__8458 (
            .O(N__38006),
            .I(N__38002));
    SRMux I__8457 (
            .O(N__38005),
            .I(N__37999));
    LocalMux I__8456 (
            .O(N__38002),
            .I(N__37996));
    LocalMux I__8455 (
            .O(N__37999),
            .I(N__37991));
    Span4Mux_v I__8454 (
            .O(N__37996),
            .I(N__37988));
    SRMux I__8453 (
            .O(N__37995),
            .I(N__37985));
    SRMux I__8452 (
            .O(N__37994),
            .I(N__37982));
    Span12Mux_v I__8451 (
            .O(N__37991),
            .I(N__37979));
    Span4Mux_h I__8450 (
            .O(N__37988),
            .I(N__37976));
    LocalMux I__8449 (
            .O(N__37985),
            .I(n10483));
    LocalMux I__8448 (
            .O(N__37982),
            .I(n10483));
    Odrv12 I__8447 (
            .O(N__37979),
            .I(n10483));
    Odrv4 I__8446 (
            .O(N__37976),
            .I(n10483));
    InMux I__8445 (
            .O(N__37967),
            .I(N__37964));
    LocalMux I__8444 (
            .O(N__37964),
            .I(N__37961));
    Span4Mux_v I__8443 (
            .O(N__37961),
            .I(N__37957));
    InMux I__8442 (
            .O(N__37960),
            .I(N__37954));
    Odrv4 I__8441 (
            .O(N__37957),
            .I(\comm_spi.n16887 ));
    LocalMux I__8440 (
            .O(N__37954),
            .I(\comm_spi.n16887 ));
    InMux I__8439 (
            .O(N__37949),
            .I(N__37946));
    LocalMux I__8438 (
            .O(N__37946),
            .I(N__37942));
    InMux I__8437 (
            .O(N__37945),
            .I(N__37939));
    Span4Mux_v I__8436 (
            .O(N__37942),
            .I(N__37934));
    LocalMux I__8435 (
            .O(N__37939),
            .I(N__37934));
    Span4Mux_v I__8434 (
            .O(N__37934),
            .I(N__37931));
    Span4Mux_h I__8433 (
            .O(N__37931),
            .I(N__37928));
    Span4Mux_h I__8432 (
            .O(N__37928),
            .I(N__37925));
    Odrv4 I__8431 (
            .O(N__37925),
            .I(n14_adj_1169));
    CascadeMux I__8430 (
            .O(N__37922),
            .I(N__37918));
    InMux I__8429 (
            .O(N__37921),
            .I(N__37912));
    InMux I__8428 (
            .O(N__37918),
            .I(N__37912));
    InMux I__8427 (
            .O(N__37917),
            .I(N__37909));
    LocalMux I__8426 (
            .O(N__37912),
            .I(N__37906));
    LocalMux I__8425 (
            .O(N__37909),
            .I(req_data_cnt_6));
    Odrv4 I__8424 (
            .O(N__37906),
            .I(req_data_cnt_6));
    InMux I__8423 (
            .O(N__37901),
            .I(N__37898));
    LocalMux I__8422 (
            .O(N__37898),
            .I(N__37895));
    Span4Mux_v I__8421 (
            .O(N__37895),
            .I(N__37892));
    Odrv4 I__8420 (
            .O(N__37892),
            .I(n4204));
    CascadeMux I__8419 (
            .O(N__37889),
            .I(n4249_cascade_));
    CascadeMux I__8418 (
            .O(N__37886),
            .I(n4259_cascade_));
    InMux I__8417 (
            .O(N__37883),
            .I(N__37879));
    InMux I__8416 (
            .O(N__37882),
            .I(N__37875));
    LocalMux I__8415 (
            .O(N__37879),
            .I(N__37871));
    InMux I__8414 (
            .O(N__37878),
            .I(N__37867));
    LocalMux I__8413 (
            .O(N__37875),
            .I(N__37864));
    InMux I__8412 (
            .O(N__37874),
            .I(N__37861));
    Span4Mux_h I__8411 (
            .O(N__37871),
            .I(N__37858));
    InMux I__8410 (
            .O(N__37870),
            .I(N__37855));
    LocalMux I__8409 (
            .O(N__37867),
            .I(N__37852));
    Span4Mux_v I__8408 (
            .O(N__37864),
            .I(N__37847));
    LocalMux I__8407 (
            .O(N__37861),
            .I(N__37847));
    Span4Mux_v I__8406 (
            .O(N__37858),
            .I(N__37844));
    LocalMux I__8405 (
            .O(N__37855),
            .I(N__37841));
    Span12Mux_h I__8404 (
            .O(N__37852),
            .I(N__37838));
    Odrv4 I__8403 (
            .O(N__37847),
            .I(comm_buf_1_5));
    Odrv4 I__8402 (
            .O(N__37844),
            .I(comm_buf_1_5));
    Odrv4 I__8401 (
            .O(N__37841),
            .I(comm_buf_1_5));
    Odrv12 I__8400 (
            .O(N__37838),
            .I(comm_buf_1_5));
    CascadeMux I__8399 (
            .O(N__37829),
            .I(N__37825));
    InMux I__8398 (
            .O(N__37828),
            .I(N__37822));
    InMux I__8397 (
            .O(N__37825),
            .I(N__37819));
    LocalMux I__8396 (
            .O(N__37822),
            .I(N__37816));
    LocalMux I__8395 (
            .O(N__37819),
            .I(data_idxvec_4));
    Odrv4 I__8394 (
            .O(N__37816),
            .I(data_idxvec_4));
    InMux I__8393 (
            .O(N__37811),
            .I(N__37807));
    InMux I__8392 (
            .O(N__37810),
            .I(N__37803));
    LocalMux I__8391 (
            .O(N__37807),
            .I(N__37800));
    InMux I__8390 (
            .O(N__37806),
            .I(N__37797));
    LocalMux I__8389 (
            .O(N__37803),
            .I(data_cntvec_4));
    Odrv4 I__8388 (
            .O(N__37800),
            .I(data_cntvec_4));
    LocalMux I__8387 (
            .O(N__37797),
            .I(data_cntvec_4));
    InMux I__8386 (
            .O(N__37790),
            .I(N__37787));
    LocalMux I__8385 (
            .O(N__37787),
            .I(N__37784));
    Span4Mux_v I__8384 (
            .O(N__37784),
            .I(N__37781));
    Span4Mux_h I__8383 (
            .O(N__37781),
            .I(N__37778));
    Odrv4 I__8382 (
            .O(N__37778),
            .I(buf_data1_12));
    CascadeMux I__8381 (
            .O(N__37775),
            .I(n4193_cascade_));
    CascadeMux I__8380 (
            .O(N__37772),
            .I(N__37768));
    CascadeMux I__8379 (
            .O(N__37771),
            .I(N__37764));
    InMux I__8378 (
            .O(N__37768),
            .I(N__37761));
    InMux I__8377 (
            .O(N__37767),
            .I(N__37758));
    InMux I__8376 (
            .O(N__37764),
            .I(N__37755));
    LocalMux I__8375 (
            .O(N__37761),
            .I(req_data_cnt_5));
    LocalMux I__8374 (
            .O(N__37758),
            .I(req_data_cnt_5));
    LocalMux I__8373 (
            .O(N__37755),
            .I(req_data_cnt_5));
    InMux I__8372 (
            .O(N__37748),
            .I(N__37745));
    LocalMux I__8371 (
            .O(N__37745),
            .I(N__37742));
    Span4Mux_h I__8370 (
            .O(N__37742),
            .I(N__37737));
    InMux I__8369 (
            .O(N__37741),
            .I(N__37732));
    InMux I__8368 (
            .O(N__37740),
            .I(N__37732));
    Odrv4 I__8367 (
            .O(N__37737),
            .I(acadc_skipCount_5));
    LocalMux I__8366 (
            .O(N__37732),
            .I(acadc_skipCount_5));
    InMux I__8365 (
            .O(N__37727),
            .I(N__37724));
    LocalMux I__8364 (
            .O(N__37724),
            .I(n4216));
    InMux I__8363 (
            .O(N__37721),
            .I(n14050));
    InMux I__8362 (
            .O(N__37718),
            .I(N__37715));
    LocalMux I__8361 (
            .O(N__37715),
            .I(N__37712));
    Span4Mux_v I__8360 (
            .O(N__37712),
            .I(N__37708));
    InMux I__8359 (
            .O(N__37711),
            .I(N__37705));
    Sp12to4 I__8358 (
            .O(N__37708),
            .I(N__37702));
    LocalMux I__8357 (
            .O(N__37705),
            .I(N__37699));
    Span12Mux_s11_h I__8356 (
            .O(N__37702),
            .I(N__37696));
    Span4Mux_h I__8355 (
            .O(N__37699),
            .I(N__37693));
    Odrv12 I__8354 (
            .O(N__37696),
            .I(n14_adj_1207));
    Odrv4 I__8353 (
            .O(N__37693),
            .I(n14_adj_1207));
    CascadeMux I__8352 (
            .O(N__37688),
            .I(N__37684));
    InMux I__8351 (
            .O(N__37687),
            .I(N__37681));
    InMux I__8350 (
            .O(N__37684),
            .I(N__37678));
    LocalMux I__8349 (
            .O(N__37681),
            .I(N__37675));
    LocalMux I__8348 (
            .O(N__37678),
            .I(data_idxvec_12));
    Odrv4 I__8347 (
            .O(N__37675),
            .I(data_idxvec_12));
    InMux I__8346 (
            .O(N__37670),
            .I(n14051));
    InMux I__8345 (
            .O(N__37667),
            .I(N__37664));
    LocalMux I__8344 (
            .O(N__37664),
            .I(N__37660));
    InMux I__8343 (
            .O(N__37663),
            .I(N__37657));
    Span4Mux_h I__8342 (
            .O(N__37660),
            .I(N__37654));
    LocalMux I__8341 (
            .O(N__37657),
            .I(n14_adj_1202));
    Odrv4 I__8340 (
            .O(N__37654),
            .I(n14_adj_1202));
    InMux I__8339 (
            .O(N__37649),
            .I(N__37645));
    InMux I__8338 (
            .O(N__37648),
            .I(N__37642));
    LocalMux I__8337 (
            .O(N__37645),
            .I(N__37639));
    LocalMux I__8336 (
            .O(N__37642),
            .I(data_idxvec_13));
    Odrv4 I__8335 (
            .O(N__37639),
            .I(data_idxvec_13));
    InMux I__8334 (
            .O(N__37634),
            .I(n14052));
    InMux I__8333 (
            .O(N__37631),
            .I(N__37627));
    InMux I__8332 (
            .O(N__37630),
            .I(N__37624));
    LocalMux I__8331 (
            .O(N__37627),
            .I(N__37621));
    LocalMux I__8330 (
            .O(N__37624),
            .I(N__37618));
    Span4Mux_h I__8329 (
            .O(N__37621),
            .I(N__37615));
    Odrv4 I__8328 (
            .O(N__37618),
            .I(n14_adj_1206));
    Odrv4 I__8327 (
            .O(N__37615),
            .I(n14_adj_1206));
    CascadeMux I__8326 (
            .O(N__37610),
            .I(N__37607));
    InMux I__8325 (
            .O(N__37607),
            .I(N__37603));
    CascadeMux I__8324 (
            .O(N__37606),
            .I(N__37600));
    LocalMux I__8323 (
            .O(N__37603),
            .I(N__37597));
    InMux I__8322 (
            .O(N__37600),
            .I(N__37594));
    Span12Mux_v I__8321 (
            .O(N__37597),
            .I(N__37591));
    LocalMux I__8320 (
            .O(N__37594),
            .I(data_idxvec_14));
    Odrv12 I__8319 (
            .O(N__37591),
            .I(data_idxvec_14));
    InMux I__8318 (
            .O(N__37586),
            .I(n14053));
    InMux I__8317 (
            .O(N__37583),
            .I(N__37579));
    InMux I__8316 (
            .O(N__37582),
            .I(N__37576));
    LocalMux I__8315 (
            .O(N__37579),
            .I(N__37573));
    LocalMux I__8314 (
            .O(N__37576),
            .I(N__37570));
    Span4Mux_h I__8313 (
            .O(N__37573),
            .I(N__37567));
    Span12Mux_h I__8312 (
            .O(N__37570),
            .I(N__37564));
    Odrv4 I__8311 (
            .O(N__37567),
            .I(n14_adj_1205));
    Odrv12 I__8310 (
            .O(N__37564),
            .I(n14_adj_1205));
    InMux I__8309 (
            .O(N__37559),
            .I(n14054));
    CEMux I__8308 (
            .O(N__37556),
            .I(N__37553));
    LocalMux I__8307 (
            .O(N__37553),
            .I(N__37549));
    CEMux I__8306 (
            .O(N__37552),
            .I(N__37546));
    Span4Mux_h I__8305 (
            .O(N__37549),
            .I(N__37542));
    LocalMux I__8304 (
            .O(N__37546),
            .I(N__37539));
    CEMux I__8303 (
            .O(N__37545),
            .I(N__37536));
    Sp12to4 I__8302 (
            .O(N__37542),
            .I(N__37533));
    Span4Mux_h I__8301 (
            .O(N__37539),
            .I(N__37530));
    LocalMux I__8300 (
            .O(N__37536),
            .I(N__37527));
    Odrv12 I__8299 (
            .O(N__37533),
            .I(n9187));
    Odrv4 I__8298 (
            .O(N__37530),
            .I(n9187));
    Odrv12 I__8297 (
            .O(N__37527),
            .I(n9187));
    InMux I__8296 (
            .O(N__37520),
            .I(N__37517));
    LocalMux I__8295 (
            .O(N__37517),
            .I(N__37513));
    InMux I__8294 (
            .O(N__37516),
            .I(N__37509));
    Span4Mux_h I__8293 (
            .O(N__37513),
            .I(N__37506));
    InMux I__8292 (
            .O(N__37512),
            .I(N__37503));
    LocalMux I__8291 (
            .O(N__37509),
            .I(buf_adcdata3_13));
    Odrv4 I__8290 (
            .O(N__37506),
            .I(buf_adcdata3_13));
    LocalMux I__8289 (
            .O(N__37503),
            .I(buf_adcdata3_13));
    InMux I__8288 (
            .O(N__37496),
            .I(N__37493));
    LocalMux I__8287 (
            .O(N__37493),
            .I(N__37489));
    InMux I__8286 (
            .O(N__37492),
            .I(N__37486));
    Span4Mux_v I__8285 (
            .O(N__37489),
            .I(N__37481));
    LocalMux I__8284 (
            .O(N__37486),
            .I(N__37481));
    Span4Mux_v I__8283 (
            .O(N__37481),
            .I(N__37478));
    Odrv4 I__8282 (
            .O(N__37478),
            .I(n14_adj_1198));
    CascadeMux I__8281 (
            .O(N__37475),
            .I(N__37472));
    InMux I__8280 (
            .O(N__37472),
            .I(N__37469));
    LocalMux I__8279 (
            .O(N__37469),
            .I(N__37466));
    Span4Mux_v I__8278 (
            .O(N__37466),
            .I(N__37463));
    Sp12to4 I__8277 (
            .O(N__37463),
            .I(N__37458));
    InMux I__8276 (
            .O(N__37462),
            .I(N__37453));
    InMux I__8275 (
            .O(N__37461),
            .I(N__37453));
    Span12Mux_h I__8274 (
            .O(N__37458),
            .I(N__37450));
    LocalMux I__8273 (
            .O(N__37453),
            .I(cmd_rdadctmp_22));
    Odrv12 I__8272 (
            .O(N__37450),
            .I(cmd_rdadctmp_22));
    InMux I__8271 (
            .O(N__37445),
            .I(N__37442));
    LocalMux I__8270 (
            .O(N__37442),
            .I(N__37438));
    InMux I__8269 (
            .O(N__37441),
            .I(N__37435));
    Span4Mux_h I__8268 (
            .O(N__37438),
            .I(N__37432));
    LocalMux I__8267 (
            .O(N__37435),
            .I(buf_adcdata1_14));
    Odrv4 I__8266 (
            .O(N__37432),
            .I(buf_adcdata1_14));
    InMux I__8265 (
            .O(N__37427),
            .I(N__37424));
    LocalMux I__8264 (
            .O(N__37424),
            .I(N__37419));
    InMux I__8263 (
            .O(N__37423),
            .I(N__37416));
    InMux I__8262 (
            .O(N__37422),
            .I(N__37413));
    Span4Mux_v I__8261 (
            .O(N__37419),
            .I(N__37408));
    LocalMux I__8260 (
            .O(N__37416),
            .I(N__37408));
    LocalMux I__8259 (
            .O(N__37413),
            .I(req_data_cnt_11));
    Odrv4 I__8258 (
            .O(N__37408),
            .I(req_data_cnt_11));
    InMux I__8257 (
            .O(N__37403),
            .I(n14042));
    InMux I__8256 (
            .O(N__37400),
            .I(N__37396));
    InMux I__8255 (
            .O(N__37399),
            .I(N__37393));
    LocalMux I__8254 (
            .O(N__37396),
            .I(N__37390));
    LocalMux I__8253 (
            .O(N__37393),
            .I(N__37387));
    Span4Mux_h I__8252 (
            .O(N__37390),
            .I(N__37384));
    Span4Mux_v I__8251 (
            .O(N__37387),
            .I(N__37381));
    Odrv4 I__8250 (
            .O(N__37384),
            .I(n14_adj_1196));
    Odrv4 I__8249 (
            .O(N__37381),
            .I(n14_adj_1196));
    InMux I__8248 (
            .O(N__37376),
            .I(n14043));
    InMux I__8247 (
            .O(N__37373),
            .I(N__37370));
    LocalMux I__8246 (
            .O(N__37370),
            .I(N__37366));
    InMux I__8245 (
            .O(N__37369),
            .I(N__37363));
    Span4Mux_h I__8244 (
            .O(N__37366),
            .I(N__37360));
    LocalMux I__8243 (
            .O(N__37363),
            .I(N__37357));
    Span4Mux_v I__8242 (
            .O(N__37360),
            .I(N__37354));
    Odrv4 I__8241 (
            .O(N__37357),
            .I(n14_adj_1213));
    Odrv4 I__8240 (
            .O(N__37354),
            .I(n14_adj_1213));
    InMux I__8239 (
            .O(N__37349),
            .I(n14044));
    InMux I__8238 (
            .O(N__37346),
            .I(N__37342));
    CascadeMux I__8237 (
            .O(N__37345),
            .I(N__37339));
    LocalMux I__8236 (
            .O(N__37342),
            .I(N__37336));
    InMux I__8235 (
            .O(N__37339),
            .I(N__37333));
    Span4Mux_h I__8234 (
            .O(N__37336),
            .I(N__37330));
    LocalMux I__8233 (
            .O(N__37333),
            .I(data_idxvec_6));
    Odrv4 I__8232 (
            .O(N__37330),
            .I(data_idxvec_6));
    InMux I__8231 (
            .O(N__37325),
            .I(n14045));
    InMux I__8230 (
            .O(N__37322),
            .I(N__37319));
    LocalMux I__8229 (
            .O(N__37319),
            .I(N__37315));
    InMux I__8228 (
            .O(N__37318),
            .I(N__37312));
    Span4Mux_h I__8227 (
            .O(N__37315),
            .I(N__37309));
    LocalMux I__8226 (
            .O(N__37312),
            .I(N__37304));
    Span4Mux_h I__8225 (
            .O(N__37309),
            .I(N__37304));
    Span4Mux_v I__8224 (
            .O(N__37304),
            .I(N__37301));
    Odrv4 I__8223 (
            .O(N__37301),
            .I(n14_adj_1168));
    InMux I__8222 (
            .O(N__37298),
            .I(N__37295));
    LocalMux I__8221 (
            .O(N__37295),
            .I(N__37291));
    InMux I__8220 (
            .O(N__37294),
            .I(N__37288));
    Span4Mux_h I__8219 (
            .O(N__37291),
            .I(N__37285));
    LocalMux I__8218 (
            .O(N__37288),
            .I(data_idxvec_7));
    Odrv4 I__8217 (
            .O(N__37285),
            .I(data_idxvec_7));
    InMux I__8216 (
            .O(N__37280),
            .I(n14046));
    InMux I__8215 (
            .O(N__37277),
            .I(N__37274));
    LocalMux I__8214 (
            .O(N__37274),
            .I(N__37269));
    InMux I__8213 (
            .O(N__37273),
            .I(N__37266));
    InMux I__8212 (
            .O(N__37272),
            .I(N__37263));
    Span4Mux_v I__8211 (
            .O(N__37269),
            .I(N__37260));
    LocalMux I__8210 (
            .O(N__37266),
            .I(N__37255));
    LocalMux I__8209 (
            .O(N__37263),
            .I(N__37255));
    Span4Mux_h I__8208 (
            .O(N__37260),
            .I(N__37252));
    Span4Mux_v I__8207 (
            .O(N__37255),
            .I(N__37249));
    Sp12to4 I__8206 (
            .O(N__37252),
            .I(N__37246));
    Odrv4 I__8205 (
            .O(N__37249),
            .I(n14_adj_1211));
    Odrv12 I__8204 (
            .O(N__37246),
            .I(n14_adj_1211));
    InMux I__8203 (
            .O(N__37241),
            .I(bfn_17_13_0_));
    InMux I__8202 (
            .O(N__37238),
            .I(N__37234));
    InMux I__8201 (
            .O(N__37237),
            .I(N__37231));
    LocalMux I__8200 (
            .O(N__37234),
            .I(N__37228));
    LocalMux I__8199 (
            .O(N__37231),
            .I(N__37225));
    Span12Mux_v I__8198 (
            .O(N__37228),
            .I(N__37222));
    Span4Mux_v I__8197 (
            .O(N__37225),
            .I(N__37219));
    Odrv12 I__8196 (
            .O(N__37222),
            .I(n14_adj_1210));
    Odrv4 I__8195 (
            .O(N__37219),
            .I(n14_adj_1210));
    CascadeMux I__8194 (
            .O(N__37214),
            .I(N__37211));
    InMux I__8193 (
            .O(N__37211),
            .I(N__37208));
    LocalMux I__8192 (
            .O(N__37208),
            .I(N__37204));
    InMux I__8191 (
            .O(N__37207),
            .I(N__37201));
    Span4Mux_h I__8190 (
            .O(N__37204),
            .I(N__37198));
    LocalMux I__8189 (
            .O(N__37201),
            .I(data_idxvec_9));
    Odrv4 I__8188 (
            .O(N__37198),
            .I(data_idxvec_9));
    InMux I__8187 (
            .O(N__37193),
            .I(n14048));
    InMux I__8186 (
            .O(N__37190),
            .I(N__37186));
    InMux I__8185 (
            .O(N__37189),
            .I(N__37183));
    LocalMux I__8184 (
            .O(N__37186),
            .I(N__37180));
    LocalMux I__8183 (
            .O(N__37183),
            .I(N__37177));
    Span4Mux_h I__8182 (
            .O(N__37180),
            .I(N__37172));
    Span4Mux_h I__8181 (
            .O(N__37177),
            .I(N__37172));
    Odrv4 I__8180 (
            .O(N__37172),
            .I(n14_adj_1209));
    CascadeMux I__8179 (
            .O(N__37169),
            .I(N__37165));
    CascadeMux I__8178 (
            .O(N__37168),
            .I(N__37162));
    InMux I__8177 (
            .O(N__37165),
            .I(N__37159));
    InMux I__8176 (
            .O(N__37162),
            .I(N__37156));
    LocalMux I__8175 (
            .O(N__37159),
            .I(N__37153));
    LocalMux I__8174 (
            .O(N__37156),
            .I(data_idxvec_10));
    Odrv4 I__8173 (
            .O(N__37153),
            .I(data_idxvec_10));
    InMux I__8172 (
            .O(N__37148),
            .I(n14049));
    InMux I__8171 (
            .O(N__37145),
            .I(N__37142));
    LocalMux I__8170 (
            .O(N__37142),
            .I(N__37139));
    Span4Mux_v I__8169 (
            .O(N__37139),
            .I(N__37136));
    Span4Mux_v I__8168 (
            .O(N__37136),
            .I(N__37133));
    Span4Mux_h I__8167 (
            .O(N__37133),
            .I(N__37130));
    Odrv4 I__8166 (
            .O(N__37130),
            .I(buf_data1_8));
    CascadeMux I__8165 (
            .O(N__37127),
            .I(n4197_cascade_));
    InMux I__8164 (
            .O(N__37124),
            .I(N__37121));
    LocalMux I__8163 (
            .O(N__37121),
            .I(N__37118));
    Span4Mux_h I__8162 (
            .O(N__37118),
            .I(N__37115));
    Odrv4 I__8161 (
            .O(N__37115),
            .I(n4221));
    CascadeMux I__8160 (
            .O(N__37112),
            .I(n4234_cascade_));
    InMux I__8159 (
            .O(N__37109),
            .I(N__37106));
    LocalMux I__8158 (
            .O(N__37106),
            .I(N__37103));
    Span4Mux_v I__8157 (
            .O(N__37103),
            .I(N__37100));
    Span4Mux_h I__8156 (
            .O(N__37100),
            .I(N__37097));
    Span4Mux_h I__8155 (
            .O(N__37097),
            .I(N__37094));
    Odrv4 I__8154 (
            .O(N__37094),
            .I(n4209));
    CascadeMux I__8153 (
            .O(N__37091),
            .I(n4254_cascade_));
    InMux I__8152 (
            .O(N__37088),
            .I(N__37085));
    LocalMux I__8151 (
            .O(N__37085),
            .I(n4264));
    CascadeMux I__8150 (
            .O(N__37082),
            .I(n32_cascade_));
    InMux I__8149 (
            .O(N__37079),
            .I(N__37076));
    LocalMux I__8148 (
            .O(N__37076),
            .I(N__37073));
    Span4Mux_h I__8147 (
            .O(N__37073),
            .I(N__37070));
    Span4Mux_h I__8146 (
            .O(N__37070),
            .I(N__37067));
    Odrv4 I__8145 (
            .O(N__37067),
            .I(n15557));
    CascadeMux I__8144 (
            .O(N__37064),
            .I(N__37061));
    InMux I__8143 (
            .O(N__37061),
            .I(N__37057));
    InMux I__8142 (
            .O(N__37060),
            .I(N__37054));
    LocalMux I__8141 (
            .O(N__37057),
            .I(data_idxvec_0));
    LocalMux I__8140 (
            .O(N__37054),
            .I(data_idxvec_0));
    InMux I__8139 (
            .O(N__37049),
            .I(N__37046));
    LocalMux I__8138 (
            .O(N__37046),
            .I(data_idxvec_15_N_673_0));
    InMux I__8137 (
            .O(N__37043),
            .I(n14040));
    CascadeMux I__8136 (
            .O(N__37040),
            .I(N__37036));
    InMux I__8135 (
            .O(N__37039),
            .I(N__37033));
    InMux I__8134 (
            .O(N__37036),
            .I(N__37030));
    LocalMux I__8133 (
            .O(N__37033),
            .I(N__37027));
    LocalMux I__8132 (
            .O(N__37030),
            .I(N__37022));
    Span4Mux_v I__8131 (
            .O(N__37027),
            .I(N__37022));
    Odrv4 I__8130 (
            .O(N__37022),
            .I(data_idxvec_2));
    InMux I__8129 (
            .O(N__37019),
            .I(n14041));
    CascadeMux I__8128 (
            .O(N__37016),
            .I(N__37013));
    InMux I__8127 (
            .O(N__37013),
            .I(N__37010));
    LocalMux I__8126 (
            .O(N__37010),
            .I(N__37007));
    Span4Mux_h I__8125 (
            .O(N__37007),
            .I(N__37004));
    Span4Mux_v I__8124 (
            .O(N__37004),
            .I(N__37001));
    Odrv4 I__8123 (
            .O(N__37001),
            .I(buf_data1_20));
    CascadeMux I__8122 (
            .O(N__36998),
            .I(n8058_cascade_));
    InMux I__8121 (
            .O(N__36995),
            .I(N__36991));
    InMux I__8120 (
            .O(N__36994),
            .I(N__36986));
    LocalMux I__8119 (
            .O(N__36991),
            .I(N__36983));
    InMux I__8118 (
            .O(N__36990),
            .I(N__36980));
    CascadeMux I__8117 (
            .O(N__36989),
            .I(N__36977));
    LocalMux I__8116 (
            .O(N__36986),
            .I(N__36974));
    Span4Mux_v I__8115 (
            .O(N__36983),
            .I(N__36969));
    LocalMux I__8114 (
            .O(N__36980),
            .I(N__36964));
    InMux I__8113 (
            .O(N__36977),
            .I(N__36961));
    Span4Mux_v I__8112 (
            .O(N__36974),
            .I(N__36957));
    InMux I__8111 (
            .O(N__36973),
            .I(N__36954));
    CascadeMux I__8110 (
            .O(N__36972),
            .I(N__36951));
    Span4Mux_h I__8109 (
            .O(N__36969),
            .I(N__36948));
    InMux I__8108 (
            .O(N__36968),
            .I(N__36943));
    InMux I__8107 (
            .O(N__36967),
            .I(N__36943));
    Span4Mux_v I__8106 (
            .O(N__36964),
            .I(N__36940));
    LocalMux I__8105 (
            .O(N__36961),
            .I(N__36937));
    InMux I__8104 (
            .O(N__36960),
            .I(N__36934));
    Span4Mux_h I__8103 (
            .O(N__36957),
            .I(N__36929));
    LocalMux I__8102 (
            .O(N__36954),
            .I(N__36929));
    InMux I__8101 (
            .O(N__36951),
            .I(N__36926));
    Span4Mux_h I__8100 (
            .O(N__36948),
            .I(N__36923));
    LocalMux I__8099 (
            .O(N__36943),
            .I(N__36920));
    Span4Mux_h I__8098 (
            .O(N__36940),
            .I(N__36915));
    Span4Mux_v I__8097 (
            .O(N__36937),
            .I(N__36915));
    LocalMux I__8096 (
            .O(N__36934),
            .I(N__36908));
    Sp12to4 I__8095 (
            .O(N__36929),
            .I(N__36908));
    LocalMux I__8094 (
            .O(N__36926),
            .I(N__36908));
    Span4Mux_v I__8093 (
            .O(N__36923),
            .I(N__36903));
    Span4Mux_h I__8092 (
            .O(N__36920),
            .I(N__36903));
    Odrv4 I__8091 (
            .O(N__36915),
            .I(comm_buf_0_4));
    Odrv12 I__8090 (
            .O(N__36908),
            .I(comm_buf_0_4));
    Odrv4 I__8089 (
            .O(N__36903),
            .I(comm_buf_0_4));
    InMux I__8088 (
            .O(N__36896),
            .I(N__36893));
    LocalMux I__8087 (
            .O(N__36893),
            .I(n15584));
    CascadeMux I__8086 (
            .O(N__36890),
            .I(n83_cascade_));
    InMux I__8085 (
            .O(N__36887),
            .I(N__36884));
    LocalMux I__8084 (
            .O(N__36884),
            .I(N__36881));
    Odrv12 I__8083 (
            .O(N__36881),
            .I(n15581));
    InMux I__8082 (
            .O(N__36878),
            .I(N__36874));
    InMux I__8081 (
            .O(N__36877),
            .I(N__36871));
    LocalMux I__8080 (
            .O(N__36874),
            .I(N__36868));
    LocalMux I__8079 (
            .O(N__36871),
            .I(N__36865));
    Span4Mux_h I__8078 (
            .O(N__36868),
            .I(N__36862));
    Span12Mux_v I__8077 (
            .O(N__36865),
            .I(N__36858));
    Span4Mux_h I__8076 (
            .O(N__36862),
            .I(N__36855));
    InMux I__8075 (
            .O(N__36861),
            .I(N__36852));
    Odrv12 I__8074 (
            .O(N__36858),
            .I(cmd_rdadctmp_29_adj_1083));
    Odrv4 I__8073 (
            .O(N__36855),
            .I(cmd_rdadctmp_29_adj_1083));
    LocalMux I__8072 (
            .O(N__36852),
            .I(cmd_rdadctmp_29_adj_1083));
    InMux I__8071 (
            .O(N__36845),
            .I(N__36840));
    CascadeMux I__8070 (
            .O(N__36844),
            .I(N__36837));
    InMux I__8069 (
            .O(N__36843),
            .I(N__36834));
    LocalMux I__8068 (
            .O(N__36840),
            .I(N__36831));
    InMux I__8067 (
            .O(N__36837),
            .I(N__36828));
    LocalMux I__8066 (
            .O(N__36834),
            .I(N__36825));
    Span4Mux_v I__8065 (
            .O(N__36831),
            .I(N__36822));
    LocalMux I__8064 (
            .O(N__36828),
            .I(N__36817));
    Span4Mux_v I__8063 (
            .O(N__36825),
            .I(N__36817));
    Span4Mux_h I__8062 (
            .O(N__36822),
            .I(N__36814));
    Sp12to4 I__8061 (
            .O(N__36817),
            .I(N__36811));
    Odrv4 I__8060 (
            .O(N__36814),
            .I(buf_adcdata3_21));
    Odrv12 I__8059 (
            .O(N__36811),
            .I(buf_adcdata3_21));
    CascadeMux I__8058 (
            .O(N__36806),
            .I(N__36803));
    InMux I__8057 (
            .O(N__36803),
            .I(N__36800));
    LocalMux I__8056 (
            .O(N__36800),
            .I(N__36797));
    Span4Mux_v I__8055 (
            .O(N__36797),
            .I(N__36794));
    Span4Mux_h I__8054 (
            .O(N__36794),
            .I(N__36790));
    CascadeMux I__8053 (
            .O(N__36793),
            .I(N__36786));
    Span4Mux_v I__8052 (
            .O(N__36790),
            .I(N__36783));
    InMux I__8051 (
            .O(N__36789),
            .I(N__36780));
    InMux I__8050 (
            .O(N__36786),
            .I(N__36777));
    Odrv4 I__8049 (
            .O(N__36783),
            .I(cmd_rdadctmp_23_adj_1089));
    LocalMux I__8048 (
            .O(N__36780),
            .I(cmd_rdadctmp_23_adj_1089));
    LocalMux I__8047 (
            .O(N__36777),
            .I(cmd_rdadctmp_23_adj_1089));
    InMux I__8046 (
            .O(N__36770),
            .I(N__36767));
    LocalMux I__8045 (
            .O(N__36767),
            .I(N__36764));
    Span4Mux_v I__8044 (
            .O(N__36764),
            .I(N__36759));
    InMux I__8043 (
            .O(N__36763),
            .I(N__36756));
    InMux I__8042 (
            .O(N__36762),
            .I(N__36753));
    Span4Mux_h I__8041 (
            .O(N__36759),
            .I(N__36748));
    LocalMux I__8040 (
            .O(N__36756),
            .I(N__36748));
    LocalMux I__8039 (
            .O(N__36753),
            .I(buf_adcdata3_15));
    Odrv4 I__8038 (
            .O(N__36748),
            .I(buf_adcdata3_15));
    InMux I__8037 (
            .O(N__36743),
            .I(N__36740));
    LocalMux I__8036 (
            .O(N__36740),
            .I(N__36737));
    Odrv12 I__8035 (
            .O(N__36737),
            .I(buf_data1_18));
    CascadeMux I__8034 (
            .O(N__36734),
            .I(N__36731));
    InMux I__8033 (
            .O(N__36731),
            .I(N__36728));
    LocalMux I__8032 (
            .O(N__36728),
            .I(N__36725));
    Span4Mux_h I__8031 (
            .O(N__36725),
            .I(N__36722));
    Span4Mux_h I__8030 (
            .O(N__36722),
            .I(N__36719));
    Odrv4 I__8029 (
            .O(N__36719),
            .I(n75_adj_1164));
    InMux I__8028 (
            .O(N__36716),
            .I(N__36709));
    InMux I__8027 (
            .O(N__36715),
            .I(N__36706));
    InMux I__8026 (
            .O(N__36714),
            .I(N__36702));
    InMux I__8025 (
            .O(N__36713),
            .I(N__36699));
    InMux I__8024 (
            .O(N__36712),
            .I(N__36696));
    LocalMux I__8023 (
            .O(N__36709),
            .I(N__36693));
    LocalMux I__8022 (
            .O(N__36706),
            .I(N__36690));
    CascadeMux I__8021 (
            .O(N__36705),
            .I(N__36687));
    LocalMux I__8020 (
            .O(N__36702),
            .I(N__36684));
    LocalMux I__8019 (
            .O(N__36699),
            .I(N__36681));
    LocalMux I__8018 (
            .O(N__36696),
            .I(N__36678));
    Span4Mux_h I__8017 (
            .O(N__36693),
            .I(N__36673));
    Span4Mux_h I__8016 (
            .O(N__36690),
            .I(N__36673));
    InMux I__8015 (
            .O(N__36687),
            .I(N__36670));
    Span4Mux_v I__8014 (
            .O(N__36684),
            .I(N__36667));
    Span4Mux_v I__8013 (
            .O(N__36681),
            .I(N__36662));
    Span4Mux_h I__8012 (
            .O(N__36678),
            .I(N__36662));
    Odrv4 I__8011 (
            .O(N__36673),
            .I(comm_buf_1_0));
    LocalMux I__8010 (
            .O(N__36670),
            .I(comm_buf_1_0));
    Odrv4 I__8009 (
            .O(N__36667),
            .I(comm_buf_1_0));
    Odrv4 I__8008 (
            .O(N__36662),
            .I(comm_buf_1_0));
    InMux I__8007 (
            .O(N__36653),
            .I(N__36650));
    LocalMux I__8006 (
            .O(N__36650),
            .I(N__36645));
    InMux I__8005 (
            .O(N__36649),
            .I(N__36642));
    InMux I__8004 (
            .O(N__36648),
            .I(N__36639));
    Span4Mux_v I__8003 (
            .O(N__36645),
            .I(N__36636));
    LocalMux I__8002 (
            .O(N__36642),
            .I(data_cntvec_0));
    LocalMux I__8001 (
            .O(N__36639),
            .I(data_cntvec_0));
    Odrv4 I__8000 (
            .O(N__36636),
            .I(data_cntvec_0));
    InMux I__7999 (
            .O(N__36629),
            .I(N__36626));
    LocalMux I__7998 (
            .O(N__36626),
            .I(N__36623));
    Odrv4 I__7997 (
            .O(N__36623),
            .I(n15527));
    CEMux I__7996 (
            .O(N__36620),
            .I(N__36617));
    LocalMux I__7995 (
            .O(N__36617),
            .I(N__36614));
    Span4Mux_h I__7994 (
            .O(N__36614),
            .I(N__36611));
    Span4Mux_h I__7993 (
            .O(N__36611),
            .I(N__36608));
    Odrv4 I__7992 (
            .O(N__36608),
            .I(n14_adj_1189));
    InMux I__7991 (
            .O(N__36605),
            .I(N__36602));
    LocalMux I__7990 (
            .O(N__36602),
            .I(n13_adj_1032));
    CascadeMux I__7989 (
            .O(N__36599),
            .I(n13_adj_1032_cascade_));
    InMux I__7988 (
            .O(N__36596),
            .I(N__36590));
    InMux I__7987 (
            .O(N__36595),
            .I(N__36590));
    LocalMux I__7986 (
            .O(N__36590),
            .I(n8519));
    InMux I__7985 (
            .O(N__36587),
            .I(N__36583));
    InMux I__7984 (
            .O(N__36586),
            .I(N__36580));
    LocalMux I__7983 (
            .O(N__36583),
            .I(N__36577));
    LocalMux I__7982 (
            .O(N__36580),
            .I(N__36574));
    Span12Mux_h I__7981 (
            .O(N__36577),
            .I(N__36571));
    Odrv4 I__7980 (
            .O(N__36574),
            .I(n22_adj_1115));
    Odrv12 I__7979 (
            .O(N__36571),
            .I(n22_adj_1115));
    CascadeMux I__7978 (
            .O(N__36566),
            .I(N__36563));
    InMux I__7977 (
            .O(N__36563),
            .I(N__36560));
    LocalMux I__7976 (
            .O(N__36560),
            .I(n15651));
    InMux I__7975 (
            .O(N__36557),
            .I(N__36554));
    LocalMux I__7974 (
            .O(N__36554),
            .I(n15526));
    CascadeMux I__7973 (
            .O(N__36551),
            .I(n15668_cascade_));
    InMux I__7972 (
            .O(N__36548),
            .I(N__36545));
    LocalMux I__7971 (
            .O(N__36545),
            .I(n1523));
    CascadeMux I__7970 (
            .O(N__36542),
            .I(n1523_cascade_));
    CascadeMux I__7969 (
            .O(N__36539),
            .I(n2_adj_1200_cascade_));
    InMux I__7968 (
            .O(N__36536),
            .I(N__36533));
    LocalMux I__7967 (
            .O(N__36533),
            .I(n16464));
    CascadeMux I__7966 (
            .O(N__36530),
            .I(n16467_cascade_));
    InMux I__7965 (
            .O(N__36527),
            .I(N__36524));
    LocalMux I__7964 (
            .O(N__36524),
            .I(n8_adj_1201));
    SRMux I__7963 (
            .O(N__36521),
            .I(N__36518));
    LocalMux I__7962 (
            .O(N__36518),
            .I(N__36515));
    Span4Mux_h I__7961 (
            .O(N__36515),
            .I(N__36512));
    Odrv4 I__7960 (
            .O(N__36512),
            .I(\ADC_VAC2.n14926 ));
    InMux I__7959 (
            .O(N__36509),
            .I(N__36506));
    LocalMux I__7958 (
            .O(N__36506),
            .I(N__36502));
    CEMux I__7957 (
            .O(N__36505),
            .I(N__36499));
    Sp12to4 I__7956 (
            .O(N__36502),
            .I(N__36496));
    LocalMux I__7955 (
            .O(N__36499),
            .I(N__36493));
    Span12Mux_v I__7954 (
            .O(N__36496),
            .I(N__36490));
    Odrv4 I__7953 (
            .O(N__36493),
            .I(\ADC_VAC2.n9413 ));
    Odrv12 I__7952 (
            .O(N__36490),
            .I(\ADC_VAC2.n9413 ));
    InMux I__7951 (
            .O(N__36485),
            .I(N__36479));
    InMux I__7950 (
            .O(N__36484),
            .I(N__36479));
    LocalMux I__7949 (
            .O(N__36479),
            .I(N__36476));
    Span4Mux_h I__7948 (
            .O(N__36476),
            .I(N__36471));
    InMux I__7947 (
            .O(N__36475),
            .I(N__36467));
    InMux I__7946 (
            .O(N__36474),
            .I(N__36463));
    Span4Mux_h I__7945 (
            .O(N__36471),
            .I(N__36460));
    CascadeMux I__7944 (
            .O(N__36470),
            .I(N__36457));
    LocalMux I__7943 (
            .O(N__36467),
            .I(N__36453));
    InMux I__7942 (
            .O(N__36466),
            .I(N__36450));
    LocalMux I__7941 (
            .O(N__36463),
            .I(N__36446));
    Span4Mux_v I__7940 (
            .O(N__36460),
            .I(N__36443));
    InMux I__7939 (
            .O(N__36457),
            .I(N__36438));
    InMux I__7938 (
            .O(N__36456),
            .I(N__36438));
    Span4Mux_v I__7937 (
            .O(N__36453),
            .I(N__36435));
    LocalMux I__7936 (
            .O(N__36450),
            .I(N__36430));
    InMux I__7935 (
            .O(N__36449),
            .I(N__36425));
    Span4Mux_v I__7934 (
            .O(N__36446),
            .I(N__36416));
    Span4Mux_v I__7933 (
            .O(N__36443),
            .I(N__36416));
    LocalMux I__7932 (
            .O(N__36438),
            .I(N__36416));
    Span4Mux_h I__7931 (
            .O(N__36435),
            .I(N__36416));
    InMux I__7930 (
            .O(N__36434),
            .I(N__36411));
    InMux I__7929 (
            .O(N__36433),
            .I(N__36411));
    Span4Mux_h I__7928 (
            .O(N__36430),
            .I(N__36407));
    InMux I__7927 (
            .O(N__36429),
            .I(N__36404));
    InMux I__7926 (
            .O(N__36428),
            .I(N__36401));
    LocalMux I__7925 (
            .O(N__36425),
            .I(N__36398));
    Sp12to4 I__7924 (
            .O(N__36416),
            .I(N__36393));
    LocalMux I__7923 (
            .O(N__36411),
            .I(N__36393));
    InMux I__7922 (
            .O(N__36410),
            .I(N__36390));
    Odrv4 I__7921 (
            .O(N__36407),
            .I(DTRIG_N_957_adj_1077));
    LocalMux I__7920 (
            .O(N__36404),
            .I(DTRIG_N_957_adj_1077));
    LocalMux I__7919 (
            .O(N__36401),
            .I(DTRIG_N_957_adj_1077));
    Odrv4 I__7918 (
            .O(N__36398),
            .I(DTRIG_N_957_adj_1077));
    Odrv12 I__7917 (
            .O(N__36393),
            .I(DTRIG_N_957_adj_1077));
    LocalMux I__7916 (
            .O(N__36390),
            .I(DTRIG_N_957_adj_1077));
    SRMux I__7915 (
            .O(N__36377),
            .I(N__36374));
    LocalMux I__7914 (
            .O(N__36374),
            .I(N__36371));
    Span4Mux_h I__7913 (
            .O(N__36371),
            .I(N__36368));
    Span4Mux_h I__7912 (
            .O(N__36368),
            .I(N__36365));
    Span4Mux_v I__7911 (
            .O(N__36365),
            .I(N__36362));
    Odrv4 I__7910 (
            .O(N__36362),
            .I(\ADC_VAC2.n10706 ));
    InMux I__7909 (
            .O(N__36359),
            .I(N__36352));
    InMux I__7908 (
            .O(N__36358),
            .I(N__36352));
    InMux I__7907 (
            .O(N__36357),
            .I(N__36349));
    LocalMux I__7906 (
            .O(N__36352),
            .I(\comm_spi.bit_cnt_2 ));
    LocalMux I__7905 (
            .O(N__36349),
            .I(\comm_spi.bit_cnt_2 ));
    InMux I__7904 (
            .O(N__36344),
            .I(N__36334));
    InMux I__7903 (
            .O(N__36343),
            .I(N__36334));
    InMux I__7902 (
            .O(N__36342),
            .I(N__36334));
    InMux I__7901 (
            .O(N__36341),
            .I(N__36331));
    LocalMux I__7900 (
            .O(N__36334),
            .I(\comm_spi.bit_cnt_1 ));
    LocalMux I__7899 (
            .O(N__36331),
            .I(\comm_spi.bit_cnt_1 ));
    CascadeMux I__7898 (
            .O(N__36326),
            .I(N__36323));
    InMux I__7897 (
            .O(N__36323),
            .I(N__36310));
    InMux I__7896 (
            .O(N__36322),
            .I(N__36310));
    InMux I__7895 (
            .O(N__36321),
            .I(N__36310));
    InMux I__7894 (
            .O(N__36320),
            .I(N__36310));
    InMux I__7893 (
            .O(N__36319),
            .I(N__36307));
    LocalMux I__7892 (
            .O(N__36310),
            .I(\comm_spi.bit_cnt_0 ));
    LocalMux I__7891 (
            .O(N__36307),
            .I(\comm_spi.bit_cnt_0 ));
    CascadeMux I__7890 (
            .O(N__36302),
            .I(N__36299));
    CascadeBuf I__7889 (
            .O(N__36299),
            .I(N__36296));
    CascadeMux I__7888 (
            .O(N__36296),
            .I(N__36293));
    CascadeBuf I__7887 (
            .O(N__36293),
            .I(N__36290));
    CascadeMux I__7886 (
            .O(N__36290),
            .I(N__36287));
    CascadeBuf I__7885 (
            .O(N__36287),
            .I(N__36284));
    CascadeMux I__7884 (
            .O(N__36284),
            .I(N__36281));
    CascadeBuf I__7883 (
            .O(N__36281),
            .I(N__36278));
    CascadeMux I__7882 (
            .O(N__36278),
            .I(N__36275));
    CascadeBuf I__7881 (
            .O(N__36275),
            .I(N__36272));
    CascadeMux I__7880 (
            .O(N__36272),
            .I(N__36269));
    CascadeBuf I__7879 (
            .O(N__36269),
            .I(N__36266));
    CascadeMux I__7878 (
            .O(N__36266),
            .I(N__36263));
    CascadeBuf I__7877 (
            .O(N__36263),
            .I(N__36259));
    CascadeMux I__7876 (
            .O(N__36262),
            .I(N__36256));
    CascadeMux I__7875 (
            .O(N__36259),
            .I(N__36253));
    CascadeBuf I__7874 (
            .O(N__36256),
            .I(N__36250));
    CascadeBuf I__7873 (
            .O(N__36253),
            .I(N__36247));
    CascadeMux I__7872 (
            .O(N__36250),
            .I(N__36244));
    CascadeMux I__7871 (
            .O(N__36247),
            .I(N__36241));
    InMux I__7870 (
            .O(N__36244),
            .I(N__36238));
    CascadeBuf I__7869 (
            .O(N__36241),
            .I(N__36235));
    LocalMux I__7868 (
            .O(N__36238),
            .I(N__36232));
    CascadeMux I__7867 (
            .O(N__36235),
            .I(N__36229));
    Span4Mux_h I__7866 (
            .O(N__36232),
            .I(N__36226));
    InMux I__7865 (
            .O(N__36229),
            .I(N__36223));
    Span4Mux_v I__7864 (
            .O(N__36226),
            .I(N__36220));
    LocalMux I__7863 (
            .O(N__36223),
            .I(N__36217));
    Sp12to4 I__7862 (
            .O(N__36220),
            .I(N__36213));
    Span4Mux_h I__7861 (
            .O(N__36217),
            .I(N__36210));
    InMux I__7860 (
            .O(N__36216),
            .I(N__36207));
    Span12Mux_v I__7859 (
            .O(N__36213),
            .I(N__36204));
    Span4Mux_h I__7858 (
            .O(N__36210),
            .I(N__36201));
    LocalMux I__7857 (
            .O(N__36207),
            .I(data_count_4));
    Odrv12 I__7856 (
            .O(N__36204),
            .I(data_count_4));
    Odrv4 I__7855 (
            .O(N__36201),
            .I(data_count_4));
    InMux I__7854 (
            .O(N__36194),
            .I(n13945));
    CascadeMux I__7853 (
            .O(N__36191),
            .I(N__36188));
    CascadeBuf I__7852 (
            .O(N__36188),
            .I(N__36185));
    CascadeMux I__7851 (
            .O(N__36185),
            .I(N__36182));
    CascadeBuf I__7850 (
            .O(N__36182),
            .I(N__36179));
    CascadeMux I__7849 (
            .O(N__36179),
            .I(N__36176));
    CascadeBuf I__7848 (
            .O(N__36176),
            .I(N__36173));
    CascadeMux I__7847 (
            .O(N__36173),
            .I(N__36170));
    CascadeBuf I__7846 (
            .O(N__36170),
            .I(N__36167));
    CascadeMux I__7845 (
            .O(N__36167),
            .I(N__36164));
    CascadeBuf I__7844 (
            .O(N__36164),
            .I(N__36161));
    CascadeMux I__7843 (
            .O(N__36161),
            .I(N__36158));
    CascadeBuf I__7842 (
            .O(N__36158),
            .I(N__36155));
    CascadeMux I__7841 (
            .O(N__36155),
            .I(N__36152));
    CascadeBuf I__7840 (
            .O(N__36152),
            .I(N__36149));
    CascadeMux I__7839 (
            .O(N__36149),
            .I(N__36145));
    CascadeMux I__7838 (
            .O(N__36148),
            .I(N__36142));
    CascadeBuf I__7837 (
            .O(N__36145),
            .I(N__36139));
    CascadeBuf I__7836 (
            .O(N__36142),
            .I(N__36136));
    CascadeMux I__7835 (
            .O(N__36139),
            .I(N__36133));
    CascadeMux I__7834 (
            .O(N__36136),
            .I(N__36130));
    CascadeBuf I__7833 (
            .O(N__36133),
            .I(N__36127));
    InMux I__7832 (
            .O(N__36130),
            .I(N__36124));
    CascadeMux I__7831 (
            .O(N__36127),
            .I(N__36121));
    LocalMux I__7830 (
            .O(N__36124),
            .I(N__36118));
    InMux I__7829 (
            .O(N__36121),
            .I(N__36115));
    Span4Mux_v I__7828 (
            .O(N__36118),
            .I(N__36112));
    LocalMux I__7827 (
            .O(N__36115),
            .I(N__36109));
    Sp12to4 I__7826 (
            .O(N__36112),
            .I(N__36105));
    Span4Mux_h I__7825 (
            .O(N__36109),
            .I(N__36102));
    InMux I__7824 (
            .O(N__36108),
            .I(N__36099));
    Span12Mux_h I__7823 (
            .O(N__36105),
            .I(N__36096));
    Span4Mux_h I__7822 (
            .O(N__36102),
            .I(N__36093));
    LocalMux I__7821 (
            .O(N__36099),
            .I(data_count_5));
    Odrv12 I__7820 (
            .O(N__36096),
            .I(data_count_5));
    Odrv4 I__7819 (
            .O(N__36093),
            .I(data_count_5));
    InMux I__7818 (
            .O(N__36086),
            .I(n13946));
    CascadeMux I__7817 (
            .O(N__36083),
            .I(N__36080));
    CascadeBuf I__7816 (
            .O(N__36080),
            .I(N__36077));
    CascadeMux I__7815 (
            .O(N__36077),
            .I(N__36074));
    CascadeBuf I__7814 (
            .O(N__36074),
            .I(N__36071));
    CascadeMux I__7813 (
            .O(N__36071),
            .I(N__36068));
    CascadeBuf I__7812 (
            .O(N__36068),
            .I(N__36065));
    CascadeMux I__7811 (
            .O(N__36065),
            .I(N__36062));
    CascadeBuf I__7810 (
            .O(N__36062),
            .I(N__36059));
    CascadeMux I__7809 (
            .O(N__36059),
            .I(N__36056));
    CascadeBuf I__7808 (
            .O(N__36056),
            .I(N__36053));
    CascadeMux I__7807 (
            .O(N__36053),
            .I(N__36050));
    CascadeBuf I__7806 (
            .O(N__36050),
            .I(N__36047));
    CascadeMux I__7805 (
            .O(N__36047),
            .I(N__36044));
    CascadeBuf I__7804 (
            .O(N__36044),
            .I(N__36041));
    CascadeMux I__7803 (
            .O(N__36041),
            .I(N__36037));
    CascadeMux I__7802 (
            .O(N__36040),
            .I(N__36034));
    CascadeBuf I__7801 (
            .O(N__36037),
            .I(N__36031));
    CascadeBuf I__7800 (
            .O(N__36034),
            .I(N__36028));
    CascadeMux I__7799 (
            .O(N__36031),
            .I(N__36025));
    CascadeMux I__7798 (
            .O(N__36028),
            .I(N__36022));
    CascadeBuf I__7797 (
            .O(N__36025),
            .I(N__36019));
    InMux I__7796 (
            .O(N__36022),
            .I(N__36016));
    CascadeMux I__7795 (
            .O(N__36019),
            .I(N__36013));
    LocalMux I__7794 (
            .O(N__36016),
            .I(N__36010));
    InMux I__7793 (
            .O(N__36013),
            .I(N__36007));
    Sp12to4 I__7792 (
            .O(N__36010),
            .I(N__36004));
    LocalMux I__7791 (
            .O(N__36007),
            .I(N__36001));
    Span12Mux_v I__7790 (
            .O(N__36004),
            .I(N__35997));
    Span4Mux_h I__7789 (
            .O(N__36001),
            .I(N__35994));
    InMux I__7788 (
            .O(N__36000),
            .I(N__35991));
    Span12Mux_h I__7787 (
            .O(N__35997),
            .I(N__35988));
    Span4Mux_h I__7786 (
            .O(N__35994),
            .I(N__35985));
    LocalMux I__7785 (
            .O(N__35991),
            .I(data_count_6));
    Odrv12 I__7784 (
            .O(N__35988),
            .I(data_count_6));
    Odrv4 I__7783 (
            .O(N__35985),
            .I(data_count_6));
    InMux I__7782 (
            .O(N__35978),
            .I(n13947));
    CascadeMux I__7781 (
            .O(N__35975),
            .I(N__35972));
    CascadeBuf I__7780 (
            .O(N__35972),
            .I(N__35969));
    CascadeMux I__7779 (
            .O(N__35969),
            .I(N__35966));
    CascadeBuf I__7778 (
            .O(N__35966),
            .I(N__35963));
    CascadeMux I__7777 (
            .O(N__35963),
            .I(N__35960));
    CascadeBuf I__7776 (
            .O(N__35960),
            .I(N__35957));
    CascadeMux I__7775 (
            .O(N__35957),
            .I(N__35954));
    CascadeBuf I__7774 (
            .O(N__35954),
            .I(N__35951));
    CascadeMux I__7773 (
            .O(N__35951),
            .I(N__35948));
    CascadeBuf I__7772 (
            .O(N__35948),
            .I(N__35945));
    CascadeMux I__7771 (
            .O(N__35945),
            .I(N__35942));
    CascadeBuf I__7770 (
            .O(N__35942),
            .I(N__35939));
    CascadeMux I__7769 (
            .O(N__35939),
            .I(N__35936));
    CascadeBuf I__7768 (
            .O(N__35936),
            .I(N__35933));
    CascadeMux I__7767 (
            .O(N__35933),
            .I(N__35930));
    CascadeBuf I__7766 (
            .O(N__35930),
            .I(N__35926));
    CascadeMux I__7765 (
            .O(N__35929),
            .I(N__35923));
    CascadeMux I__7764 (
            .O(N__35926),
            .I(N__35920));
    CascadeBuf I__7763 (
            .O(N__35923),
            .I(N__35917));
    CascadeBuf I__7762 (
            .O(N__35920),
            .I(N__35914));
    CascadeMux I__7761 (
            .O(N__35917),
            .I(N__35911));
    CascadeMux I__7760 (
            .O(N__35914),
            .I(N__35908));
    InMux I__7759 (
            .O(N__35911),
            .I(N__35905));
    InMux I__7758 (
            .O(N__35908),
            .I(N__35902));
    LocalMux I__7757 (
            .O(N__35905),
            .I(N__35899));
    LocalMux I__7756 (
            .O(N__35902),
            .I(N__35896));
    Span12Mux_v I__7755 (
            .O(N__35899),
            .I(N__35892));
    Span4Mux_h I__7754 (
            .O(N__35896),
            .I(N__35889));
    InMux I__7753 (
            .O(N__35895),
            .I(N__35886));
    Span12Mux_h I__7752 (
            .O(N__35892),
            .I(N__35883));
    Span4Mux_h I__7751 (
            .O(N__35889),
            .I(N__35880));
    LocalMux I__7750 (
            .O(N__35886),
            .I(data_count_7));
    Odrv12 I__7749 (
            .O(N__35883),
            .I(data_count_7));
    Odrv4 I__7748 (
            .O(N__35880),
            .I(data_count_7));
    InMux I__7747 (
            .O(N__35873),
            .I(n13948));
    InMux I__7746 (
            .O(N__35870),
            .I(bfn_16_19_0_));
    CascadeMux I__7745 (
            .O(N__35867),
            .I(N__35864));
    CascadeBuf I__7744 (
            .O(N__35864),
            .I(N__35861));
    CascadeMux I__7743 (
            .O(N__35861),
            .I(N__35858));
    CascadeBuf I__7742 (
            .O(N__35858),
            .I(N__35855));
    CascadeMux I__7741 (
            .O(N__35855),
            .I(N__35852));
    CascadeBuf I__7740 (
            .O(N__35852),
            .I(N__35849));
    CascadeMux I__7739 (
            .O(N__35849),
            .I(N__35846));
    CascadeBuf I__7738 (
            .O(N__35846),
            .I(N__35843));
    CascadeMux I__7737 (
            .O(N__35843),
            .I(N__35840));
    CascadeBuf I__7736 (
            .O(N__35840),
            .I(N__35837));
    CascadeMux I__7735 (
            .O(N__35837),
            .I(N__35834));
    CascadeBuf I__7734 (
            .O(N__35834),
            .I(N__35831));
    CascadeMux I__7733 (
            .O(N__35831),
            .I(N__35828));
    CascadeBuf I__7732 (
            .O(N__35828),
            .I(N__35825));
    CascadeMux I__7731 (
            .O(N__35825),
            .I(N__35822));
    CascadeBuf I__7730 (
            .O(N__35822),
            .I(N__35818));
    CascadeMux I__7729 (
            .O(N__35821),
            .I(N__35815));
    CascadeMux I__7728 (
            .O(N__35818),
            .I(N__35812));
    CascadeBuf I__7727 (
            .O(N__35815),
            .I(N__35809));
    CascadeBuf I__7726 (
            .O(N__35812),
            .I(N__35806));
    CascadeMux I__7725 (
            .O(N__35809),
            .I(N__35803));
    CascadeMux I__7724 (
            .O(N__35806),
            .I(N__35800));
    InMux I__7723 (
            .O(N__35803),
            .I(N__35797));
    InMux I__7722 (
            .O(N__35800),
            .I(N__35794));
    LocalMux I__7721 (
            .O(N__35797),
            .I(N__35791));
    LocalMux I__7720 (
            .O(N__35794),
            .I(N__35788));
    Span12Mux_v I__7719 (
            .O(N__35791),
            .I(N__35784));
    Span4Mux_h I__7718 (
            .O(N__35788),
            .I(N__35781));
    InMux I__7717 (
            .O(N__35787),
            .I(N__35778));
    Span12Mux_h I__7716 (
            .O(N__35784),
            .I(N__35775));
    Span4Mux_h I__7715 (
            .O(N__35781),
            .I(N__35772));
    LocalMux I__7714 (
            .O(N__35778),
            .I(data_count_8));
    Odrv12 I__7713 (
            .O(N__35775),
            .I(data_count_8));
    Odrv4 I__7712 (
            .O(N__35772),
            .I(data_count_8));
    InMux I__7711 (
            .O(N__35765),
            .I(N__35760));
    CascadeMux I__7710 (
            .O(N__35764),
            .I(N__35756));
    CascadeMux I__7709 (
            .O(N__35763),
            .I(N__35749));
    LocalMux I__7708 (
            .O(N__35760),
            .I(N__35743));
    CascadeMux I__7707 (
            .O(N__35759),
            .I(N__35738));
    InMux I__7706 (
            .O(N__35756),
            .I(N__35711));
    InMux I__7705 (
            .O(N__35755),
            .I(N__35711));
    InMux I__7704 (
            .O(N__35754),
            .I(N__35711));
    InMux I__7703 (
            .O(N__35753),
            .I(N__35711));
    InMux I__7702 (
            .O(N__35752),
            .I(N__35711));
    InMux I__7701 (
            .O(N__35749),
            .I(N__35711));
    InMux I__7700 (
            .O(N__35748),
            .I(N__35711));
    InMux I__7699 (
            .O(N__35747),
            .I(N__35711));
    InMux I__7698 (
            .O(N__35746),
            .I(N__35708));
    Span4Mux_h I__7697 (
            .O(N__35743),
            .I(N__35705));
    InMux I__7696 (
            .O(N__35742),
            .I(N__35688));
    InMux I__7695 (
            .O(N__35741),
            .I(N__35688));
    InMux I__7694 (
            .O(N__35738),
            .I(N__35688));
    InMux I__7693 (
            .O(N__35737),
            .I(N__35688));
    InMux I__7692 (
            .O(N__35736),
            .I(N__35688));
    InMux I__7691 (
            .O(N__35735),
            .I(N__35688));
    InMux I__7690 (
            .O(N__35734),
            .I(N__35688));
    InMux I__7689 (
            .O(N__35733),
            .I(N__35688));
    InMux I__7688 (
            .O(N__35732),
            .I(N__35677));
    InMux I__7687 (
            .O(N__35731),
            .I(N__35677));
    InMux I__7686 (
            .O(N__35730),
            .I(N__35677));
    InMux I__7685 (
            .O(N__35729),
            .I(N__35677));
    InMux I__7684 (
            .O(N__35728),
            .I(N__35677));
    LocalMux I__7683 (
            .O(N__35711),
            .I(N__35674));
    LocalMux I__7682 (
            .O(N__35708),
            .I(N__35671));
    Span4Mux_h I__7681 (
            .O(N__35705),
            .I(N__35662));
    LocalMux I__7680 (
            .O(N__35688),
            .I(N__35662));
    LocalMux I__7679 (
            .O(N__35677),
            .I(N__35662));
    Span12Mux_v I__7678 (
            .O(N__35674),
            .I(N__35659));
    Span4Mux_h I__7677 (
            .O(N__35671),
            .I(N__35656));
    InMux I__7676 (
            .O(N__35670),
            .I(N__35653));
    InMux I__7675 (
            .O(N__35669),
            .I(N__35650));
    Sp12to4 I__7674 (
            .O(N__35662),
            .I(N__35647));
    Odrv12 I__7673 (
            .O(N__35659),
            .I(dds_state_2));
    Odrv4 I__7672 (
            .O(N__35656),
            .I(dds_state_2));
    LocalMux I__7671 (
            .O(N__35653),
            .I(dds_state_2));
    LocalMux I__7670 (
            .O(N__35650),
            .I(dds_state_2));
    Odrv12 I__7669 (
            .O(N__35647),
            .I(dds_state_2));
    InMux I__7668 (
            .O(N__35636),
            .I(N__35633));
    LocalMux I__7667 (
            .O(N__35633),
            .I(N__35630));
    Span4Mux_h I__7666 (
            .O(N__35630),
            .I(N__35627));
    Span4Mux_v I__7665 (
            .O(N__35627),
            .I(N__35624));
    Span4Mux_v I__7664 (
            .O(N__35624),
            .I(N__35621));
    Odrv4 I__7663 (
            .O(N__35621),
            .I(\ADC_VAC2.n15280 ));
    InMux I__7662 (
            .O(N__35618),
            .I(N__35613));
    InMux I__7661 (
            .O(N__35617),
            .I(N__35610));
    InMux I__7660 (
            .O(N__35616),
            .I(N__35605));
    LocalMux I__7659 (
            .O(N__35613),
            .I(N__35600));
    LocalMux I__7658 (
            .O(N__35610),
            .I(N__35600));
    InMux I__7657 (
            .O(N__35609),
            .I(N__35592));
    InMux I__7656 (
            .O(N__35608),
            .I(N__35589));
    LocalMux I__7655 (
            .O(N__35605),
            .I(N__35586));
    Span4Mux_h I__7654 (
            .O(N__35600),
            .I(N__35583));
    InMux I__7653 (
            .O(N__35599),
            .I(N__35572));
    InMux I__7652 (
            .O(N__35598),
            .I(N__35572));
    InMux I__7651 (
            .O(N__35597),
            .I(N__35572));
    InMux I__7650 (
            .O(N__35596),
            .I(N__35572));
    InMux I__7649 (
            .O(N__35595),
            .I(N__35572));
    LocalMux I__7648 (
            .O(N__35592),
            .I(N__35569));
    LocalMux I__7647 (
            .O(N__35589),
            .I(N__35565));
    Span4Mux_h I__7646 (
            .O(N__35586),
            .I(N__35562));
    Span4Mux_h I__7645 (
            .O(N__35583),
            .I(N__35557));
    LocalMux I__7644 (
            .O(N__35572),
            .I(N__35557));
    Span4Mux_v I__7643 (
            .O(N__35569),
            .I(N__35554));
    InMux I__7642 (
            .O(N__35568),
            .I(N__35551));
    Span12Mux_s8_h I__7641 (
            .O(N__35565),
            .I(N__35546));
    Sp12to4 I__7640 (
            .O(N__35562),
            .I(N__35546));
    Span4Mux_h I__7639 (
            .O(N__35557),
            .I(N__35543));
    Sp12to4 I__7638 (
            .O(N__35554),
            .I(N__35540));
    LocalMux I__7637 (
            .O(N__35551),
            .I(N__35536));
    Span12Mux_v I__7636 (
            .O(N__35546),
            .I(N__35533));
    Span4Mux_h I__7635 (
            .O(N__35543),
            .I(N__35530));
    Span12Mux_h I__7634 (
            .O(N__35540),
            .I(N__35527));
    InMux I__7633 (
            .O(N__35539),
            .I(N__35524));
    Span12Mux_h I__7632 (
            .O(N__35536),
            .I(N__35517));
    Span12Mux_h I__7631 (
            .O(N__35533),
            .I(N__35517));
    Sp12to4 I__7630 (
            .O(N__35530),
            .I(N__35517));
    Odrv12 I__7629 (
            .O(N__35527),
            .I(adc_state_1_adj_1043));
    LocalMux I__7628 (
            .O(N__35524),
            .I(adc_state_1_adj_1043));
    Odrv12 I__7627 (
            .O(N__35517),
            .I(adc_state_1_adj_1043));
    CEMux I__7626 (
            .O(N__35510),
            .I(N__35507));
    LocalMux I__7625 (
            .O(N__35507),
            .I(N__35504));
    Span4Mux_h I__7624 (
            .O(N__35504),
            .I(N__35500));
    CEMux I__7623 (
            .O(N__35503),
            .I(N__35497));
    Span4Mux_v I__7622 (
            .O(N__35500),
            .I(N__35494));
    LocalMux I__7621 (
            .O(N__35497),
            .I(N__35491));
    Span4Mux_v I__7620 (
            .O(N__35494),
            .I(N__35488));
    Span4Mux_h I__7619 (
            .O(N__35491),
            .I(N__35485));
    Span4Mux_h I__7618 (
            .O(N__35488),
            .I(N__35480));
    Span4Mux_h I__7617 (
            .O(N__35485),
            .I(N__35480));
    Odrv4 I__7616 (
            .O(N__35480),
            .I(\ADC_VAC2.n12 ));
    CascadeMux I__7615 (
            .O(N__35477),
            .I(N__35474));
    InMux I__7614 (
            .O(N__35474),
            .I(N__35471));
    LocalMux I__7613 (
            .O(N__35471),
            .I(N__35467));
    InMux I__7612 (
            .O(N__35470),
            .I(N__35464));
    Span4Mux_h I__7611 (
            .O(N__35467),
            .I(N__35461));
    LocalMux I__7610 (
            .O(N__35464),
            .I(data_cntvec_12));
    Odrv4 I__7609 (
            .O(N__35461),
            .I(data_cntvec_12));
    InMux I__7608 (
            .O(N__35456),
            .I(n13962));
    CascadeMux I__7607 (
            .O(N__35453),
            .I(N__35450));
    InMux I__7606 (
            .O(N__35450),
            .I(N__35447));
    LocalMux I__7605 (
            .O(N__35447),
            .I(N__35443));
    InMux I__7604 (
            .O(N__35446),
            .I(N__35440));
    Span4Mux_v I__7603 (
            .O(N__35443),
            .I(N__35437));
    LocalMux I__7602 (
            .O(N__35440),
            .I(data_cntvec_13));
    Odrv4 I__7601 (
            .O(N__35437),
            .I(data_cntvec_13));
    InMux I__7600 (
            .O(N__35432),
            .I(n13963));
    CascadeMux I__7599 (
            .O(N__35429),
            .I(N__35426));
    InMux I__7598 (
            .O(N__35426),
            .I(N__35423));
    LocalMux I__7597 (
            .O(N__35423),
            .I(N__35419));
    InMux I__7596 (
            .O(N__35422),
            .I(N__35416));
    Span4Mux_h I__7595 (
            .O(N__35419),
            .I(N__35413));
    LocalMux I__7594 (
            .O(N__35416),
            .I(data_cntvec_14));
    Odrv4 I__7593 (
            .O(N__35413),
            .I(data_cntvec_14));
    InMux I__7592 (
            .O(N__35408),
            .I(n13964));
    InMux I__7591 (
            .O(N__35405),
            .I(n13965));
    CascadeMux I__7590 (
            .O(N__35402),
            .I(N__35399));
    InMux I__7589 (
            .O(N__35399),
            .I(N__35396));
    LocalMux I__7588 (
            .O(N__35396),
            .I(N__35392));
    InMux I__7587 (
            .O(N__35395),
            .I(N__35389));
    Span4Mux_h I__7586 (
            .O(N__35392),
            .I(N__35386));
    LocalMux I__7585 (
            .O(N__35389),
            .I(N__35381));
    Span4Mux_v I__7584 (
            .O(N__35386),
            .I(N__35381));
    Odrv4 I__7583 (
            .O(N__35381),
            .I(data_cntvec_15));
    CascadeMux I__7582 (
            .O(N__35378),
            .I(N__35375));
    CascadeBuf I__7581 (
            .O(N__35375),
            .I(N__35372));
    CascadeMux I__7580 (
            .O(N__35372),
            .I(N__35369));
    CascadeBuf I__7579 (
            .O(N__35369),
            .I(N__35366));
    CascadeMux I__7578 (
            .O(N__35366),
            .I(N__35363));
    CascadeBuf I__7577 (
            .O(N__35363),
            .I(N__35360));
    CascadeMux I__7576 (
            .O(N__35360),
            .I(N__35357));
    CascadeBuf I__7575 (
            .O(N__35357),
            .I(N__35354));
    CascadeMux I__7574 (
            .O(N__35354),
            .I(N__35351));
    CascadeBuf I__7573 (
            .O(N__35351),
            .I(N__35348));
    CascadeMux I__7572 (
            .O(N__35348),
            .I(N__35345));
    CascadeBuf I__7571 (
            .O(N__35345),
            .I(N__35342));
    CascadeMux I__7570 (
            .O(N__35342),
            .I(N__35339));
    CascadeBuf I__7569 (
            .O(N__35339),
            .I(N__35336));
    CascadeMux I__7568 (
            .O(N__35336),
            .I(N__35333));
    CascadeBuf I__7567 (
            .O(N__35333),
            .I(N__35329));
    CascadeMux I__7566 (
            .O(N__35332),
            .I(N__35326));
    CascadeMux I__7565 (
            .O(N__35329),
            .I(N__35323));
    CascadeBuf I__7564 (
            .O(N__35326),
            .I(N__35320));
    CascadeBuf I__7563 (
            .O(N__35323),
            .I(N__35317));
    CascadeMux I__7562 (
            .O(N__35320),
            .I(N__35314));
    CascadeMux I__7561 (
            .O(N__35317),
            .I(N__35311));
    InMux I__7560 (
            .O(N__35314),
            .I(N__35308));
    InMux I__7559 (
            .O(N__35311),
            .I(N__35305));
    LocalMux I__7558 (
            .O(N__35308),
            .I(N__35302));
    LocalMux I__7557 (
            .O(N__35305),
            .I(N__35299));
    Span12Mux_v I__7556 (
            .O(N__35302),
            .I(N__35295));
    Span4Mux_h I__7555 (
            .O(N__35299),
            .I(N__35292));
    InMux I__7554 (
            .O(N__35298),
            .I(N__35289));
    Span12Mux_h I__7553 (
            .O(N__35295),
            .I(N__35286));
    Span4Mux_h I__7552 (
            .O(N__35292),
            .I(N__35283));
    LocalMux I__7551 (
            .O(N__35289),
            .I(data_count_0));
    Odrv12 I__7550 (
            .O(N__35286),
            .I(data_count_0));
    Odrv4 I__7549 (
            .O(N__35283),
            .I(data_count_0));
    InMux I__7548 (
            .O(N__35276),
            .I(bfn_16_18_0_));
    CascadeMux I__7547 (
            .O(N__35273),
            .I(N__35270));
    CascadeBuf I__7546 (
            .O(N__35270),
            .I(N__35267));
    CascadeMux I__7545 (
            .O(N__35267),
            .I(N__35264));
    CascadeBuf I__7544 (
            .O(N__35264),
            .I(N__35261));
    CascadeMux I__7543 (
            .O(N__35261),
            .I(N__35258));
    CascadeBuf I__7542 (
            .O(N__35258),
            .I(N__35255));
    CascadeMux I__7541 (
            .O(N__35255),
            .I(N__35252));
    CascadeBuf I__7540 (
            .O(N__35252),
            .I(N__35249));
    CascadeMux I__7539 (
            .O(N__35249),
            .I(N__35246));
    CascadeBuf I__7538 (
            .O(N__35246),
            .I(N__35243));
    CascadeMux I__7537 (
            .O(N__35243),
            .I(N__35240));
    CascadeBuf I__7536 (
            .O(N__35240),
            .I(N__35237));
    CascadeMux I__7535 (
            .O(N__35237),
            .I(N__35234));
    CascadeBuf I__7534 (
            .O(N__35234),
            .I(N__35231));
    CascadeMux I__7533 (
            .O(N__35231),
            .I(N__35228));
    CascadeBuf I__7532 (
            .O(N__35228),
            .I(N__35224));
    CascadeMux I__7531 (
            .O(N__35227),
            .I(N__35221));
    CascadeMux I__7530 (
            .O(N__35224),
            .I(N__35218));
    CascadeBuf I__7529 (
            .O(N__35221),
            .I(N__35215));
    CascadeBuf I__7528 (
            .O(N__35218),
            .I(N__35212));
    CascadeMux I__7527 (
            .O(N__35215),
            .I(N__35209));
    CascadeMux I__7526 (
            .O(N__35212),
            .I(N__35206));
    InMux I__7525 (
            .O(N__35209),
            .I(N__35203));
    InMux I__7524 (
            .O(N__35206),
            .I(N__35200));
    LocalMux I__7523 (
            .O(N__35203),
            .I(N__35197));
    LocalMux I__7522 (
            .O(N__35200),
            .I(N__35194));
    Span12Mux_v I__7521 (
            .O(N__35197),
            .I(N__35190));
    Span4Mux_h I__7520 (
            .O(N__35194),
            .I(N__35187));
    InMux I__7519 (
            .O(N__35193),
            .I(N__35184));
    Span12Mux_h I__7518 (
            .O(N__35190),
            .I(N__35181));
    Span4Mux_h I__7517 (
            .O(N__35187),
            .I(N__35178));
    LocalMux I__7516 (
            .O(N__35184),
            .I(data_count_1));
    Odrv12 I__7515 (
            .O(N__35181),
            .I(data_count_1));
    Odrv4 I__7514 (
            .O(N__35178),
            .I(data_count_1));
    InMux I__7513 (
            .O(N__35171),
            .I(n13942));
    CascadeMux I__7512 (
            .O(N__35168),
            .I(N__35165));
    CascadeBuf I__7511 (
            .O(N__35165),
            .I(N__35162));
    CascadeMux I__7510 (
            .O(N__35162),
            .I(N__35159));
    CascadeBuf I__7509 (
            .O(N__35159),
            .I(N__35156));
    CascadeMux I__7508 (
            .O(N__35156),
            .I(N__35153));
    CascadeBuf I__7507 (
            .O(N__35153),
            .I(N__35150));
    CascadeMux I__7506 (
            .O(N__35150),
            .I(N__35147));
    CascadeBuf I__7505 (
            .O(N__35147),
            .I(N__35144));
    CascadeMux I__7504 (
            .O(N__35144),
            .I(N__35141));
    CascadeBuf I__7503 (
            .O(N__35141),
            .I(N__35138));
    CascadeMux I__7502 (
            .O(N__35138),
            .I(N__35135));
    CascadeBuf I__7501 (
            .O(N__35135),
            .I(N__35132));
    CascadeMux I__7500 (
            .O(N__35132),
            .I(N__35129));
    CascadeBuf I__7499 (
            .O(N__35129),
            .I(N__35126));
    CascadeMux I__7498 (
            .O(N__35126),
            .I(N__35123));
    CascadeBuf I__7497 (
            .O(N__35123),
            .I(N__35119));
    CascadeMux I__7496 (
            .O(N__35122),
            .I(N__35116));
    CascadeMux I__7495 (
            .O(N__35119),
            .I(N__35113));
    CascadeBuf I__7494 (
            .O(N__35116),
            .I(N__35110));
    CascadeBuf I__7493 (
            .O(N__35113),
            .I(N__35107));
    CascadeMux I__7492 (
            .O(N__35110),
            .I(N__35104));
    CascadeMux I__7491 (
            .O(N__35107),
            .I(N__35101));
    InMux I__7490 (
            .O(N__35104),
            .I(N__35098));
    InMux I__7489 (
            .O(N__35101),
            .I(N__35095));
    LocalMux I__7488 (
            .O(N__35098),
            .I(N__35092));
    LocalMux I__7487 (
            .O(N__35095),
            .I(N__35089));
    Span12Mux_v I__7486 (
            .O(N__35092),
            .I(N__35085));
    Span4Mux_v I__7485 (
            .O(N__35089),
            .I(N__35082));
    InMux I__7484 (
            .O(N__35088),
            .I(N__35079));
    Span12Mux_h I__7483 (
            .O(N__35085),
            .I(N__35076));
    Span4Mux_h I__7482 (
            .O(N__35082),
            .I(N__35073));
    LocalMux I__7481 (
            .O(N__35079),
            .I(data_count_2));
    Odrv12 I__7480 (
            .O(N__35076),
            .I(data_count_2));
    Odrv4 I__7479 (
            .O(N__35073),
            .I(data_count_2));
    InMux I__7478 (
            .O(N__35066),
            .I(n13943));
    CascadeMux I__7477 (
            .O(N__35063),
            .I(N__35060));
    CascadeBuf I__7476 (
            .O(N__35060),
            .I(N__35057));
    CascadeMux I__7475 (
            .O(N__35057),
            .I(N__35054));
    CascadeBuf I__7474 (
            .O(N__35054),
            .I(N__35051));
    CascadeMux I__7473 (
            .O(N__35051),
            .I(N__35048));
    CascadeBuf I__7472 (
            .O(N__35048),
            .I(N__35045));
    CascadeMux I__7471 (
            .O(N__35045),
            .I(N__35042));
    CascadeBuf I__7470 (
            .O(N__35042),
            .I(N__35039));
    CascadeMux I__7469 (
            .O(N__35039),
            .I(N__35036));
    CascadeBuf I__7468 (
            .O(N__35036),
            .I(N__35033));
    CascadeMux I__7467 (
            .O(N__35033),
            .I(N__35030));
    CascadeBuf I__7466 (
            .O(N__35030),
            .I(N__35027));
    CascadeMux I__7465 (
            .O(N__35027),
            .I(N__35024));
    CascadeBuf I__7464 (
            .O(N__35024),
            .I(N__35021));
    CascadeMux I__7463 (
            .O(N__35021),
            .I(N__35017));
    CascadeMux I__7462 (
            .O(N__35020),
            .I(N__35014));
    CascadeBuf I__7461 (
            .O(N__35017),
            .I(N__35011));
    CascadeBuf I__7460 (
            .O(N__35014),
            .I(N__35008));
    CascadeMux I__7459 (
            .O(N__35011),
            .I(N__35005));
    CascadeMux I__7458 (
            .O(N__35008),
            .I(N__35002));
    CascadeBuf I__7457 (
            .O(N__35005),
            .I(N__34999));
    InMux I__7456 (
            .O(N__35002),
            .I(N__34996));
    CascadeMux I__7455 (
            .O(N__34999),
            .I(N__34993));
    LocalMux I__7454 (
            .O(N__34996),
            .I(N__34990));
    InMux I__7453 (
            .O(N__34993),
            .I(N__34987));
    Sp12to4 I__7452 (
            .O(N__34990),
            .I(N__34984));
    LocalMux I__7451 (
            .O(N__34987),
            .I(N__34981));
    Span12Mux_v I__7450 (
            .O(N__34984),
            .I(N__34977));
    Span4Mux_v I__7449 (
            .O(N__34981),
            .I(N__34974));
    InMux I__7448 (
            .O(N__34980),
            .I(N__34971));
    Span12Mux_h I__7447 (
            .O(N__34977),
            .I(N__34968));
    Span4Mux_h I__7446 (
            .O(N__34974),
            .I(N__34965));
    LocalMux I__7445 (
            .O(N__34971),
            .I(data_count_3));
    Odrv12 I__7444 (
            .O(N__34968),
            .I(data_count_3));
    Odrv4 I__7443 (
            .O(N__34965),
            .I(data_count_3));
    InMux I__7442 (
            .O(N__34958),
            .I(n13944));
    InMux I__7441 (
            .O(N__34955),
            .I(n13953));
    InMux I__7440 (
            .O(N__34952),
            .I(n13954));
    InMux I__7439 (
            .O(N__34949),
            .I(n13955));
    InMux I__7438 (
            .O(N__34946),
            .I(N__34941));
    InMux I__7437 (
            .O(N__34945),
            .I(N__34938));
    InMux I__7436 (
            .O(N__34944),
            .I(N__34935));
    LocalMux I__7435 (
            .O(N__34941),
            .I(data_cntvec_6));
    LocalMux I__7434 (
            .O(N__34938),
            .I(data_cntvec_6));
    LocalMux I__7433 (
            .O(N__34935),
            .I(data_cntvec_6));
    InMux I__7432 (
            .O(N__34928),
            .I(n13956));
    InMux I__7431 (
            .O(N__34925),
            .I(N__34922));
    LocalMux I__7430 (
            .O(N__34922),
            .I(N__34917));
    InMux I__7429 (
            .O(N__34921),
            .I(N__34914));
    InMux I__7428 (
            .O(N__34920),
            .I(N__34911));
    Span4Mux_h I__7427 (
            .O(N__34917),
            .I(N__34908));
    LocalMux I__7426 (
            .O(N__34914),
            .I(N__34905));
    LocalMux I__7425 (
            .O(N__34911),
            .I(N__34900));
    Span4Mux_v I__7424 (
            .O(N__34908),
            .I(N__34900));
    Span4Mux_v I__7423 (
            .O(N__34905),
            .I(N__34897));
    Odrv4 I__7422 (
            .O(N__34900),
            .I(data_cntvec_7));
    Odrv4 I__7421 (
            .O(N__34897),
            .I(data_cntvec_7));
    InMux I__7420 (
            .O(N__34892),
            .I(n13957));
    InMux I__7419 (
            .O(N__34889),
            .I(N__34885));
    InMux I__7418 (
            .O(N__34888),
            .I(N__34882));
    LocalMux I__7417 (
            .O(N__34885),
            .I(N__34878));
    LocalMux I__7416 (
            .O(N__34882),
            .I(N__34875));
    InMux I__7415 (
            .O(N__34881),
            .I(N__34872));
    Span4Mux_v I__7414 (
            .O(N__34878),
            .I(N__34869));
    Span4Mux_h I__7413 (
            .O(N__34875),
            .I(N__34866));
    LocalMux I__7412 (
            .O(N__34872),
            .I(data_cntvec_8));
    Odrv4 I__7411 (
            .O(N__34869),
            .I(data_cntvec_8));
    Odrv4 I__7410 (
            .O(N__34866),
            .I(data_cntvec_8));
    InMux I__7409 (
            .O(N__34859),
            .I(bfn_16_17_0_));
    InMux I__7408 (
            .O(N__34856),
            .I(N__34852));
    InMux I__7407 (
            .O(N__34855),
            .I(N__34849));
    LocalMux I__7406 (
            .O(N__34852),
            .I(N__34846));
    LocalMux I__7405 (
            .O(N__34849),
            .I(N__34842));
    Span4Mux_h I__7404 (
            .O(N__34846),
            .I(N__34839));
    InMux I__7403 (
            .O(N__34845),
            .I(N__34836));
    Span4Mux_h I__7402 (
            .O(N__34842),
            .I(N__34833));
    Span4Mux_v I__7401 (
            .O(N__34839),
            .I(N__34830));
    LocalMux I__7400 (
            .O(N__34836),
            .I(data_cntvec_9));
    Odrv4 I__7399 (
            .O(N__34833),
            .I(data_cntvec_9));
    Odrv4 I__7398 (
            .O(N__34830),
            .I(data_cntvec_9));
    InMux I__7397 (
            .O(N__34823),
            .I(n13959));
    InMux I__7396 (
            .O(N__34820),
            .I(N__34816));
    InMux I__7395 (
            .O(N__34819),
            .I(N__34813));
    LocalMux I__7394 (
            .O(N__34816),
            .I(N__34809));
    LocalMux I__7393 (
            .O(N__34813),
            .I(N__34806));
    InMux I__7392 (
            .O(N__34812),
            .I(N__34803));
    Span4Mux_h I__7391 (
            .O(N__34809),
            .I(N__34800));
    Span12Mux_v I__7390 (
            .O(N__34806),
            .I(N__34797));
    LocalMux I__7389 (
            .O(N__34803),
            .I(data_cntvec_10));
    Odrv4 I__7388 (
            .O(N__34800),
            .I(data_cntvec_10));
    Odrv12 I__7387 (
            .O(N__34797),
            .I(data_cntvec_10));
    InMux I__7386 (
            .O(N__34790),
            .I(n13960));
    InMux I__7385 (
            .O(N__34787),
            .I(N__34783));
    InMux I__7384 (
            .O(N__34786),
            .I(N__34779));
    LocalMux I__7383 (
            .O(N__34783),
            .I(N__34776));
    InMux I__7382 (
            .O(N__34782),
            .I(N__34773));
    LocalMux I__7381 (
            .O(N__34779),
            .I(N__34768));
    Span4Mux_h I__7380 (
            .O(N__34776),
            .I(N__34768));
    LocalMux I__7379 (
            .O(N__34773),
            .I(data_cntvec_11));
    Odrv4 I__7378 (
            .O(N__34768),
            .I(data_cntvec_11));
    InMux I__7377 (
            .O(N__34763),
            .I(n13961));
    InMux I__7376 (
            .O(N__34760),
            .I(N__34755));
    InMux I__7375 (
            .O(N__34759),
            .I(N__34752));
    InMux I__7374 (
            .O(N__34758),
            .I(N__34749));
    LocalMux I__7373 (
            .O(N__34755),
            .I(N__34746));
    LocalMux I__7372 (
            .O(N__34752),
            .I(acadc_skipCount_6));
    LocalMux I__7371 (
            .O(N__34749),
            .I(acadc_skipCount_6));
    Odrv4 I__7370 (
            .O(N__34746),
            .I(acadc_skipCount_6));
    InMux I__7369 (
            .O(N__34739),
            .I(N__34736));
    LocalMux I__7368 (
            .O(N__34736),
            .I(N__34733));
    Span4Mux_h I__7367 (
            .O(N__34733),
            .I(N__34730));
    Span4Mux_h I__7366 (
            .O(N__34730),
            .I(N__34727));
    Odrv4 I__7365 (
            .O(N__34727),
            .I(buf_data1_14));
    CascadeMux I__7364 (
            .O(N__34724),
            .I(n4191_cascade_));
    InMux I__7363 (
            .O(N__34721),
            .I(N__34718));
    LocalMux I__7362 (
            .O(N__34718),
            .I(n4215));
    CascadeMux I__7361 (
            .O(N__34715),
            .I(n4228_cascade_));
    InMux I__7360 (
            .O(N__34712),
            .I(N__34709));
    LocalMux I__7359 (
            .O(N__34709),
            .I(n4203));
    CascadeMux I__7358 (
            .O(N__34706),
            .I(n4248_cascade_));
    InMux I__7357 (
            .O(N__34703),
            .I(N__34700));
    LocalMux I__7356 (
            .O(N__34700),
            .I(N__34697));
    Odrv12 I__7355 (
            .O(N__34697),
            .I(n4258));
    InMux I__7354 (
            .O(N__34694),
            .I(bfn_16_16_0_));
    InMux I__7353 (
            .O(N__34691),
            .I(n13951));
    InMux I__7352 (
            .O(N__34688),
            .I(N__34685));
    LocalMux I__7351 (
            .O(N__34685),
            .I(N__34680));
    InMux I__7350 (
            .O(N__34684),
            .I(N__34677));
    InMux I__7349 (
            .O(N__34683),
            .I(N__34674));
    Span4Mux_h I__7348 (
            .O(N__34680),
            .I(N__34671));
    LocalMux I__7347 (
            .O(N__34677),
            .I(N__34668));
    LocalMux I__7346 (
            .O(N__34674),
            .I(data_cntvec_2));
    Odrv4 I__7345 (
            .O(N__34671),
            .I(data_cntvec_2));
    Odrv4 I__7344 (
            .O(N__34668),
            .I(data_cntvec_2));
    InMux I__7343 (
            .O(N__34661),
            .I(n13952));
    InMux I__7342 (
            .O(N__34658),
            .I(N__34654));
    CascadeMux I__7341 (
            .O(N__34657),
            .I(N__34650));
    LocalMux I__7340 (
            .O(N__34654),
            .I(N__34647));
    InMux I__7339 (
            .O(N__34653),
            .I(N__34644));
    InMux I__7338 (
            .O(N__34650),
            .I(N__34641));
    Odrv4 I__7337 (
            .O(N__34647),
            .I(req_data_cnt_4));
    LocalMux I__7336 (
            .O(N__34644),
            .I(req_data_cnt_4));
    LocalMux I__7335 (
            .O(N__34641),
            .I(req_data_cnt_4));
    InMux I__7334 (
            .O(N__34634),
            .I(N__34631));
    LocalMux I__7333 (
            .O(N__34631),
            .I(n18_adj_1217));
    InMux I__7332 (
            .O(N__34628),
            .I(N__34625));
    LocalMux I__7331 (
            .O(N__34625),
            .I(N__34621));
    CascadeMux I__7330 (
            .O(N__34624),
            .I(N__34618));
    Span4Mux_h I__7329 (
            .O(N__34621),
            .I(N__34614));
    InMux I__7328 (
            .O(N__34618),
            .I(N__34611));
    InMux I__7327 (
            .O(N__34617),
            .I(N__34608));
    Span4Mux_v I__7326 (
            .O(N__34614),
            .I(N__34605));
    LocalMux I__7325 (
            .O(N__34611),
            .I(N__34602));
    LocalMux I__7324 (
            .O(N__34608),
            .I(buf_dds_6));
    Odrv4 I__7323 (
            .O(N__34605),
            .I(buf_dds_6));
    Odrv12 I__7322 (
            .O(N__34602),
            .I(buf_dds_6));
    InMux I__7321 (
            .O(N__34595),
            .I(N__34587));
    InMux I__7320 (
            .O(N__34594),
            .I(N__34584));
    InMux I__7319 (
            .O(N__34593),
            .I(N__34581));
    InMux I__7318 (
            .O(N__34592),
            .I(N__34578));
    InMux I__7317 (
            .O(N__34591),
            .I(N__34575));
    InMux I__7316 (
            .O(N__34590),
            .I(N__34572));
    LocalMux I__7315 (
            .O(N__34587),
            .I(N__34567));
    LocalMux I__7314 (
            .O(N__34584),
            .I(N__34567));
    LocalMux I__7313 (
            .O(N__34581),
            .I(N__34564));
    LocalMux I__7312 (
            .O(N__34578),
            .I(N__34561));
    LocalMux I__7311 (
            .O(N__34575),
            .I(N__34551));
    LocalMux I__7310 (
            .O(N__34572),
            .I(N__34551));
    Span4Mux_h I__7309 (
            .O(N__34567),
            .I(N__34551));
    Span4Mux_h I__7308 (
            .O(N__34564),
            .I(N__34551));
    Span4Mux_v I__7307 (
            .O(N__34561),
            .I(N__34547));
    InMux I__7306 (
            .O(N__34560),
            .I(N__34544));
    Span4Mux_h I__7305 (
            .O(N__34551),
            .I(N__34541));
    InMux I__7304 (
            .O(N__34550),
            .I(N__34538));
    Span4Mux_h I__7303 (
            .O(N__34547),
            .I(N__34535));
    LocalMux I__7302 (
            .O(N__34544),
            .I(N__34532));
    Odrv4 I__7301 (
            .O(N__34541),
            .I(comm_buf_0_1));
    LocalMux I__7300 (
            .O(N__34538),
            .I(comm_buf_0_1));
    Odrv4 I__7299 (
            .O(N__34535),
            .I(comm_buf_0_1));
    Odrv12 I__7298 (
            .O(N__34532),
            .I(comm_buf_0_1));
    InMux I__7297 (
            .O(N__34523),
            .I(N__34520));
    LocalMux I__7296 (
            .O(N__34520),
            .I(N__34516));
    InMux I__7295 (
            .O(N__34519),
            .I(N__34513));
    Odrv4 I__7294 (
            .O(N__34516),
            .I(n7485));
    LocalMux I__7293 (
            .O(N__34513),
            .I(n7485));
    InMux I__7292 (
            .O(N__34508),
            .I(N__34503));
    InMux I__7291 (
            .O(N__34507),
            .I(N__34499));
    InMux I__7290 (
            .O(N__34506),
            .I(N__34496));
    LocalMux I__7289 (
            .O(N__34503),
            .I(N__34493));
    InMux I__7288 (
            .O(N__34502),
            .I(N__34490));
    LocalMux I__7287 (
            .O(N__34499),
            .I(N__34487));
    LocalMux I__7286 (
            .O(N__34496),
            .I(N__34480));
    Span4Mux_v I__7285 (
            .O(N__34493),
            .I(N__34480));
    LocalMux I__7284 (
            .O(N__34490),
            .I(N__34480));
    Odrv12 I__7283 (
            .O(N__34487),
            .I(eis_stop));
    Odrv4 I__7282 (
            .O(N__34480),
            .I(eis_stop));
    InMux I__7281 (
            .O(N__34475),
            .I(N__34471));
    CascadeMux I__7280 (
            .O(N__34474),
            .I(N__34467));
    LocalMux I__7279 (
            .O(N__34471),
            .I(N__34464));
    CascadeMux I__7278 (
            .O(N__34470),
            .I(N__34461));
    InMux I__7277 (
            .O(N__34467),
            .I(N__34458));
    Span4Mux_h I__7276 (
            .O(N__34464),
            .I(N__34455));
    InMux I__7275 (
            .O(N__34461),
            .I(N__34452));
    LocalMux I__7274 (
            .O(N__34458),
            .I(cmd_rdadctmp_23_adj_1053));
    Odrv4 I__7273 (
            .O(N__34455),
            .I(cmd_rdadctmp_23_adj_1053));
    LocalMux I__7272 (
            .O(N__34452),
            .I(cmd_rdadctmp_23_adj_1053));
    InMux I__7271 (
            .O(N__34445),
            .I(N__34442));
    LocalMux I__7270 (
            .O(N__34442),
            .I(N__34438));
    InMux I__7269 (
            .O(N__34441),
            .I(N__34435));
    Span4Mux_v I__7268 (
            .O(N__34438),
            .I(N__34432));
    LocalMux I__7267 (
            .O(N__34435),
            .I(N__34427));
    Sp12to4 I__7266 (
            .O(N__34432),
            .I(N__34427));
    Odrv12 I__7265 (
            .O(N__34427),
            .I(buf_adcdata2_15));
    InMux I__7264 (
            .O(N__34424),
            .I(N__34420));
    InMux I__7263 (
            .O(N__34423),
            .I(N__34416));
    LocalMux I__7262 (
            .O(N__34420),
            .I(N__34413));
    InMux I__7261 (
            .O(N__34419),
            .I(N__34410));
    LocalMux I__7260 (
            .O(N__34416),
            .I(N__34400));
    Span4Mux_v I__7259 (
            .O(N__34413),
            .I(N__34400));
    LocalMux I__7258 (
            .O(N__34410),
            .I(N__34400));
    InMux I__7257 (
            .O(N__34409),
            .I(N__34397));
    InMux I__7256 (
            .O(N__34408),
            .I(N__34393));
    InMux I__7255 (
            .O(N__34407),
            .I(N__34390));
    Span4Mux_v I__7254 (
            .O(N__34400),
            .I(N__34385));
    LocalMux I__7253 (
            .O(N__34397),
            .I(N__34385));
    InMux I__7252 (
            .O(N__34396),
            .I(N__34382));
    LocalMux I__7251 (
            .O(N__34393),
            .I(N__34377));
    LocalMux I__7250 (
            .O(N__34390),
            .I(N__34377));
    Span4Mux_v I__7249 (
            .O(N__34385),
            .I(N__34374));
    LocalMux I__7248 (
            .O(N__34382),
            .I(N__34370));
    Span4Mux_v I__7247 (
            .O(N__34377),
            .I(N__34365));
    Span4Mux_h I__7246 (
            .O(N__34374),
            .I(N__34365));
    InMux I__7245 (
            .O(N__34373),
            .I(N__34362));
    Span4Mux_h I__7244 (
            .O(N__34370),
            .I(N__34359));
    Odrv4 I__7243 (
            .O(N__34365),
            .I(comm_buf_0_2));
    LocalMux I__7242 (
            .O(N__34362),
            .I(comm_buf_0_2));
    Odrv4 I__7241 (
            .O(N__34359),
            .I(comm_buf_0_2));
    InMux I__7240 (
            .O(N__34352),
            .I(N__34349));
    LocalMux I__7239 (
            .O(N__34349),
            .I(N__34345));
    InMux I__7238 (
            .O(N__34348),
            .I(N__34342));
    Span4Mux_v I__7237 (
            .O(N__34345),
            .I(N__34338));
    LocalMux I__7236 (
            .O(N__34342),
            .I(N__34335));
    InMux I__7235 (
            .O(N__34341),
            .I(N__34332));
    Span4Mux_v I__7234 (
            .O(N__34338),
            .I(N__34327));
    Span4Mux_v I__7233 (
            .O(N__34335),
            .I(N__34327));
    LocalMux I__7232 (
            .O(N__34332),
            .I(buf_dds_10));
    Odrv4 I__7231 (
            .O(N__34327),
            .I(buf_dds_10));
    InMux I__7230 (
            .O(N__34322),
            .I(N__34319));
    LocalMux I__7229 (
            .O(N__34319),
            .I(N__34315));
    InMux I__7228 (
            .O(N__34318),
            .I(N__34311));
    Span4Mux_h I__7227 (
            .O(N__34315),
            .I(N__34308));
    InMux I__7226 (
            .O(N__34314),
            .I(N__34305));
    LocalMux I__7225 (
            .O(N__34311),
            .I(acadc_skipCount_0));
    Odrv4 I__7224 (
            .O(N__34308),
            .I(acadc_skipCount_0));
    LocalMux I__7223 (
            .O(N__34305),
            .I(acadc_skipCount_0));
    InMux I__7222 (
            .O(N__34298),
            .I(N__34295));
    LocalMux I__7221 (
            .O(N__34295),
            .I(n17_adj_1214));
    CascadeMux I__7220 (
            .O(N__34292),
            .I(N__34289));
    InMux I__7219 (
            .O(N__34289),
            .I(N__34286));
    LocalMux I__7218 (
            .O(N__34286),
            .I(N__34281));
    InMux I__7217 (
            .O(N__34285),
            .I(N__34278));
    InMux I__7216 (
            .O(N__34284),
            .I(N__34275));
    Odrv4 I__7215 (
            .O(N__34281),
            .I(req_data_cnt_0));
    LocalMux I__7214 (
            .O(N__34278),
            .I(req_data_cnt_0));
    LocalMux I__7213 (
            .O(N__34275),
            .I(req_data_cnt_0));
    CascadeMux I__7212 (
            .O(N__34268),
            .I(N__34265));
    InMux I__7211 (
            .O(N__34265),
            .I(N__34262));
    LocalMux I__7210 (
            .O(N__34262),
            .I(N__34259));
    Span12Mux_v I__7209 (
            .O(N__34259),
            .I(N__34256));
    Odrv12 I__7208 (
            .O(N__34256),
            .I(buf_data1_21));
    InMux I__7207 (
            .O(N__34253),
            .I(N__34250));
    LocalMux I__7206 (
            .O(N__34250),
            .I(N__34247));
    Span4Mux_v I__7205 (
            .O(N__34247),
            .I(N__34244));
    Span4Mux_h I__7204 (
            .O(N__34244),
            .I(N__34241));
    Odrv4 I__7203 (
            .O(N__34241),
            .I(n66_adj_1158));
    CascadeMux I__7202 (
            .O(N__34238),
            .I(N__34235));
    InMux I__7201 (
            .O(N__34235),
            .I(N__34230));
    InMux I__7200 (
            .O(N__34234),
            .I(N__34227));
    InMux I__7199 (
            .O(N__34233),
            .I(N__34224));
    LocalMux I__7198 (
            .O(N__34230),
            .I(N__34221));
    LocalMux I__7197 (
            .O(N__34227),
            .I(buf_dds_5));
    LocalMux I__7196 (
            .O(N__34224),
            .I(buf_dds_5));
    Odrv12 I__7195 (
            .O(N__34221),
            .I(buf_dds_5));
    InMux I__7194 (
            .O(N__34214),
            .I(N__34211));
    LocalMux I__7193 (
            .O(N__34211),
            .I(N__34207));
    InMux I__7192 (
            .O(N__34210),
            .I(N__34203));
    Span4Mux_h I__7191 (
            .O(N__34207),
            .I(N__34200));
    InMux I__7190 (
            .O(N__34206),
            .I(N__34197));
    LocalMux I__7189 (
            .O(N__34203),
            .I(acadc_skipCount_10));
    Odrv4 I__7188 (
            .O(N__34200),
            .I(acadc_skipCount_10));
    LocalMux I__7187 (
            .O(N__34197),
            .I(acadc_skipCount_10));
    CascadeMux I__7186 (
            .O(N__34190),
            .I(n7485_cascade_));
    InMux I__7185 (
            .O(N__34187),
            .I(N__34181));
    InMux I__7184 (
            .O(N__34186),
            .I(N__34181));
    LocalMux I__7183 (
            .O(N__34181),
            .I(tacadc_rst));
    InMux I__7182 (
            .O(N__34178),
            .I(N__34173));
    InMux I__7181 (
            .O(N__34177),
            .I(N__34168));
    InMux I__7180 (
            .O(N__34176),
            .I(N__34168));
    LocalMux I__7179 (
            .O(N__34173),
            .I(req_data_cnt_10));
    LocalMux I__7178 (
            .O(N__34168),
            .I(req_data_cnt_10));
    CascadeMux I__7177 (
            .O(N__34163),
            .I(N__34160));
    InMux I__7176 (
            .O(N__34160),
            .I(N__34157));
    LocalMux I__7175 (
            .O(N__34157),
            .I(n90_adj_1167));
    InMux I__7174 (
            .O(N__34154),
            .I(N__34151));
    LocalMux I__7173 (
            .O(N__34151),
            .I(N__34148));
    Span4Mux_h I__7172 (
            .O(N__34148),
            .I(N__34145));
    Odrv4 I__7171 (
            .O(N__34145),
            .I(n72_adj_1162));
    InMux I__7170 (
            .O(N__34142),
            .I(N__34138));
    CascadeMux I__7169 (
            .O(N__34141),
            .I(N__34135));
    LocalMux I__7168 (
            .O(N__34138),
            .I(N__34130));
    InMux I__7167 (
            .O(N__34135),
            .I(N__34125));
    InMux I__7166 (
            .O(N__34134),
            .I(N__34125));
    InMux I__7165 (
            .O(N__34133),
            .I(N__34121));
    Span4Mux_h I__7164 (
            .O(N__34130),
            .I(N__34113));
    LocalMux I__7163 (
            .O(N__34125),
            .I(N__34113));
    InMux I__7162 (
            .O(N__34124),
            .I(N__34110));
    LocalMux I__7161 (
            .O(N__34121),
            .I(N__34107));
    InMux I__7160 (
            .O(N__34120),
            .I(N__34102));
    InMux I__7159 (
            .O(N__34119),
            .I(N__34102));
    InMux I__7158 (
            .O(N__34118),
            .I(N__34099));
    Span4Mux_v I__7157 (
            .O(N__34113),
            .I(N__34094));
    LocalMux I__7156 (
            .O(N__34110),
            .I(N__34094));
    Span4Mux_v I__7155 (
            .O(N__34107),
            .I(N__34089));
    LocalMux I__7154 (
            .O(N__34102),
            .I(N__34089));
    LocalMux I__7153 (
            .O(N__34099),
            .I(N__34084));
    Span4Mux_h I__7152 (
            .O(N__34094),
            .I(N__34084));
    Span4Mux_h I__7151 (
            .O(N__34089),
            .I(N__34081));
    Span4Mux_v I__7150 (
            .O(N__34084),
            .I(N__34078));
    Span4Mux_v I__7149 (
            .O(N__34081),
            .I(N__34075));
    Odrv4 I__7148 (
            .O(N__34078),
            .I(comm_buf_0_0));
    Odrv4 I__7147 (
            .O(N__34075),
            .I(comm_buf_0_0));
    CascadeMux I__7146 (
            .O(N__34070),
            .I(n14_adj_1202_cascade_));
    InMux I__7145 (
            .O(N__34067),
            .I(N__34064));
    LocalMux I__7144 (
            .O(N__34064),
            .I(N__34061));
    Span4Mux_v I__7143 (
            .O(N__34061),
            .I(N__34056));
    InMux I__7142 (
            .O(N__34060),
            .I(N__34051));
    InMux I__7141 (
            .O(N__34059),
            .I(N__34051));
    Odrv4 I__7140 (
            .O(N__34056),
            .I(buf_dds_13));
    LocalMux I__7139 (
            .O(N__34051),
            .I(buf_dds_13));
    InMux I__7138 (
            .O(N__34046),
            .I(N__34043));
    LocalMux I__7137 (
            .O(N__34043),
            .I(N__34040));
    Odrv12 I__7136 (
            .O(N__34040),
            .I(n15690));
    InMux I__7135 (
            .O(N__34037),
            .I(N__34034));
    LocalMux I__7134 (
            .O(N__34034),
            .I(N__34031));
    Span4Mux_h I__7133 (
            .O(N__34031),
            .I(N__34026));
    InMux I__7132 (
            .O(N__34030),
            .I(N__34023));
    InMux I__7131 (
            .O(N__34029),
            .I(N__34020));
    Span4Mux_h I__7130 (
            .O(N__34026),
            .I(N__34015));
    LocalMux I__7129 (
            .O(N__34023),
            .I(N__34015));
    LocalMux I__7128 (
            .O(N__34020),
            .I(req_data_cnt_12));
    Odrv4 I__7127 (
            .O(N__34015),
            .I(req_data_cnt_12));
    InMux I__7126 (
            .O(N__34010),
            .I(N__34007));
    LocalMux I__7125 (
            .O(N__34007),
            .I(N__34004));
    Odrv4 I__7124 (
            .O(N__34004),
            .I(n13_adj_1026));
    InMux I__7123 (
            .O(N__34001),
            .I(N__33998));
    LocalMux I__7122 (
            .O(N__33998),
            .I(N__33995));
    Odrv12 I__7121 (
            .O(N__33995),
            .I(buf_data1_17));
    CascadeMux I__7120 (
            .O(N__33992),
            .I(n78_cascade_));
    InMux I__7119 (
            .O(N__33989),
            .I(N__33986));
    LocalMux I__7118 (
            .O(N__33986),
            .I(N__33983));
    Span4Mux_h I__7117 (
            .O(N__33983),
            .I(N__33980));
    Odrv4 I__7116 (
            .O(N__33980),
            .I(n99_adj_1024));
    InMux I__7115 (
            .O(N__33977),
            .I(N__33974));
    LocalMux I__7114 (
            .O(N__33974),
            .I(n4257));
    InMux I__7113 (
            .O(N__33971),
            .I(N__33966));
    InMux I__7112 (
            .O(N__33970),
            .I(N__33963));
    InMux I__7111 (
            .O(N__33969),
            .I(N__33958));
    LocalMux I__7110 (
            .O(N__33966),
            .I(N__33953));
    LocalMux I__7109 (
            .O(N__33963),
            .I(N__33953));
    InMux I__7108 (
            .O(N__33962),
            .I(N__33950));
    InMux I__7107 (
            .O(N__33961),
            .I(N__33947));
    LocalMux I__7106 (
            .O(N__33958),
            .I(N__33944));
    Span4Mux_v I__7105 (
            .O(N__33953),
            .I(N__33941));
    LocalMux I__7104 (
            .O(N__33950),
            .I(N__33938));
    LocalMux I__7103 (
            .O(N__33947),
            .I(N__33933));
    Span4Mux_h I__7102 (
            .O(N__33944),
            .I(N__33933));
    Span4Mux_h I__7101 (
            .O(N__33941),
            .I(N__33930));
    Span12Mux_h I__7100 (
            .O(N__33938),
            .I(N__33927));
    Sp12to4 I__7099 (
            .O(N__33933),
            .I(N__33924));
    Span4Mux_h I__7098 (
            .O(N__33930),
            .I(N__33921));
    Odrv12 I__7097 (
            .O(N__33927),
            .I(comm_buf_1_6));
    Odrv12 I__7096 (
            .O(N__33924),
            .I(comm_buf_1_6));
    Odrv4 I__7095 (
            .O(N__33921),
            .I(comm_buf_1_6));
    InMux I__7094 (
            .O(N__33914),
            .I(N__33911));
    LocalMux I__7093 (
            .O(N__33911),
            .I(n8133));
    CascadeMux I__7092 (
            .O(N__33908),
            .I(N__33904));
    CascadeMux I__7091 (
            .O(N__33907),
            .I(N__33900));
    InMux I__7090 (
            .O(N__33904),
            .I(N__33897));
    CascadeMux I__7089 (
            .O(N__33903),
            .I(N__33893));
    InMux I__7088 (
            .O(N__33900),
            .I(N__33890));
    LocalMux I__7087 (
            .O(N__33897),
            .I(N__33887));
    InMux I__7086 (
            .O(N__33896),
            .I(N__33882));
    InMux I__7085 (
            .O(N__33893),
            .I(N__33882));
    LocalMux I__7084 (
            .O(N__33890),
            .I(trig_dds));
    Odrv12 I__7083 (
            .O(N__33887),
            .I(trig_dds));
    LocalMux I__7082 (
            .O(N__33882),
            .I(trig_dds));
    CascadeMux I__7081 (
            .O(N__33875),
            .I(N__33872));
    InMux I__7080 (
            .O(N__33872),
            .I(N__33867));
    InMux I__7079 (
            .O(N__33871),
            .I(N__33864));
    InMux I__7078 (
            .O(N__33870),
            .I(N__33861));
    LocalMux I__7077 (
            .O(N__33867),
            .I(N__33856));
    LocalMux I__7076 (
            .O(N__33864),
            .I(N__33856));
    LocalMux I__7075 (
            .O(N__33861),
            .I(buf_dds_0));
    Odrv12 I__7074 (
            .O(N__33856),
            .I(buf_dds_0));
    InMux I__7073 (
            .O(N__33851),
            .I(N__33846));
    CascadeMux I__7072 (
            .O(N__33850),
            .I(N__33843));
    InMux I__7071 (
            .O(N__33849),
            .I(N__33840));
    LocalMux I__7070 (
            .O(N__33846),
            .I(N__33837));
    InMux I__7069 (
            .O(N__33843),
            .I(N__33834));
    LocalMux I__7068 (
            .O(N__33840),
            .I(N__33831));
    Span4Mux_h I__7067 (
            .O(N__33837),
            .I(N__33828));
    LocalMux I__7066 (
            .O(N__33834),
            .I(buf_dds_8));
    Odrv4 I__7065 (
            .O(N__33831),
            .I(buf_dds_8));
    Odrv4 I__7064 (
            .O(N__33828),
            .I(buf_dds_8));
    InMux I__7063 (
            .O(N__33821),
            .I(N__33818));
    LocalMux I__7062 (
            .O(N__33818),
            .I(N__33815));
    Span12Mux_v I__7061 (
            .O(N__33815),
            .I(N__33812));
    Odrv12 I__7060 (
            .O(N__33812),
            .I(buf_data1_15));
    CascadeMux I__7059 (
            .O(N__33809),
            .I(n4190_cascade_));
    InMux I__7058 (
            .O(N__33806),
            .I(N__33803));
    LocalMux I__7057 (
            .O(N__33803),
            .I(n4227));
    InMux I__7056 (
            .O(N__33800),
            .I(N__33797));
    LocalMux I__7055 (
            .O(N__33797),
            .I(n4262));
    CascadeMux I__7054 (
            .O(N__33794),
            .I(N__33790));
    InMux I__7053 (
            .O(N__33793),
            .I(N__33786));
    InMux I__7052 (
            .O(N__33790),
            .I(N__33782));
    InMux I__7051 (
            .O(N__33789),
            .I(N__33779));
    LocalMux I__7050 (
            .O(N__33786),
            .I(N__33776));
    InMux I__7049 (
            .O(N__33785),
            .I(N__33772));
    LocalMux I__7048 (
            .O(N__33782),
            .I(N__33765));
    LocalMux I__7047 (
            .O(N__33779),
            .I(N__33765));
    Span4Mux_v I__7046 (
            .O(N__33776),
            .I(N__33765));
    InMux I__7045 (
            .O(N__33775),
            .I(N__33762));
    LocalMux I__7044 (
            .O(N__33772),
            .I(N__33759));
    Span4Mux_v I__7043 (
            .O(N__33765),
            .I(N__33756));
    LocalMux I__7042 (
            .O(N__33762),
            .I(N__33753));
    Span4Mux_v I__7041 (
            .O(N__33759),
            .I(N__33749));
    Span4Mux_h I__7040 (
            .O(N__33756),
            .I(N__33744));
    Span4Mux_h I__7039 (
            .O(N__33753),
            .I(N__33744));
    InMux I__7038 (
            .O(N__33752),
            .I(N__33741));
    Span4Mux_v I__7037 (
            .O(N__33749),
            .I(N__33736));
    Span4Mux_h I__7036 (
            .O(N__33744),
            .I(N__33736));
    LocalMux I__7035 (
            .O(N__33741),
            .I(comm_buf_0_5));
    Odrv4 I__7034 (
            .O(N__33736),
            .I(comm_buf_0_5));
    CascadeMux I__7033 (
            .O(N__33731),
            .I(n13_cascade_));
    InMux I__7032 (
            .O(N__33728),
            .I(N__33725));
    LocalMux I__7031 (
            .O(N__33725),
            .I(n6_adj_1273));
    InMux I__7030 (
            .O(N__33722),
            .I(N__33719));
    LocalMux I__7029 (
            .O(N__33719),
            .I(n5_adj_1282));
    InMux I__7028 (
            .O(N__33716),
            .I(N__33712));
    InMux I__7027 (
            .O(N__33715),
            .I(N__33709));
    LocalMux I__7026 (
            .O(N__33712),
            .I(comm_length_0));
    LocalMux I__7025 (
            .O(N__33709),
            .I(comm_length_0));
    SRMux I__7024 (
            .O(N__33704),
            .I(N__33701));
    LocalMux I__7023 (
            .O(N__33701),
            .I(N__33697));
    SRMux I__7022 (
            .O(N__33700),
            .I(N__33694));
    Span4Mux_h I__7021 (
            .O(N__33697),
            .I(N__33689));
    LocalMux I__7020 (
            .O(N__33694),
            .I(N__33686));
    SRMux I__7019 (
            .O(N__33693),
            .I(N__33683));
    SRMux I__7018 (
            .O(N__33692),
            .I(N__33680));
    Span4Mux_h I__7017 (
            .O(N__33689),
            .I(N__33677));
    Span4Mux_v I__7016 (
            .O(N__33686),
            .I(N__33674));
    LocalMux I__7015 (
            .O(N__33683),
            .I(N__33669));
    LocalMux I__7014 (
            .O(N__33680),
            .I(N__33669));
    Span4Mux_h I__7013 (
            .O(N__33677),
            .I(N__33666));
    Span4Mux_h I__7012 (
            .O(N__33674),
            .I(N__33661));
    Span4Mux_v I__7011 (
            .O(N__33669),
            .I(N__33661));
    Odrv4 I__7010 (
            .O(N__33666),
            .I(n10566));
    Odrv4 I__7009 (
            .O(N__33661),
            .I(n10566));
    InMux I__7008 (
            .O(N__33656),
            .I(N__33653));
    LocalMux I__7007 (
            .O(N__33653),
            .I(n13));
    CascadeMux I__7006 (
            .O(N__33650),
            .I(N__33646));
    InMux I__7005 (
            .O(N__33649),
            .I(N__33641));
    InMux I__7004 (
            .O(N__33646),
            .I(N__33641));
    LocalMux I__7003 (
            .O(N__33641),
            .I(N__33638));
    Odrv4 I__7002 (
            .O(N__33638),
            .I(n12649));
    CascadeMux I__7001 (
            .O(N__33635),
            .I(n8525_cascade_));
    InMux I__7000 (
            .O(N__33632),
            .I(N__33629));
    LocalMux I__6999 (
            .O(N__33629),
            .I(N__33622));
    InMux I__6998 (
            .O(N__33628),
            .I(N__33617));
    InMux I__6997 (
            .O(N__33627),
            .I(N__33617));
    InMux I__6996 (
            .O(N__33626),
            .I(N__33614));
    InMux I__6995 (
            .O(N__33625),
            .I(N__33611));
    Span4Mux_v I__6994 (
            .O(N__33622),
            .I(N__33608));
    LocalMux I__6993 (
            .O(N__33617),
            .I(N__33603));
    LocalMux I__6992 (
            .O(N__33614),
            .I(N__33603));
    LocalMux I__6991 (
            .O(N__33611),
            .I(n4075));
    Odrv4 I__6990 (
            .O(N__33608),
            .I(n4075));
    Odrv12 I__6989 (
            .O(N__33603),
            .I(n4075));
    CascadeMux I__6988 (
            .O(N__33596),
            .I(n15460_cascade_));
    CascadeMux I__6987 (
            .O(N__33593),
            .I(n19_cascade_));
    InMux I__6986 (
            .O(N__33590),
            .I(N__33587));
    LocalMux I__6985 (
            .O(N__33587),
            .I(n15463));
    InMux I__6984 (
            .O(N__33584),
            .I(N__33581));
    LocalMux I__6983 (
            .O(N__33581),
            .I(N__33578));
    Span4Mux_v I__6982 (
            .O(N__33578),
            .I(N__33575));
    Span4Mux_h I__6981 (
            .O(N__33575),
            .I(N__33572));
    Odrv4 I__6980 (
            .O(N__33572),
            .I(n23));
    CascadeMux I__6979 (
            .O(N__33569),
            .I(n19_adj_1151_cascade_));
    InMux I__6978 (
            .O(N__33566),
            .I(N__33563));
    LocalMux I__6977 (
            .O(N__33563),
            .I(N__33560));
    Span4Mux_v I__6976 (
            .O(N__33560),
            .I(N__33556));
    CascadeMux I__6975 (
            .O(N__33559),
            .I(N__33552));
    Span4Mux_h I__6974 (
            .O(N__33556),
            .I(N__33548));
    InMux I__6973 (
            .O(N__33555),
            .I(N__33541));
    InMux I__6972 (
            .O(N__33552),
            .I(N__33541));
    InMux I__6971 (
            .O(N__33551),
            .I(N__33541));
    Odrv4 I__6970 (
            .O(N__33548),
            .I(comm_length_2));
    LocalMux I__6969 (
            .O(N__33541),
            .I(comm_length_2));
    InMux I__6968 (
            .O(N__33536),
            .I(N__33526));
    InMux I__6967 (
            .O(N__33535),
            .I(N__33526));
    InMux I__6966 (
            .O(N__33534),
            .I(N__33513));
    InMux I__6965 (
            .O(N__33533),
            .I(N__33513));
    InMux I__6964 (
            .O(N__33532),
            .I(N__33513));
    InMux I__6963 (
            .O(N__33531),
            .I(N__33510));
    LocalMux I__6962 (
            .O(N__33526),
            .I(N__33507));
    InMux I__6961 (
            .O(N__33525),
            .I(N__33502));
    InMux I__6960 (
            .O(N__33524),
            .I(N__33502));
    InMux I__6959 (
            .O(N__33523),
            .I(N__33495));
    InMux I__6958 (
            .O(N__33522),
            .I(N__33495));
    InMux I__6957 (
            .O(N__33521),
            .I(N__33495));
    InMux I__6956 (
            .O(N__33520),
            .I(N__33492));
    LocalMux I__6955 (
            .O(N__33513),
            .I(N__33480));
    LocalMux I__6954 (
            .O(N__33510),
            .I(N__33471));
    Span4Mux_h I__6953 (
            .O(N__33507),
            .I(N__33471));
    LocalMux I__6952 (
            .O(N__33502),
            .I(N__33471));
    LocalMux I__6951 (
            .O(N__33495),
            .I(N__33471));
    LocalMux I__6950 (
            .O(N__33492),
            .I(N__33468));
    InMux I__6949 (
            .O(N__33491),
            .I(N__33461));
    InMux I__6948 (
            .O(N__33490),
            .I(N__33461));
    InMux I__6947 (
            .O(N__33489),
            .I(N__33461));
    CascadeMux I__6946 (
            .O(N__33488),
            .I(N__33456));
    InMux I__6945 (
            .O(N__33487),
            .I(N__33453));
    InMux I__6944 (
            .O(N__33486),
            .I(N__33450));
    InMux I__6943 (
            .O(N__33485),
            .I(N__33441));
    InMux I__6942 (
            .O(N__33484),
            .I(N__33441));
    InMux I__6941 (
            .O(N__33483),
            .I(N__33441));
    Span4Mux_v I__6940 (
            .O(N__33480),
            .I(N__33436));
    Span4Mux_v I__6939 (
            .O(N__33471),
            .I(N__33436));
    Span4Mux_v I__6938 (
            .O(N__33468),
            .I(N__33431));
    LocalMux I__6937 (
            .O(N__33461),
            .I(N__33431));
    InMux I__6936 (
            .O(N__33460),
            .I(N__33424));
    InMux I__6935 (
            .O(N__33459),
            .I(N__33424));
    InMux I__6934 (
            .O(N__33456),
            .I(N__33424));
    LocalMux I__6933 (
            .O(N__33453),
            .I(N__33419));
    LocalMux I__6932 (
            .O(N__33450),
            .I(N__33419));
    CascadeMux I__6931 (
            .O(N__33449),
            .I(N__33416));
    InMux I__6930 (
            .O(N__33448),
            .I(N__33411));
    LocalMux I__6929 (
            .O(N__33441),
            .I(N__33408));
    Span4Mux_h I__6928 (
            .O(N__33436),
            .I(N__33405));
    Span4Mux_h I__6927 (
            .O(N__33431),
            .I(N__33400));
    LocalMux I__6926 (
            .O(N__33424),
            .I(N__33400));
    Span4Mux_h I__6925 (
            .O(N__33419),
            .I(N__33397));
    InMux I__6924 (
            .O(N__33416),
            .I(N__33394));
    InMux I__6923 (
            .O(N__33415),
            .I(N__33389));
    InMux I__6922 (
            .O(N__33414),
            .I(N__33389));
    LocalMux I__6921 (
            .O(N__33411),
            .I(comm_index_2));
    Odrv12 I__6920 (
            .O(N__33408),
            .I(comm_index_2));
    Odrv4 I__6919 (
            .O(N__33405),
            .I(comm_index_2));
    Odrv4 I__6918 (
            .O(N__33400),
            .I(comm_index_2));
    Odrv4 I__6917 (
            .O(N__33397),
            .I(comm_index_2));
    LocalMux I__6916 (
            .O(N__33394),
            .I(comm_index_2));
    LocalMux I__6915 (
            .O(N__33389),
            .I(comm_index_2));
    CascadeMux I__6914 (
            .O(N__33374),
            .I(N__33368));
    InMux I__6913 (
            .O(N__33373),
            .I(N__33363));
    InMux I__6912 (
            .O(N__33372),
            .I(N__33363));
    InMux I__6911 (
            .O(N__33371),
            .I(N__33358));
    InMux I__6910 (
            .O(N__33368),
            .I(N__33358));
    LocalMux I__6909 (
            .O(N__33363),
            .I(comm_length_3));
    LocalMux I__6908 (
            .O(N__33358),
            .I(comm_length_3));
    InMux I__6907 (
            .O(N__33353),
            .I(N__33343));
    InMux I__6906 (
            .O(N__33352),
            .I(N__33340));
    InMux I__6905 (
            .O(N__33351),
            .I(N__33337));
    InMux I__6904 (
            .O(N__33350),
            .I(N__33332));
    InMux I__6903 (
            .O(N__33349),
            .I(N__33332));
    InMux I__6902 (
            .O(N__33348),
            .I(N__33325));
    InMux I__6901 (
            .O(N__33347),
            .I(N__33322));
    InMux I__6900 (
            .O(N__33346),
            .I(N__33317));
    LocalMux I__6899 (
            .O(N__33343),
            .I(N__33312));
    LocalMux I__6898 (
            .O(N__33340),
            .I(N__33312));
    LocalMux I__6897 (
            .O(N__33337),
            .I(N__33307));
    LocalMux I__6896 (
            .O(N__33332),
            .I(N__33307));
    InMux I__6895 (
            .O(N__33331),
            .I(N__33302));
    InMux I__6894 (
            .O(N__33330),
            .I(N__33302));
    CascadeMux I__6893 (
            .O(N__33329),
            .I(N__33299));
    CascadeMux I__6892 (
            .O(N__33328),
            .I(N__33296));
    LocalMux I__6891 (
            .O(N__33325),
            .I(N__33291));
    LocalMux I__6890 (
            .O(N__33322),
            .I(N__33288));
    InMux I__6889 (
            .O(N__33321),
            .I(N__33285));
    InMux I__6888 (
            .O(N__33320),
            .I(N__33282));
    LocalMux I__6887 (
            .O(N__33317),
            .I(N__33279));
    Span4Mux_h I__6886 (
            .O(N__33312),
            .I(N__33272));
    Span4Mux_v I__6885 (
            .O(N__33307),
            .I(N__33272));
    LocalMux I__6884 (
            .O(N__33302),
            .I(N__33272));
    InMux I__6883 (
            .O(N__33299),
            .I(N__33269));
    InMux I__6882 (
            .O(N__33296),
            .I(N__33262));
    InMux I__6881 (
            .O(N__33295),
            .I(N__33262));
    InMux I__6880 (
            .O(N__33294),
            .I(N__33262));
    Span4Mux_v I__6879 (
            .O(N__33291),
            .I(N__33255));
    Span4Mux_v I__6878 (
            .O(N__33288),
            .I(N__33255));
    LocalMux I__6877 (
            .O(N__33285),
            .I(N__33255));
    LocalMux I__6876 (
            .O(N__33282),
            .I(N__33252));
    Span4Mux_v I__6875 (
            .O(N__33279),
            .I(N__33246));
    Span4Mux_h I__6874 (
            .O(N__33272),
            .I(N__33239));
    LocalMux I__6873 (
            .O(N__33269),
            .I(N__33239));
    LocalMux I__6872 (
            .O(N__33262),
            .I(N__33239));
    Span4Mux_h I__6871 (
            .O(N__33255),
            .I(N__33234));
    Span4Mux_v I__6870 (
            .O(N__33252),
            .I(N__33234));
    InMux I__6869 (
            .O(N__33251),
            .I(N__33229));
    InMux I__6868 (
            .O(N__33250),
            .I(N__33229));
    InMux I__6867 (
            .O(N__33249),
            .I(N__33226));
    Odrv4 I__6866 (
            .O(N__33246),
            .I(comm_index_3));
    Odrv4 I__6865 (
            .O(N__33239),
            .I(comm_index_3));
    Odrv4 I__6864 (
            .O(N__33234),
            .I(comm_index_3));
    LocalMux I__6863 (
            .O(N__33229),
            .I(comm_index_3));
    LocalMux I__6862 (
            .O(N__33226),
            .I(comm_index_3));
    CascadeMux I__6861 (
            .O(N__33215),
            .I(n6_adj_1281_cascade_));
    InMux I__6860 (
            .O(N__33212),
            .I(N__33202));
    InMux I__6859 (
            .O(N__33211),
            .I(N__33195));
    InMux I__6858 (
            .O(N__33210),
            .I(N__33195));
    InMux I__6857 (
            .O(N__33209),
            .I(N__33195));
    InMux I__6856 (
            .O(N__33208),
            .I(N__33188));
    InMux I__6855 (
            .O(N__33207),
            .I(N__33188));
    InMux I__6854 (
            .O(N__33206),
            .I(N__33188));
    InMux I__6853 (
            .O(N__33205),
            .I(N__33185));
    LocalMux I__6852 (
            .O(N__33202),
            .I(N__33163));
    LocalMux I__6851 (
            .O(N__33195),
            .I(N__33163));
    LocalMux I__6850 (
            .O(N__33188),
            .I(N__33160));
    LocalMux I__6849 (
            .O(N__33185),
            .I(N__33157));
    InMux I__6848 (
            .O(N__33184),
            .I(N__33146));
    InMux I__6847 (
            .O(N__33183),
            .I(N__33146));
    InMux I__6846 (
            .O(N__33182),
            .I(N__33146));
    InMux I__6845 (
            .O(N__33181),
            .I(N__33146));
    InMux I__6844 (
            .O(N__33180),
            .I(N__33146));
    InMux I__6843 (
            .O(N__33179),
            .I(N__33141));
    InMux I__6842 (
            .O(N__33178),
            .I(N__33141));
    InMux I__6841 (
            .O(N__33177),
            .I(N__33138));
    InMux I__6840 (
            .O(N__33176),
            .I(N__33133));
    InMux I__6839 (
            .O(N__33175),
            .I(N__33133));
    InMux I__6838 (
            .O(N__33174),
            .I(N__33121));
    InMux I__6837 (
            .O(N__33173),
            .I(N__33121));
    InMux I__6836 (
            .O(N__33172),
            .I(N__33121));
    InMux I__6835 (
            .O(N__33171),
            .I(N__33121));
    InMux I__6834 (
            .O(N__33170),
            .I(N__33118));
    CascadeMux I__6833 (
            .O(N__33169),
            .I(N__33113));
    CascadeMux I__6832 (
            .O(N__33168),
            .I(N__33107));
    Span4Mux_v I__6831 (
            .O(N__33163),
            .I(N__33091));
    Span4Mux_v I__6830 (
            .O(N__33160),
            .I(N__33091));
    Span4Mux_v I__6829 (
            .O(N__33157),
            .I(N__33086));
    LocalMux I__6828 (
            .O(N__33146),
            .I(N__33086));
    LocalMux I__6827 (
            .O(N__33141),
            .I(N__33080));
    LocalMux I__6826 (
            .O(N__33138),
            .I(N__33080));
    LocalMux I__6825 (
            .O(N__33133),
            .I(N__33077));
    InMux I__6824 (
            .O(N__33132),
            .I(N__33070));
    InMux I__6823 (
            .O(N__33131),
            .I(N__33070));
    InMux I__6822 (
            .O(N__33130),
            .I(N__33070));
    LocalMux I__6821 (
            .O(N__33121),
            .I(N__33065));
    LocalMux I__6820 (
            .O(N__33118),
            .I(N__33065));
    InMux I__6819 (
            .O(N__33117),
            .I(N__33062));
    InMux I__6818 (
            .O(N__33116),
            .I(N__33059));
    InMux I__6817 (
            .O(N__33113),
            .I(N__33052));
    InMux I__6816 (
            .O(N__33112),
            .I(N__33052));
    InMux I__6815 (
            .O(N__33111),
            .I(N__33052));
    InMux I__6814 (
            .O(N__33110),
            .I(N__33041));
    InMux I__6813 (
            .O(N__33107),
            .I(N__33041));
    InMux I__6812 (
            .O(N__33106),
            .I(N__33041));
    InMux I__6811 (
            .O(N__33105),
            .I(N__33041));
    InMux I__6810 (
            .O(N__33104),
            .I(N__33041));
    InMux I__6809 (
            .O(N__33103),
            .I(N__33038));
    InMux I__6808 (
            .O(N__33102),
            .I(N__33031));
    InMux I__6807 (
            .O(N__33101),
            .I(N__33031));
    InMux I__6806 (
            .O(N__33100),
            .I(N__33031));
    InMux I__6805 (
            .O(N__33099),
            .I(N__33028));
    InMux I__6804 (
            .O(N__33098),
            .I(N__33021));
    InMux I__6803 (
            .O(N__33097),
            .I(N__33021));
    InMux I__6802 (
            .O(N__33096),
            .I(N__33021));
    Span4Mux_h I__6801 (
            .O(N__33091),
            .I(N__33015));
    Span4Mux_h I__6800 (
            .O(N__33086),
            .I(N__33015));
    InMux I__6799 (
            .O(N__33085),
            .I(N__33012));
    Span4Mux_v I__6798 (
            .O(N__33080),
            .I(N__33007));
    Span4Mux_v I__6797 (
            .O(N__33077),
            .I(N__33007));
    LocalMux I__6796 (
            .O(N__33070),
            .I(N__33002));
    Span4Mux_v I__6795 (
            .O(N__33065),
            .I(N__33002));
    LocalMux I__6794 (
            .O(N__33062),
            .I(N__32997));
    LocalMux I__6793 (
            .O(N__33059),
            .I(N__32997));
    LocalMux I__6792 (
            .O(N__33052),
            .I(N__32994));
    LocalMux I__6791 (
            .O(N__33041),
            .I(N__32991));
    LocalMux I__6790 (
            .O(N__33038),
            .I(N__32982));
    LocalMux I__6789 (
            .O(N__33031),
            .I(N__32982));
    LocalMux I__6788 (
            .O(N__33028),
            .I(N__32982));
    LocalMux I__6787 (
            .O(N__33021),
            .I(N__32982));
    InMux I__6786 (
            .O(N__33020),
            .I(N__32979));
    Span4Mux_h I__6785 (
            .O(N__33015),
            .I(N__32976));
    LocalMux I__6784 (
            .O(N__33012),
            .I(N__32973));
    Span4Mux_h I__6783 (
            .O(N__33007),
            .I(N__32964));
    Span4Mux_h I__6782 (
            .O(N__33002),
            .I(N__32964));
    Span4Mux_v I__6781 (
            .O(N__32997),
            .I(N__32964));
    Span4Mux_v I__6780 (
            .O(N__32994),
            .I(N__32964));
    Span12Mux_h I__6779 (
            .O(N__32991),
            .I(N__32959));
    Span12Mux_v I__6778 (
            .O(N__32982),
            .I(N__32959));
    LocalMux I__6777 (
            .O(N__32979),
            .I(comm_index_1));
    Odrv4 I__6776 (
            .O(N__32976),
            .I(comm_index_1));
    Odrv4 I__6775 (
            .O(N__32973),
            .I(comm_index_1));
    Odrv4 I__6774 (
            .O(N__32964),
            .I(comm_index_1));
    Odrv12 I__6773 (
            .O(N__32959),
            .I(comm_index_1));
    InMux I__6772 (
            .O(N__32948),
            .I(N__32945));
    LocalMux I__6771 (
            .O(N__32945),
            .I(n2));
    CascadeMux I__6770 (
            .O(N__32942),
            .I(n15119_cascade_));
    InMux I__6769 (
            .O(N__32939),
            .I(N__32933));
    InMux I__6768 (
            .O(N__32938),
            .I(N__32933));
    LocalMux I__6767 (
            .O(N__32933),
            .I(comm_length_1));
    InMux I__6766 (
            .O(N__32930),
            .I(N__32927));
    LocalMux I__6765 (
            .O(N__32927),
            .I(N__32920));
    InMux I__6764 (
            .O(N__32926),
            .I(N__32917));
    InMux I__6763 (
            .O(N__32925),
            .I(N__32913));
    CascadeMux I__6762 (
            .O(N__32924),
            .I(N__32908));
    CascadeMux I__6761 (
            .O(N__32923),
            .I(N__32905));
    Span4Mux_v I__6760 (
            .O(N__32920),
            .I(N__32900));
    LocalMux I__6759 (
            .O(N__32917),
            .I(N__32900));
    CascadeMux I__6758 (
            .O(N__32916),
            .I(N__32896));
    LocalMux I__6757 (
            .O(N__32913),
            .I(N__32893));
    CascadeMux I__6756 (
            .O(N__32912),
            .I(N__32890));
    InMux I__6755 (
            .O(N__32911),
            .I(N__32882));
    InMux I__6754 (
            .O(N__32908),
            .I(N__32882));
    InMux I__6753 (
            .O(N__32905),
            .I(N__32882));
    Span4Mux_h I__6752 (
            .O(N__32900),
            .I(N__32879));
    InMux I__6751 (
            .O(N__32899),
            .I(N__32872));
    InMux I__6750 (
            .O(N__32896),
            .I(N__32872));
    Span4Mux_v I__6749 (
            .O(N__32893),
            .I(N__32869));
    InMux I__6748 (
            .O(N__32890),
            .I(N__32866));
    InMux I__6747 (
            .O(N__32889),
            .I(N__32863));
    LocalMux I__6746 (
            .O(N__32882),
            .I(N__32858));
    Span4Mux_v I__6745 (
            .O(N__32879),
            .I(N__32858));
    InMux I__6744 (
            .O(N__32878),
            .I(N__32853));
    InMux I__6743 (
            .O(N__32877),
            .I(N__32853));
    LocalMux I__6742 (
            .O(N__32872),
            .I(eis_state_0));
    Odrv4 I__6741 (
            .O(N__32869),
            .I(eis_state_0));
    LocalMux I__6740 (
            .O(N__32866),
            .I(eis_state_0));
    LocalMux I__6739 (
            .O(N__32863),
            .I(eis_state_0));
    Odrv4 I__6738 (
            .O(N__32858),
            .I(eis_state_0));
    LocalMux I__6737 (
            .O(N__32853),
            .I(eis_state_0));
    CascadeMux I__6736 (
            .O(N__32840),
            .I(N__32837));
    InMux I__6735 (
            .O(N__32837),
            .I(N__32826));
    InMux I__6734 (
            .O(N__32836),
            .I(N__32826));
    InMux I__6733 (
            .O(N__32835),
            .I(N__32826));
    InMux I__6732 (
            .O(N__32834),
            .I(N__32823));
    InMux I__6731 (
            .O(N__32833),
            .I(N__32820));
    LocalMux I__6730 (
            .O(N__32826),
            .I(N__32815));
    LocalMux I__6729 (
            .O(N__32823),
            .I(N__32815));
    LocalMux I__6728 (
            .O(N__32820),
            .I(N__32803));
    Span4Mux_v I__6727 (
            .O(N__32815),
            .I(N__32803));
    InMux I__6726 (
            .O(N__32814),
            .I(N__32798));
    InMux I__6725 (
            .O(N__32813),
            .I(N__32798));
    InMux I__6724 (
            .O(N__32812),
            .I(N__32795));
    InMux I__6723 (
            .O(N__32811),
            .I(N__32790));
    InMux I__6722 (
            .O(N__32810),
            .I(N__32790));
    InMux I__6721 (
            .O(N__32809),
            .I(N__32785));
    InMux I__6720 (
            .O(N__32808),
            .I(N__32785));
    Span4Mux_v I__6719 (
            .O(N__32803),
            .I(N__32782));
    LocalMux I__6718 (
            .O(N__32798),
            .I(eis_end_N_770));
    LocalMux I__6717 (
            .O(N__32795),
            .I(eis_end_N_770));
    LocalMux I__6716 (
            .O(N__32790),
            .I(eis_end_N_770));
    LocalMux I__6715 (
            .O(N__32785),
            .I(eis_end_N_770));
    Odrv4 I__6714 (
            .O(N__32782),
            .I(eis_end_N_770));
    InMux I__6713 (
            .O(N__32771),
            .I(N__32768));
    LocalMux I__6712 (
            .O(N__32768),
            .I(N__32764));
    CascadeMux I__6711 (
            .O(N__32767),
            .I(N__32760));
    Span4Mux_v I__6710 (
            .O(N__32764),
            .I(N__32757));
    CascadeMux I__6709 (
            .O(N__32763),
            .I(N__32754));
    InMux I__6708 (
            .O(N__32760),
            .I(N__32750));
    Span4Mux_h I__6707 (
            .O(N__32757),
            .I(N__32747));
    InMux I__6706 (
            .O(N__32754),
            .I(N__32744));
    SRMux I__6705 (
            .O(N__32753),
            .I(N__32741));
    LocalMux I__6704 (
            .O(N__32750),
            .I(N__32738));
    Span4Mux_h I__6703 (
            .O(N__32747),
            .I(N__32730));
    LocalMux I__6702 (
            .O(N__32744),
            .I(N__32730));
    LocalMux I__6701 (
            .O(N__32741),
            .I(N__32725));
    Span4Mux_h I__6700 (
            .O(N__32738),
            .I(N__32722));
    InMux I__6699 (
            .O(N__32737),
            .I(N__32715));
    InMux I__6698 (
            .O(N__32736),
            .I(N__32715));
    InMux I__6697 (
            .O(N__32735),
            .I(N__32715));
    Span4Mux_v I__6696 (
            .O(N__32730),
            .I(N__32712));
    InMux I__6695 (
            .O(N__32729),
            .I(N__32707));
    InMux I__6694 (
            .O(N__32728),
            .I(N__32707));
    Span4Mux_v I__6693 (
            .O(N__32725),
            .I(N__32704));
    Span4Mux_v I__6692 (
            .O(N__32722),
            .I(N__32699));
    LocalMux I__6691 (
            .O(N__32715),
            .I(N__32699));
    Sp12to4 I__6690 (
            .O(N__32712),
            .I(N__32696));
    LocalMux I__6689 (
            .O(N__32707),
            .I(N__32693));
    Span4Mux_v I__6688 (
            .O(N__32704),
            .I(N__32688));
    Span4Mux_v I__6687 (
            .O(N__32699),
            .I(N__32688));
    Span12Mux_h I__6686 (
            .O(N__32696),
            .I(N__32685));
    Span12Mux_v I__6685 (
            .O(N__32693),
            .I(N__32682));
    Sp12to4 I__6684 (
            .O(N__32688),
            .I(N__32679));
    Span12Mux_v I__6683 (
            .O(N__32685),
            .I(N__32676));
    Span12Mux_v I__6682 (
            .O(N__32682),
            .I(N__32673));
    Span12Mux_h I__6681 (
            .O(N__32679),
            .I(N__32670));
    Span12Mux_v I__6680 (
            .O(N__32676),
            .I(N__32667));
    Span12Mux_h I__6679 (
            .O(N__32673),
            .I(N__32662));
    Span12Mux_v I__6678 (
            .O(N__32670),
            .I(N__32662));
    Odrv12 I__6677 (
            .O(N__32667),
            .I(ICE_GPMO_0));
    Odrv12 I__6676 (
            .O(N__32662),
            .I(ICE_GPMO_0));
    InMux I__6675 (
            .O(N__32657),
            .I(N__32652));
    InMux I__6674 (
            .O(N__32656),
            .I(N__32647));
    InMux I__6673 (
            .O(N__32655),
            .I(N__32647));
    LocalMux I__6672 (
            .O(N__32652),
            .I(N__32644));
    LocalMux I__6671 (
            .O(N__32647),
            .I(N__32641));
    Span4Mux_h I__6670 (
            .O(N__32644),
            .I(N__32636));
    Span4Mux_h I__6669 (
            .O(N__32641),
            .I(N__32636));
    Odrv4 I__6668 (
            .O(N__32636),
            .I(data_index_8));
    InMux I__6667 (
            .O(N__32633),
            .I(N__32630));
    LocalMux I__6666 (
            .O(N__32630),
            .I(N__32627));
    Odrv12 I__6665 (
            .O(N__32627),
            .I(buf_data1_3));
    InMux I__6664 (
            .O(N__32624),
            .I(N__32620));
    InMux I__6663 (
            .O(N__32623),
            .I(N__32616));
    LocalMux I__6662 (
            .O(N__32620),
            .I(N__32613));
    CascadeMux I__6661 (
            .O(N__32619),
            .I(N__32610));
    LocalMux I__6660 (
            .O(N__32616),
            .I(N__32607));
    Span12Mux_v I__6659 (
            .O(N__32613),
            .I(N__32604));
    InMux I__6658 (
            .O(N__32610),
            .I(N__32601));
    Sp12to4 I__6657 (
            .O(N__32607),
            .I(N__32598));
    Span12Mux_h I__6656 (
            .O(N__32604),
            .I(N__32595));
    LocalMux I__6655 (
            .O(N__32601),
            .I(N__32590));
    Span12Mux_v I__6654 (
            .O(N__32598),
            .I(N__32590));
    Span12Mux_v I__6653 (
            .O(N__32595),
            .I(N__32587));
    Odrv12 I__6652 (
            .O(N__32590),
            .I(buf_adcdata3_3));
    Odrv12 I__6651 (
            .O(N__32587),
            .I(buf_adcdata3_3));
    InMux I__6650 (
            .O(N__32582),
            .I(N__32579));
    LocalMux I__6649 (
            .O(N__32579),
            .I(N__32576));
    Span4Mux_v I__6648 (
            .O(N__32576),
            .I(N__32573));
    Span4Mux_h I__6647 (
            .O(N__32573),
            .I(N__32570));
    Span4Mux_h I__6646 (
            .O(N__32570),
            .I(N__32567));
    Odrv4 I__6645 (
            .O(N__32567),
            .I(n4149));
    InMux I__6644 (
            .O(N__32564),
            .I(N__32559));
    InMux I__6643 (
            .O(N__32563),
            .I(N__32554));
    InMux I__6642 (
            .O(N__32562),
            .I(N__32554));
    LocalMux I__6641 (
            .O(N__32559),
            .I(N__32551));
    LocalMux I__6640 (
            .O(N__32554),
            .I(N__32548));
    Span4Mux_h I__6639 (
            .O(N__32551),
            .I(N__32543));
    Span4Mux_v I__6638 (
            .O(N__32548),
            .I(N__32543));
    Span4Mux_h I__6637 (
            .O(N__32543),
            .I(N__32540));
    Odrv4 I__6636 (
            .O(N__32540),
            .I(comm_tx_buf_5));
    SRMux I__6635 (
            .O(N__32537),
            .I(N__32534));
    LocalMux I__6634 (
            .O(N__32534),
            .I(N__32531));
    Span4Mux_v I__6633 (
            .O(N__32531),
            .I(N__32528));
    Sp12to4 I__6632 (
            .O(N__32528),
            .I(N__32525));
    Odrv12 I__6631 (
            .O(N__32525),
            .I(\comm_spi.data_tx_7__N_819 ));
    CEMux I__6630 (
            .O(N__32522),
            .I(N__32519));
    LocalMux I__6629 (
            .O(N__32519),
            .I(N__32515));
    CEMux I__6628 (
            .O(N__32518),
            .I(N__32512));
    Span4Mux_h I__6627 (
            .O(N__32515),
            .I(N__32509));
    LocalMux I__6626 (
            .O(N__32512),
            .I(N__32506));
    Odrv4 I__6625 (
            .O(N__32509),
            .I(n8561));
    Odrv4 I__6624 (
            .O(N__32506),
            .I(n8561));
    InMux I__6623 (
            .O(N__32501),
            .I(N__32497));
    InMux I__6622 (
            .O(N__32500),
            .I(N__32494));
    LocalMux I__6621 (
            .O(N__32497),
            .I(n8_adj_1229));
    LocalMux I__6620 (
            .O(N__32494),
            .I(n8_adj_1229));
    InMux I__6619 (
            .O(N__32489),
            .I(N__32485));
    InMux I__6618 (
            .O(N__32488),
            .I(N__32482));
    LocalMux I__6617 (
            .O(N__32485),
            .I(n7_adj_1228));
    LocalMux I__6616 (
            .O(N__32482),
            .I(n7_adj_1228));
    CascadeMux I__6615 (
            .O(N__32477),
            .I(N__32474));
    CascadeBuf I__6614 (
            .O(N__32474),
            .I(N__32471));
    CascadeMux I__6613 (
            .O(N__32471),
            .I(N__32468));
    CascadeBuf I__6612 (
            .O(N__32468),
            .I(N__32465));
    CascadeMux I__6611 (
            .O(N__32465),
            .I(N__32462));
    CascadeBuf I__6610 (
            .O(N__32462),
            .I(N__32459));
    CascadeMux I__6609 (
            .O(N__32459),
            .I(N__32456));
    CascadeBuf I__6608 (
            .O(N__32456),
            .I(N__32453));
    CascadeMux I__6607 (
            .O(N__32453),
            .I(N__32450));
    CascadeBuf I__6606 (
            .O(N__32450),
            .I(N__32447));
    CascadeMux I__6605 (
            .O(N__32447),
            .I(N__32444));
    CascadeBuf I__6604 (
            .O(N__32444),
            .I(N__32441));
    CascadeMux I__6603 (
            .O(N__32441),
            .I(N__32437));
    CascadeMux I__6602 (
            .O(N__32440),
            .I(N__32434));
    CascadeBuf I__6601 (
            .O(N__32437),
            .I(N__32431));
    CascadeBuf I__6600 (
            .O(N__32434),
            .I(N__32428));
    CascadeMux I__6599 (
            .O(N__32431),
            .I(N__32425));
    CascadeMux I__6598 (
            .O(N__32428),
            .I(N__32422));
    CascadeBuf I__6597 (
            .O(N__32425),
            .I(N__32419));
    InMux I__6596 (
            .O(N__32422),
            .I(N__32416));
    CascadeMux I__6595 (
            .O(N__32419),
            .I(N__32413));
    LocalMux I__6594 (
            .O(N__32416),
            .I(N__32410));
    CascadeBuf I__6593 (
            .O(N__32413),
            .I(N__32407));
    Span4Mux_h I__6592 (
            .O(N__32410),
            .I(N__32404));
    CascadeMux I__6591 (
            .O(N__32407),
            .I(N__32401));
    Span4Mux_v I__6590 (
            .O(N__32404),
            .I(N__32398));
    InMux I__6589 (
            .O(N__32401),
            .I(N__32395));
    Span4Mux_v I__6588 (
            .O(N__32398),
            .I(N__32392));
    LocalMux I__6587 (
            .O(N__32395),
            .I(N__32389));
    Span4Mux_h I__6586 (
            .O(N__32392),
            .I(N__32386));
    Span4Mux_h I__6585 (
            .O(N__32389),
            .I(N__32383));
    Span4Mux_h I__6584 (
            .O(N__32386),
            .I(N__32378));
    Span4Mux_h I__6583 (
            .O(N__32383),
            .I(N__32378));
    Odrv4 I__6582 (
            .O(N__32378),
            .I(data_index_9_N_258_3));
    CEMux I__6581 (
            .O(N__32375),
            .I(N__32372));
    LocalMux I__6580 (
            .O(N__32372),
            .I(N__32368));
    CEMux I__6579 (
            .O(N__32371),
            .I(N__32364));
    Span4Mux_h I__6578 (
            .O(N__32368),
            .I(N__32361));
    CEMux I__6577 (
            .O(N__32367),
            .I(N__32358));
    LocalMux I__6576 (
            .O(N__32364),
            .I(N__32355));
    Span4Mux_h I__6575 (
            .O(N__32361),
            .I(N__32352));
    LocalMux I__6574 (
            .O(N__32358),
            .I(N__32349));
    Span4Mux_h I__6573 (
            .O(N__32355),
            .I(N__32346));
    Span4Mux_h I__6572 (
            .O(N__32352),
            .I(N__32342));
    Span4Mux_h I__6571 (
            .O(N__32349),
            .I(N__32339));
    Span4Mux_h I__6570 (
            .O(N__32346),
            .I(N__32336));
    InMux I__6569 (
            .O(N__32345),
            .I(N__32333));
    Odrv4 I__6568 (
            .O(N__32342),
            .I(n8456));
    Odrv4 I__6567 (
            .O(N__32339),
            .I(n8456));
    Odrv4 I__6566 (
            .O(N__32336),
            .I(n8456));
    LocalMux I__6565 (
            .O(N__32333),
            .I(n8456));
    InMux I__6564 (
            .O(N__32324),
            .I(N__32320));
    InMux I__6563 (
            .O(N__32323),
            .I(N__32317));
    LocalMux I__6562 (
            .O(N__32320),
            .I(N__32312));
    LocalMux I__6561 (
            .O(N__32317),
            .I(N__32312));
    Odrv4 I__6560 (
            .O(N__32312),
            .I(acadc_skipcnt_3));
    CascadeMux I__6559 (
            .O(N__32309),
            .I(N__32306));
    InMux I__6558 (
            .O(N__32306),
            .I(N__32302));
    InMux I__6557 (
            .O(N__32305),
            .I(N__32299));
    LocalMux I__6556 (
            .O(N__32302),
            .I(N__32296));
    LocalMux I__6555 (
            .O(N__32299),
            .I(acadc_skipcnt_5));
    Odrv4 I__6554 (
            .O(N__32296),
            .I(acadc_skipcnt_5));
    InMux I__6553 (
            .O(N__32291),
            .I(N__32287));
    InMux I__6552 (
            .O(N__32290),
            .I(N__32284));
    LocalMux I__6551 (
            .O(N__32287),
            .I(N__32281));
    LocalMux I__6550 (
            .O(N__32284),
            .I(acadc_skipcnt_8));
    Odrv4 I__6549 (
            .O(N__32281),
            .I(acadc_skipcnt_8));
    InMux I__6548 (
            .O(N__32276),
            .I(N__32273));
    LocalMux I__6547 (
            .O(N__32273),
            .I(N__32268));
    InMux I__6546 (
            .O(N__32272),
            .I(N__32265));
    InMux I__6545 (
            .O(N__32271),
            .I(N__32262));
    Span4Mux_v I__6544 (
            .O(N__32268),
            .I(N__32259));
    LocalMux I__6543 (
            .O(N__32265),
            .I(N__32256));
    LocalMux I__6542 (
            .O(N__32262),
            .I(acadc_skipCount_8));
    Odrv4 I__6541 (
            .O(N__32259),
            .I(acadc_skipCount_8));
    Odrv4 I__6540 (
            .O(N__32256),
            .I(acadc_skipCount_8));
    CascadeMux I__6539 (
            .O(N__32249),
            .I(n20_cascade_));
    InMux I__6538 (
            .O(N__32246),
            .I(N__32243));
    LocalMux I__6537 (
            .O(N__32243),
            .I(N__32240));
    Span4Mux_h I__6536 (
            .O(N__32240),
            .I(N__32237));
    Odrv4 I__6535 (
            .O(N__32237),
            .I(n26));
    InMux I__6534 (
            .O(N__32234),
            .I(N__32231));
    LocalMux I__6533 (
            .O(N__32231),
            .I(N__32227));
    InMux I__6532 (
            .O(N__32230),
            .I(N__32224));
    Span4Mux_h I__6531 (
            .O(N__32227),
            .I(N__32221));
    LocalMux I__6530 (
            .O(N__32224),
            .I(acadc_skipcnt_13));
    Odrv4 I__6529 (
            .O(N__32221),
            .I(acadc_skipcnt_13));
    InMux I__6528 (
            .O(N__32216),
            .I(N__32212));
    CascadeMux I__6527 (
            .O(N__32215),
            .I(N__32209));
    LocalMux I__6526 (
            .O(N__32212),
            .I(N__32206));
    InMux I__6525 (
            .O(N__32209),
            .I(N__32202));
    Span12Mux_h I__6524 (
            .O(N__32206),
            .I(N__32199));
    InMux I__6523 (
            .O(N__32205),
            .I(N__32196));
    LocalMux I__6522 (
            .O(N__32202),
            .I(acadc_skipCount_13));
    Odrv12 I__6521 (
            .O(N__32199),
            .I(acadc_skipCount_13));
    LocalMux I__6520 (
            .O(N__32196),
            .I(acadc_skipCount_13));
    InMux I__6519 (
            .O(N__32189),
            .I(N__32186));
    LocalMux I__6518 (
            .O(N__32186),
            .I(n14_adj_1160));
    CascadeMux I__6517 (
            .O(N__32183),
            .I(N__32180));
    InMux I__6516 (
            .O(N__32180),
            .I(N__32177));
    LocalMux I__6515 (
            .O(N__32177),
            .I(N__32174));
    Span4Mux_v I__6514 (
            .O(N__32174),
            .I(N__32170));
    InMux I__6513 (
            .O(N__32173),
            .I(N__32167));
    Span4Mux_h I__6512 (
            .O(N__32170),
            .I(N__32161));
    LocalMux I__6511 (
            .O(N__32167),
            .I(N__32161));
    CascadeMux I__6510 (
            .O(N__32166),
            .I(N__32158));
    Span4Mux_h I__6509 (
            .O(N__32161),
            .I(N__32155));
    InMux I__6508 (
            .O(N__32158),
            .I(N__32152));
    Odrv4 I__6507 (
            .O(N__32155),
            .I(cmd_rdadctmp_16));
    LocalMux I__6506 (
            .O(N__32152),
            .I(cmd_rdadctmp_16));
    InMux I__6505 (
            .O(N__32147),
            .I(N__32144));
    LocalMux I__6504 (
            .O(N__32144),
            .I(N__32141));
    Span4Mux_h I__6503 (
            .O(N__32141),
            .I(N__32137));
    InMux I__6502 (
            .O(N__32140),
            .I(N__32134));
    Span4Mux_h I__6501 (
            .O(N__32137),
            .I(N__32131));
    LocalMux I__6500 (
            .O(N__32134),
            .I(buf_adcdata1_8));
    Odrv4 I__6499 (
            .O(N__32131),
            .I(buf_adcdata1_8));
    InMux I__6498 (
            .O(N__32126),
            .I(N__32122));
    InMux I__6497 (
            .O(N__32125),
            .I(N__32119));
    LocalMux I__6496 (
            .O(N__32122),
            .I(N__32115));
    LocalMux I__6495 (
            .O(N__32119),
            .I(N__32112));
    InMux I__6494 (
            .O(N__32118),
            .I(N__32109));
    Span4Mux_v I__6493 (
            .O(N__32115),
            .I(N__32105));
    Span4Mux_v I__6492 (
            .O(N__32112),
            .I(N__32101));
    LocalMux I__6491 (
            .O(N__32109),
            .I(N__32098));
    InMux I__6490 (
            .O(N__32108),
            .I(N__32095));
    Span4Mux_h I__6489 (
            .O(N__32105),
            .I(N__32091));
    InMux I__6488 (
            .O(N__32104),
            .I(N__32088));
    Span4Mux_h I__6487 (
            .O(N__32101),
            .I(N__32081));
    Span4Mux_v I__6486 (
            .O(N__32098),
            .I(N__32081));
    LocalMux I__6485 (
            .O(N__32095),
            .I(N__32081));
    InMux I__6484 (
            .O(N__32094),
            .I(N__32078));
    Odrv4 I__6483 (
            .O(N__32091),
            .I(n84));
    LocalMux I__6482 (
            .O(N__32088),
            .I(n84));
    Odrv4 I__6481 (
            .O(N__32081),
            .I(n84));
    LocalMux I__6480 (
            .O(N__32078),
            .I(n84));
    InMux I__6479 (
            .O(N__32069),
            .I(N__32066));
    LocalMux I__6478 (
            .O(N__32066),
            .I(N__32063));
    Span4Mux_h I__6477 (
            .O(N__32063),
            .I(N__32060));
    Odrv4 I__6476 (
            .O(N__32060),
            .I(n15546));
    InMux I__6475 (
            .O(N__32057),
            .I(N__32052));
    InMux I__6474 (
            .O(N__32056),
            .I(N__32049));
    InMux I__6473 (
            .O(N__32055),
            .I(N__32046));
    LocalMux I__6472 (
            .O(N__32052),
            .I(data_index_5));
    LocalMux I__6471 (
            .O(N__32049),
            .I(data_index_5));
    LocalMux I__6470 (
            .O(N__32046),
            .I(data_index_5));
    InMux I__6469 (
            .O(N__32039),
            .I(N__32035));
    InMux I__6468 (
            .O(N__32038),
            .I(N__32032));
    LocalMux I__6467 (
            .O(N__32035),
            .I(N__32026));
    LocalMux I__6466 (
            .O(N__32032),
            .I(N__32026));
    CascadeMux I__6465 (
            .O(N__32031),
            .I(N__32023));
    Span4Mux_v I__6464 (
            .O(N__32026),
            .I(N__32020));
    InMux I__6463 (
            .O(N__32023),
            .I(N__32017));
    Span4Mux_v I__6462 (
            .O(N__32020),
            .I(N__32014));
    LocalMux I__6461 (
            .O(N__32017),
            .I(buf_dds_12));
    Odrv4 I__6460 (
            .O(N__32014),
            .I(buf_dds_12));
    InMux I__6459 (
            .O(N__32009),
            .I(N__32006));
    LocalMux I__6458 (
            .O(N__32006),
            .I(N__32002));
    InMux I__6457 (
            .O(N__32005),
            .I(N__31999));
    Span4Mux_v I__6456 (
            .O(N__32002),
            .I(N__31996));
    LocalMux I__6455 (
            .O(N__31999),
            .I(acadc_skipcnt_2));
    Odrv4 I__6454 (
            .O(N__31996),
            .I(acadc_skipcnt_2));
    InMux I__6453 (
            .O(N__31991),
            .I(N__31988));
    LocalMux I__6452 (
            .O(N__31988),
            .I(N__31983));
    InMux I__6451 (
            .O(N__31987),
            .I(N__31980));
    InMux I__6450 (
            .O(N__31986),
            .I(N__31977));
    Sp12to4 I__6449 (
            .O(N__31983),
            .I(N__31972));
    LocalMux I__6448 (
            .O(N__31980),
            .I(N__31972));
    LocalMux I__6447 (
            .O(N__31977),
            .I(acadc_skipCount_7));
    Odrv12 I__6446 (
            .O(N__31972),
            .I(acadc_skipCount_7));
    CascadeMux I__6445 (
            .O(N__31967),
            .I(N__31964));
    InMux I__6444 (
            .O(N__31964),
            .I(N__31961));
    LocalMux I__6443 (
            .O(N__31961),
            .I(N__31957));
    InMux I__6442 (
            .O(N__31960),
            .I(N__31954));
    Span4Mux_h I__6441 (
            .O(N__31957),
            .I(N__31951));
    LocalMux I__6440 (
            .O(N__31954),
            .I(acadc_skipcnt_7));
    Odrv4 I__6439 (
            .O(N__31951),
            .I(acadc_skipcnt_7));
    InMux I__6438 (
            .O(N__31946),
            .I(N__31942));
    CascadeMux I__6437 (
            .O(N__31945),
            .I(N__31939));
    LocalMux I__6436 (
            .O(N__31942),
            .I(N__31936));
    InMux I__6435 (
            .O(N__31939),
            .I(N__31932));
    Span4Mux_h I__6434 (
            .O(N__31936),
            .I(N__31929));
    InMux I__6433 (
            .O(N__31935),
            .I(N__31926));
    LocalMux I__6432 (
            .O(N__31932),
            .I(acadc_skipCount_2));
    Odrv4 I__6431 (
            .O(N__31929),
            .I(acadc_skipCount_2));
    LocalMux I__6430 (
            .O(N__31926),
            .I(acadc_skipCount_2));
    InMux I__6429 (
            .O(N__31919),
            .I(N__31916));
    LocalMux I__6428 (
            .O(N__31916),
            .I(n22_adj_1170));
    InMux I__6427 (
            .O(N__31913),
            .I(N__31908));
    InMux I__6426 (
            .O(N__31912),
            .I(N__31903));
    InMux I__6425 (
            .O(N__31911),
            .I(N__31903));
    LocalMux I__6424 (
            .O(N__31908),
            .I(N__31900));
    LocalMux I__6423 (
            .O(N__31903),
            .I(req_data_cnt_14));
    Odrv4 I__6422 (
            .O(N__31900),
            .I(req_data_cnt_14));
    InMux I__6421 (
            .O(N__31895),
            .I(N__31892));
    LocalMux I__6420 (
            .O(N__31892),
            .I(n23_adj_1194));
    InMux I__6419 (
            .O(N__31889),
            .I(N__31886));
    LocalMux I__6418 (
            .O(N__31886),
            .I(N__31881));
    InMux I__6417 (
            .O(N__31885),
            .I(N__31876));
    InMux I__6416 (
            .O(N__31884),
            .I(N__31876));
    Odrv4 I__6415 (
            .O(N__31881),
            .I(acadc_skipCount_4));
    LocalMux I__6414 (
            .O(N__31876),
            .I(acadc_skipCount_4));
    InMux I__6413 (
            .O(N__31871),
            .I(N__31866));
    CascadeMux I__6412 (
            .O(N__31870),
            .I(N__31863));
    InMux I__6411 (
            .O(N__31869),
            .I(N__31859));
    LocalMux I__6410 (
            .O(N__31866),
            .I(N__31856));
    InMux I__6409 (
            .O(N__31863),
            .I(N__31853));
    InMux I__6408 (
            .O(N__31862),
            .I(N__31850));
    LocalMux I__6407 (
            .O(N__31859),
            .I(N__31843));
    Span4Mux_h I__6406 (
            .O(N__31856),
            .I(N__31838));
    LocalMux I__6405 (
            .O(N__31853),
            .I(N__31838));
    LocalMux I__6404 (
            .O(N__31850),
            .I(N__31835));
    InMux I__6403 (
            .O(N__31849),
            .I(N__31832));
    InMux I__6402 (
            .O(N__31848),
            .I(N__31829));
    InMux I__6401 (
            .O(N__31847),
            .I(N__31824));
    InMux I__6400 (
            .O(N__31846),
            .I(N__31824));
    Span4Mux_v I__6399 (
            .O(N__31843),
            .I(N__31819));
    Span4Mux_v I__6398 (
            .O(N__31838),
            .I(N__31819));
    Span4Mux_v I__6397 (
            .O(N__31835),
            .I(N__31816));
    LocalMux I__6396 (
            .O(N__31832),
            .I(n9224));
    LocalMux I__6395 (
            .O(N__31829),
            .I(n9224));
    LocalMux I__6394 (
            .O(N__31824),
            .I(n9224));
    Odrv4 I__6393 (
            .O(N__31819),
            .I(n9224));
    Odrv4 I__6392 (
            .O(N__31816),
            .I(n9224));
    InMux I__6391 (
            .O(N__31805),
            .I(N__31802));
    LocalMux I__6390 (
            .O(N__31802),
            .I(N__31799));
    Span4Mux_h I__6389 (
            .O(N__31799),
            .I(N__31795));
    InMux I__6388 (
            .O(N__31798),
            .I(N__31792));
    Span4Mux_v I__6387 (
            .O(N__31795),
            .I(N__31789));
    LocalMux I__6386 (
            .O(N__31792),
            .I(buf_device_acadc_5));
    Odrv4 I__6385 (
            .O(N__31789),
            .I(buf_device_acadc_5));
    InMux I__6384 (
            .O(N__31784),
            .I(N__31775));
    InMux I__6383 (
            .O(N__31783),
            .I(N__31775));
    InMux I__6382 (
            .O(N__31782),
            .I(N__31775));
    LocalMux I__6381 (
            .O(N__31775),
            .I(acadc_skipCount_9));
    InMux I__6380 (
            .O(N__31772),
            .I(N__31769));
    LocalMux I__6379 (
            .O(N__31769),
            .I(N__31766));
    Span4Mux_h I__6378 (
            .O(N__31766),
            .I(N__31763));
    Odrv4 I__6377 (
            .O(N__31763),
            .I(n15834));
    InMux I__6376 (
            .O(N__31760),
            .I(N__31757));
    LocalMux I__6375 (
            .O(N__31757),
            .I(N__31754));
    Span4Mux_v I__6374 (
            .O(N__31754),
            .I(N__31751));
    Span4Mux_h I__6373 (
            .O(N__31751),
            .I(N__31748));
    Odrv4 I__6372 (
            .O(N__31748),
            .I(n19_adj_1234));
    CascadeMux I__6371 (
            .O(N__31745),
            .I(n20_adj_1253_cascade_));
    InMux I__6370 (
            .O(N__31742),
            .I(N__31739));
    LocalMux I__6369 (
            .O(N__31739),
            .I(N__31736));
    Span4Mux_h I__6368 (
            .O(N__31736),
            .I(N__31733));
    Odrv4 I__6367 (
            .O(N__31733),
            .I(n29));
    InMux I__6366 (
            .O(N__31730),
            .I(N__31723));
    InMux I__6365 (
            .O(N__31729),
            .I(N__31723));
    InMux I__6364 (
            .O(N__31728),
            .I(N__31720));
    LocalMux I__6363 (
            .O(N__31723),
            .I(N__31717));
    LocalMux I__6362 (
            .O(N__31720),
            .I(buf_dds_7));
    Odrv4 I__6361 (
            .O(N__31717),
            .I(buf_dds_7));
    CascadeMux I__6360 (
            .O(N__31712),
            .I(N__31709));
    InMux I__6359 (
            .O(N__31709),
            .I(N__31706));
    LocalMux I__6358 (
            .O(N__31706),
            .I(N__31696));
    CascadeMux I__6357 (
            .O(N__31705),
            .I(N__31693));
    CascadeMux I__6356 (
            .O(N__31704),
            .I(N__31690));
    CascadeMux I__6355 (
            .O(N__31703),
            .I(N__31687));
    CascadeMux I__6354 (
            .O(N__31702),
            .I(N__31684));
    CascadeMux I__6353 (
            .O(N__31701),
            .I(N__31681));
    CascadeMux I__6352 (
            .O(N__31700),
            .I(N__31678));
    CascadeMux I__6351 (
            .O(N__31699),
            .I(N__31675));
    Span4Mux_v I__6350 (
            .O(N__31696),
            .I(N__31670));
    InMux I__6349 (
            .O(N__31693),
            .I(N__31663));
    InMux I__6348 (
            .O(N__31690),
            .I(N__31663));
    InMux I__6347 (
            .O(N__31687),
            .I(N__31663));
    InMux I__6346 (
            .O(N__31684),
            .I(N__31654));
    InMux I__6345 (
            .O(N__31681),
            .I(N__31654));
    InMux I__6344 (
            .O(N__31678),
            .I(N__31654));
    InMux I__6343 (
            .O(N__31675),
            .I(N__31654));
    InMux I__6342 (
            .O(N__31674),
            .I(N__31651));
    InMux I__6341 (
            .O(N__31673),
            .I(N__31648));
    Span4Mux_h I__6340 (
            .O(N__31670),
            .I(N__31641));
    LocalMux I__6339 (
            .O(N__31663),
            .I(N__31641));
    LocalMux I__6338 (
            .O(N__31654),
            .I(N__31641));
    LocalMux I__6337 (
            .O(N__31651),
            .I(N__31634));
    LocalMux I__6336 (
            .O(N__31648),
            .I(N__31634));
    Span4Mux_v I__6335 (
            .O(N__31641),
            .I(N__31634));
    Odrv4 I__6334 (
            .O(N__31634),
            .I(n7567));
    InMux I__6333 (
            .O(N__31631),
            .I(N__31628));
    LocalMux I__6332 (
            .O(N__31628),
            .I(n21_adj_1204));
    CascadeMux I__6331 (
            .O(N__31625),
            .I(N__31621));
    InMux I__6330 (
            .O(N__31624),
            .I(N__31618));
    InMux I__6329 (
            .O(N__31621),
            .I(N__31614));
    LocalMux I__6328 (
            .O(N__31618),
            .I(N__31611));
    InMux I__6327 (
            .O(N__31617),
            .I(N__31608));
    LocalMux I__6326 (
            .O(N__31614),
            .I(N__31605));
    Span4Mux_v I__6325 (
            .O(N__31611),
            .I(N__31602));
    LocalMux I__6324 (
            .O(N__31608),
            .I(N__31599));
    Span4Mux_v I__6323 (
            .O(N__31605),
            .I(N__31594));
    Span4Mux_h I__6322 (
            .O(N__31602),
            .I(N__31589));
    Span4Mux_v I__6321 (
            .O(N__31599),
            .I(N__31589));
    InMux I__6320 (
            .O(N__31598),
            .I(N__31584));
    InMux I__6319 (
            .O(N__31597),
            .I(N__31584));
    Odrv4 I__6318 (
            .O(N__31594),
            .I(comm_buf_1_4));
    Odrv4 I__6317 (
            .O(N__31589),
            .I(comm_buf_1_4));
    LocalMux I__6316 (
            .O(N__31584),
            .I(comm_buf_1_4));
    InMux I__6315 (
            .O(N__31577),
            .I(N__31572));
    InMux I__6314 (
            .O(N__31576),
            .I(N__31569));
    InMux I__6313 (
            .O(N__31575),
            .I(N__31566));
    LocalMux I__6312 (
            .O(N__31572),
            .I(N__31563));
    LocalMux I__6311 (
            .O(N__31569),
            .I(N__31560));
    LocalMux I__6310 (
            .O(N__31566),
            .I(buf_dds_4));
    Odrv12 I__6309 (
            .O(N__31563),
            .I(buf_dds_4));
    Odrv4 I__6308 (
            .O(N__31560),
            .I(buf_dds_4));
    CascadeMux I__6307 (
            .O(N__31553),
            .I(N__31550));
    InMux I__6306 (
            .O(N__31550),
            .I(N__31546));
    InMux I__6305 (
            .O(N__31549),
            .I(N__31543));
    LocalMux I__6304 (
            .O(N__31546),
            .I(N__31540));
    LocalMux I__6303 (
            .O(N__31543),
            .I(buf_control_5));
    Odrv4 I__6302 (
            .O(N__31540),
            .I(buf_control_5));
    InMux I__6301 (
            .O(N__31535),
            .I(N__31532));
    LocalMux I__6300 (
            .O(N__31532),
            .I(N__31529));
    Span4Mux_h I__6299 (
            .O(N__31529),
            .I(N__31526));
    Span4Mux_h I__6298 (
            .O(N__31526),
            .I(N__31523));
    Odrv4 I__6297 (
            .O(N__31523),
            .I(buf_data1_10));
    CascadeMux I__6296 (
            .O(N__31520),
            .I(n4195_cascade_));
    InMux I__6295 (
            .O(N__31517),
            .I(N__31514));
    LocalMux I__6294 (
            .O(N__31514),
            .I(n4232));
    InMux I__6293 (
            .O(N__31511),
            .I(N__31508));
    LocalMux I__6292 (
            .O(N__31508),
            .I(N__31504));
    InMux I__6291 (
            .O(N__31507),
            .I(N__31501));
    Span4Mux_h I__6290 (
            .O(N__31504),
            .I(N__31498));
    LocalMux I__6289 (
            .O(N__31501),
            .I(acadc_skipcnt_9));
    Odrv4 I__6288 (
            .O(N__31498),
            .I(acadc_skipcnt_9));
    CascadeMux I__6287 (
            .O(N__31493),
            .I(N__31490));
    InMux I__6286 (
            .O(N__31490),
            .I(N__31487));
    LocalMux I__6285 (
            .O(N__31487),
            .I(N__31483));
    InMux I__6284 (
            .O(N__31486),
            .I(N__31480));
    Span12Mux_v I__6283 (
            .O(N__31483),
            .I(N__31477));
    LocalMux I__6282 (
            .O(N__31480),
            .I(acadc_skipcnt_15));
    Odrv12 I__6281 (
            .O(N__31477),
            .I(acadc_skipcnt_15));
    InMux I__6280 (
            .O(N__31472),
            .I(N__31469));
    LocalMux I__6279 (
            .O(N__31469),
            .I(n24_adj_1174));
    InMux I__6278 (
            .O(N__31466),
            .I(N__31463));
    LocalMux I__6277 (
            .O(N__31463),
            .I(n4247));
    InMux I__6276 (
            .O(N__31460),
            .I(N__31457));
    LocalMux I__6275 (
            .O(N__31457),
            .I(N__31453));
    InMux I__6274 (
            .O(N__31456),
            .I(N__31449));
    Span4Mux_v I__6273 (
            .O(N__31453),
            .I(N__31446));
    InMux I__6272 (
            .O(N__31452),
            .I(N__31443));
    LocalMux I__6271 (
            .O(N__31449),
            .I(N__31440));
    Span4Mux_v I__6270 (
            .O(N__31446),
            .I(N__31437));
    LocalMux I__6269 (
            .O(N__31443),
            .I(buf_dds_15));
    Odrv4 I__6268 (
            .O(N__31440),
            .I(buf_dds_15));
    Odrv4 I__6267 (
            .O(N__31437),
            .I(buf_dds_15));
    InMux I__6266 (
            .O(N__31430),
            .I(N__31427));
    LocalMux I__6265 (
            .O(N__31427),
            .I(N__31424));
    Span12Mux_v I__6264 (
            .O(N__31424),
            .I(N__31419));
    InMux I__6263 (
            .O(N__31423),
            .I(N__31414));
    InMux I__6262 (
            .O(N__31422),
            .I(N__31414));
    Odrv12 I__6261 (
            .O(N__31419),
            .I(req_data_cnt_13));
    LocalMux I__6260 (
            .O(N__31414),
            .I(req_data_cnt_13));
    InMux I__6259 (
            .O(N__31409),
            .I(N__31404));
    InMux I__6258 (
            .O(N__31408),
            .I(N__31399));
    InMux I__6257 (
            .O(N__31407),
            .I(N__31399));
    LocalMux I__6256 (
            .O(N__31404),
            .I(req_data_cnt_8));
    LocalMux I__6255 (
            .O(N__31399),
            .I(req_data_cnt_8));
    CascadeMux I__6254 (
            .O(N__31394),
            .I(N__31391));
    InMux I__6253 (
            .O(N__31391),
            .I(N__31388));
    LocalMux I__6252 (
            .O(N__31388),
            .I(N__31385));
    Odrv12 I__6251 (
            .O(N__31385),
            .I(n15812));
    InMux I__6250 (
            .O(N__31382),
            .I(N__31379));
    LocalMux I__6249 (
            .O(N__31379),
            .I(N__31375));
    InMux I__6248 (
            .O(N__31378),
            .I(N__31372));
    Span4Mux_v I__6247 (
            .O(N__31375),
            .I(N__31369));
    LocalMux I__6246 (
            .O(N__31372),
            .I(buf_device_acadc_6));
    Odrv4 I__6245 (
            .O(N__31369),
            .I(buf_device_acadc_6));
    CascadeMux I__6244 (
            .O(N__31364),
            .I(N__31361));
    InMux I__6243 (
            .O(N__31361),
            .I(N__31358));
    LocalMux I__6242 (
            .O(N__31358),
            .I(N__31355));
    Span4Mux_h I__6241 (
            .O(N__31355),
            .I(N__31352));
    Odrv4 I__6240 (
            .O(N__31352),
            .I(buf_data1_16));
    InMux I__6239 (
            .O(N__31349),
            .I(N__31346));
    LocalMux I__6238 (
            .O(N__31346),
            .I(N__31343));
    Span4Mux_h I__6237 (
            .O(N__31343),
            .I(N__31340));
    Odrv4 I__6236 (
            .O(N__31340),
            .I(n99));
    CascadeMux I__6235 (
            .O(N__31337),
            .I(N__31332));
    InMux I__6234 (
            .O(N__31336),
            .I(N__31329));
    InMux I__6233 (
            .O(N__31335),
            .I(N__31326));
    InMux I__6232 (
            .O(N__31332),
            .I(N__31323));
    LocalMux I__6231 (
            .O(N__31329),
            .I(req_data_cnt_7));
    LocalMux I__6230 (
            .O(N__31326),
            .I(req_data_cnt_7));
    LocalMux I__6229 (
            .O(N__31323),
            .I(req_data_cnt_7));
    InMux I__6228 (
            .O(N__31316),
            .I(N__31313));
    LocalMux I__6227 (
            .O(N__31313),
            .I(N__31310));
    Odrv4 I__6226 (
            .O(N__31310),
            .I(n4214));
    CascadeMux I__6225 (
            .O(N__31307),
            .I(N__31304));
    InMux I__6224 (
            .O(N__31304),
            .I(N__31301));
    LocalMux I__6223 (
            .O(N__31301),
            .I(N__31298));
    Span4Mux_v I__6222 (
            .O(N__31298),
            .I(N__31295));
    Odrv4 I__6221 (
            .O(N__31295),
            .I(n15556));
    InMux I__6220 (
            .O(N__31292),
            .I(N__31289));
    LocalMux I__6219 (
            .O(N__31289),
            .I(N__31286));
    Span12Mux_h I__6218 (
            .O(N__31286),
            .I(N__31283));
    Odrv12 I__6217 (
            .O(N__31283),
            .I(n60_adj_1157));
    InMux I__6216 (
            .O(N__31280),
            .I(N__31277));
    LocalMux I__6215 (
            .O(N__31277),
            .I(N__31274));
    Odrv4 I__6214 (
            .O(N__31274),
            .I(n4252));
    CascadeMux I__6213 (
            .O(N__31271),
            .I(N__31268));
    InMux I__6212 (
            .O(N__31268),
            .I(N__31265));
    LocalMux I__6211 (
            .O(N__31265),
            .I(n4202));
    CascadeMux I__6210 (
            .O(N__31262),
            .I(N__31259));
    InMux I__6209 (
            .O(N__31259),
            .I(N__31256));
    LocalMux I__6208 (
            .O(N__31256),
            .I(\CLOCK_DDS.tmp_buf_2 ));
    InMux I__6207 (
            .O(N__31253),
            .I(N__31250));
    LocalMux I__6206 (
            .O(N__31250),
            .I(N__31247));
    Odrv4 I__6205 (
            .O(N__31247),
            .I(\CLOCK_DDS.tmp_buf_3 ));
    CascadeMux I__6204 (
            .O(N__31244),
            .I(N__31241));
    InMux I__6203 (
            .O(N__31241),
            .I(N__31238));
    LocalMux I__6202 (
            .O(N__31238),
            .I(\CLOCK_DDS.tmp_buf_4 ));
    CascadeMux I__6201 (
            .O(N__31235),
            .I(N__31232));
    InMux I__6200 (
            .O(N__31232),
            .I(N__31229));
    LocalMux I__6199 (
            .O(N__31229),
            .I(\CLOCK_DDS.tmp_buf_5 ));
    CascadeMux I__6198 (
            .O(N__31226),
            .I(N__31223));
    InMux I__6197 (
            .O(N__31223),
            .I(N__31220));
    LocalMux I__6196 (
            .O(N__31220),
            .I(\CLOCK_DDS.tmp_buf_6 ));
    InMux I__6195 (
            .O(N__31217),
            .I(N__31214));
    LocalMux I__6194 (
            .O(N__31214),
            .I(\CLOCK_DDS.tmp_buf_7 ));
    CEMux I__6193 (
            .O(N__31211),
            .I(N__31206));
    CEMux I__6192 (
            .O(N__31210),
            .I(N__31203));
    CEMux I__6191 (
            .O(N__31209),
            .I(N__31200));
    LocalMux I__6190 (
            .O(N__31206),
            .I(\CLOCK_DDS.n9759 ));
    LocalMux I__6189 (
            .O(N__31203),
            .I(\CLOCK_DDS.n9759 ));
    LocalMux I__6188 (
            .O(N__31200),
            .I(\CLOCK_DDS.n9759 ));
    SRMux I__6187 (
            .O(N__31193),
            .I(N__31190));
    LocalMux I__6186 (
            .O(N__31190),
            .I(N__31186));
    InMux I__6185 (
            .O(N__31189),
            .I(N__31183));
    Span4Mux_v I__6184 (
            .O(N__31186),
            .I(N__31180));
    LocalMux I__6183 (
            .O(N__31183),
            .I(N__31177));
    Span4Mux_h I__6182 (
            .O(N__31180),
            .I(N__31174));
    Span4Mux_h I__6181 (
            .O(N__31177),
            .I(N__31171));
    Odrv4 I__6180 (
            .O(N__31174),
            .I(n10823));
    Odrv4 I__6179 (
            .O(N__31171),
            .I(n10823));
    CEMux I__6178 (
            .O(N__31166),
            .I(N__31163));
    LocalMux I__6177 (
            .O(N__31163),
            .I(N__31160));
    Span4Mux_h I__6176 (
            .O(N__31160),
            .I(N__31157));
    Span4Mux_v I__6175 (
            .O(N__31157),
            .I(N__31154));
    Odrv4 I__6174 (
            .O(N__31154),
            .I(\CLOCK_DDS.n9_adj_1021 ));
    InMux I__6173 (
            .O(N__31151),
            .I(N__31148));
    LocalMux I__6172 (
            .O(N__31148),
            .I(N__31145));
    Span4Mux_v I__6171 (
            .O(N__31145),
            .I(N__31139));
    InMux I__6170 (
            .O(N__31144),
            .I(N__31132));
    InMux I__6169 (
            .O(N__31143),
            .I(N__31132));
    InMux I__6168 (
            .O(N__31142),
            .I(N__31132));
    Span4Mux_h I__6167 (
            .O(N__31139),
            .I(N__31129));
    LocalMux I__6166 (
            .O(N__31132),
            .I(bit_cnt_1));
    Odrv4 I__6165 (
            .O(N__31129),
            .I(bit_cnt_1));
    InMux I__6164 (
            .O(N__31124),
            .I(N__31120));
    InMux I__6163 (
            .O(N__31123),
            .I(N__31117));
    LocalMux I__6162 (
            .O(N__31120),
            .I(N__31112));
    LocalMux I__6161 (
            .O(N__31117),
            .I(N__31112));
    Odrv12 I__6160 (
            .O(N__31112),
            .I(n15176));
    InMux I__6159 (
            .O(N__31109),
            .I(N__31106));
    LocalMux I__6158 (
            .O(N__31106),
            .I(N__31103));
    Span4Mux_v I__6157 (
            .O(N__31103),
            .I(N__31100));
    Sp12to4 I__6156 (
            .O(N__31100),
            .I(N__31097));
    Odrv12 I__6155 (
            .O(N__31097),
            .I(n15396));
    CascadeMux I__6154 (
            .O(N__31094),
            .I(N__31091));
    InMux I__6153 (
            .O(N__31091),
            .I(N__31088));
    LocalMux I__6152 (
            .O(N__31088),
            .I(N__31085));
    Odrv4 I__6151 (
            .O(N__31085),
            .I(n15670));
    InMux I__6150 (
            .O(N__31082),
            .I(N__31079));
    LocalMux I__6149 (
            .O(N__31079),
            .I(N__31076));
    Span4Mux_h I__6148 (
            .O(N__31076),
            .I(N__31070));
    InMux I__6147 (
            .O(N__31075),
            .I(N__31065));
    InMux I__6146 (
            .O(N__31074),
            .I(N__31065));
    InMux I__6145 (
            .O(N__31073),
            .I(N__31062));
    Odrv4 I__6144 (
            .O(N__31070),
            .I(n13475));
    LocalMux I__6143 (
            .O(N__31065),
            .I(n13475));
    LocalMux I__6142 (
            .O(N__31062),
            .I(n13475));
    InMux I__6141 (
            .O(N__31055),
            .I(N__31052));
    LocalMux I__6140 (
            .O(N__31052),
            .I(N__31049));
    Odrv4 I__6139 (
            .O(N__31049),
            .I(n15_adj_1203));
    InMux I__6138 (
            .O(N__31046),
            .I(N__31043));
    LocalMux I__6137 (
            .O(N__31043),
            .I(N__31040));
    Span4Mux_v I__6136 (
            .O(N__31040),
            .I(N__31037));
    Span4Mux_h I__6135 (
            .O(N__31037),
            .I(N__31033));
    InMux I__6134 (
            .O(N__31036),
            .I(N__31030));
    Odrv4 I__6133 (
            .O(N__31033),
            .I(tmp_buf_15));
    LocalMux I__6132 (
            .O(N__31030),
            .I(tmp_buf_15));
    CascadeMux I__6131 (
            .O(N__31025),
            .I(N__31022));
    InMux I__6130 (
            .O(N__31022),
            .I(N__31019));
    LocalMux I__6129 (
            .O(N__31019),
            .I(\CLOCK_DDS.tmp_buf_0 ));
    CascadeMux I__6128 (
            .O(N__31016),
            .I(N__31013));
    InMux I__6127 (
            .O(N__31013),
            .I(N__31010));
    LocalMux I__6126 (
            .O(N__31010),
            .I(\CLOCK_DDS.tmp_buf_1 ));
    SRMux I__6125 (
            .O(N__31007),
            .I(N__31004));
    LocalMux I__6124 (
            .O(N__31004),
            .I(N__31001));
    Span4Mux_v I__6123 (
            .O(N__31001),
            .I(N__30997));
    SRMux I__6122 (
            .O(N__31000),
            .I(N__30993));
    Sp12to4 I__6121 (
            .O(N__30997),
            .I(N__30990));
    SRMux I__6120 (
            .O(N__30996),
            .I(N__30987));
    LocalMux I__6119 (
            .O(N__30993),
            .I(N__30984));
    Span12Mux_h I__6118 (
            .O(N__30990),
            .I(N__30979));
    LocalMux I__6117 (
            .O(N__30987),
            .I(N__30979));
    Span4Mux_h I__6116 (
            .O(N__30984),
            .I(N__30976));
    Odrv12 I__6115 (
            .O(N__30979),
            .I(\comm_spi.data_tx_7__N_813 ));
    Odrv4 I__6114 (
            .O(N__30976),
            .I(\comm_spi.data_tx_7__N_813 ));
    InMux I__6113 (
            .O(N__30971),
            .I(N__30968));
    LocalMux I__6112 (
            .O(N__30968),
            .I(N__30964));
    InMux I__6111 (
            .O(N__30967),
            .I(N__30961));
    Span4Mux_v I__6110 (
            .O(N__30964),
            .I(N__30958));
    LocalMux I__6109 (
            .O(N__30961),
            .I(N__30955));
    Span4Mux_h I__6108 (
            .O(N__30958),
            .I(N__30951));
    Span4Mux_v I__6107 (
            .O(N__30955),
            .I(N__30948));
    InMux I__6106 (
            .O(N__30954),
            .I(N__30945));
    Sp12to4 I__6105 (
            .O(N__30951),
            .I(N__30938));
    Sp12to4 I__6104 (
            .O(N__30948),
            .I(N__30938));
    LocalMux I__6103 (
            .O(N__30945),
            .I(N__30938));
    Span12Mux_h I__6102 (
            .O(N__30938),
            .I(N__30935));
    Odrv12 I__6101 (
            .O(N__30935),
            .I(comm_tx_buf_3));
    SRMux I__6100 (
            .O(N__30932),
            .I(N__30929));
    LocalMux I__6099 (
            .O(N__30929),
            .I(N__30926));
    Span4Mux_v I__6098 (
            .O(N__30926),
            .I(N__30923));
    Span4Mux_h I__6097 (
            .O(N__30923),
            .I(N__30920));
    Odrv4 I__6096 (
            .O(N__30920),
            .I(\comm_spi.data_tx_7__N_825 ));
    InMux I__6095 (
            .O(N__30917),
            .I(N__30914));
    LocalMux I__6094 (
            .O(N__30914),
            .I(N__30911));
    Span4Mux_v I__6093 (
            .O(N__30911),
            .I(N__30908));
    Span4Mux_h I__6092 (
            .O(N__30908),
            .I(N__30905));
    Odrv4 I__6091 (
            .O(N__30905),
            .I(buf_data1_22));
    InMux I__6090 (
            .O(N__30902),
            .I(N__30899));
    LocalMux I__6089 (
            .O(N__30899),
            .I(N__30896));
    Span12Mux_h I__6088 (
            .O(N__30896),
            .I(N__30893));
    Odrv12 I__6087 (
            .O(N__30893),
            .I(n66));
    InMux I__6086 (
            .O(N__30890),
            .I(N__30887));
    LocalMux I__6085 (
            .O(N__30887),
            .I(N__30883));
    InMux I__6084 (
            .O(N__30886),
            .I(N__30880));
    Span4Mux_h I__6083 (
            .O(N__30883),
            .I(N__30877));
    LocalMux I__6082 (
            .O(N__30880),
            .I(N__30874));
    Span4Mux_h I__6081 (
            .O(N__30877),
            .I(N__30871));
    Span12Mux_h I__6080 (
            .O(N__30874),
            .I(N__30868));
    Odrv4 I__6079 (
            .O(N__30871),
            .I(\comm_spi.n10452 ));
    Odrv12 I__6078 (
            .O(N__30868),
            .I(\comm_spi.n10452 ));
    InMux I__6077 (
            .O(N__30863),
            .I(N__30860));
    LocalMux I__6076 (
            .O(N__30860),
            .I(N__30857));
    Span4Mux_v I__6075 (
            .O(N__30857),
            .I(N__30853));
    InMux I__6074 (
            .O(N__30856),
            .I(N__30850));
    Odrv4 I__6073 (
            .O(N__30853),
            .I(\comm_spi.n10451 ));
    LocalMux I__6072 (
            .O(N__30850),
            .I(\comm_spi.n10451 ));
    InMux I__6071 (
            .O(N__30845),
            .I(N__30839));
    InMux I__6070 (
            .O(N__30844),
            .I(N__30836));
    InMux I__6069 (
            .O(N__30843),
            .I(N__30831));
    InMux I__6068 (
            .O(N__30842),
            .I(N__30828));
    LocalMux I__6067 (
            .O(N__30839),
            .I(N__30825));
    LocalMux I__6066 (
            .O(N__30836),
            .I(N__30822));
    InMux I__6065 (
            .O(N__30835),
            .I(N__30819));
    InMux I__6064 (
            .O(N__30834),
            .I(N__30816));
    LocalMux I__6063 (
            .O(N__30831),
            .I(N__30813));
    LocalMux I__6062 (
            .O(N__30828),
            .I(N__30810));
    Span12Mux_v I__6061 (
            .O(N__30825),
            .I(N__30807));
    Span4Mux_v I__6060 (
            .O(N__30822),
            .I(N__30800));
    LocalMux I__6059 (
            .O(N__30819),
            .I(N__30800));
    LocalMux I__6058 (
            .O(N__30816),
            .I(N__30800));
    Span4Mux_v I__6057 (
            .O(N__30813),
            .I(N__30795));
    Span4Mux_h I__6056 (
            .O(N__30810),
            .I(N__30795));
    Odrv12 I__6055 (
            .O(N__30807),
            .I(\comm_spi.n10444 ));
    Odrv4 I__6054 (
            .O(N__30800),
            .I(\comm_spi.n10444 ));
    Odrv4 I__6053 (
            .O(N__30795),
            .I(\comm_spi.n10444 ));
    InMux I__6052 (
            .O(N__30788),
            .I(N__30785));
    LocalMux I__6051 (
            .O(N__30785),
            .I(N__30782));
    Odrv4 I__6050 (
            .O(N__30782),
            .I(\comm_spi.n10445 ));
    SRMux I__6049 (
            .O(N__30779),
            .I(N__30775));
    SRMux I__6048 (
            .O(N__30778),
            .I(N__30772));
    LocalMux I__6047 (
            .O(N__30775),
            .I(N__30769));
    LocalMux I__6046 (
            .O(N__30772),
            .I(N__30765));
    Span4Mux_h I__6045 (
            .O(N__30769),
            .I(N__30762));
    SRMux I__6044 (
            .O(N__30768),
            .I(N__30759));
    Span4Mux_h I__6043 (
            .O(N__30765),
            .I(N__30756));
    Span4Mux_h I__6042 (
            .O(N__30762),
            .I(N__30751));
    LocalMux I__6041 (
            .O(N__30759),
            .I(N__30751));
    Span4Mux_h I__6040 (
            .O(N__30756),
            .I(N__30748));
    Odrv4 I__6039 (
            .O(N__30751),
            .I(\comm_spi.data_tx_7__N_805 ));
    Odrv4 I__6038 (
            .O(N__30748),
            .I(\comm_spi.data_tx_7__N_805 ));
    SRMux I__6037 (
            .O(N__30743),
            .I(N__30740));
    LocalMux I__6036 (
            .O(N__30740),
            .I(N__30737));
    Span4Mux_h I__6035 (
            .O(N__30737),
            .I(N__30733));
    SRMux I__6034 (
            .O(N__30736),
            .I(N__30730));
    Span4Mux_h I__6033 (
            .O(N__30733),
            .I(N__30727));
    LocalMux I__6032 (
            .O(N__30730),
            .I(N__30724));
    Span4Mux_h I__6031 (
            .O(N__30727),
            .I(N__30721));
    Span4Mux_h I__6030 (
            .O(N__30724),
            .I(N__30718));
    Sp12to4 I__6029 (
            .O(N__30721),
            .I(N__30715));
    Span4Mux_h I__6028 (
            .O(N__30718),
            .I(N__30712));
    Odrv12 I__6027 (
            .O(N__30715),
            .I(n10640));
    Odrv4 I__6026 (
            .O(N__30712),
            .I(n10640));
    SRMux I__6025 (
            .O(N__30707),
            .I(N__30704));
    LocalMux I__6024 (
            .O(N__30704),
            .I(N__30700));
    SRMux I__6023 (
            .O(N__30703),
            .I(N__30697));
    Span4Mux_v I__6022 (
            .O(N__30700),
            .I(N__30692));
    LocalMux I__6021 (
            .O(N__30697),
            .I(N__30692));
    Sp12to4 I__6020 (
            .O(N__30692),
            .I(N__30689));
    Odrv12 I__6019 (
            .O(N__30689),
            .I(n10532));
    SRMux I__6018 (
            .O(N__30686),
            .I(N__30683));
    LocalMux I__6017 (
            .O(N__30683),
            .I(N__30680));
    Span4Mux_h I__6016 (
            .O(N__30680),
            .I(N__30677));
    Odrv4 I__6015 (
            .O(N__30677),
            .I(n15344));
    InMux I__6014 (
            .O(N__30674),
            .I(N__30671));
    LocalMux I__6013 (
            .O(N__30671),
            .I(N__30668));
    Span12Mux_h I__6012 (
            .O(N__30668),
            .I(N__30665));
    Odrv12 I__6011 (
            .O(N__30665),
            .I(n15171));
    CascadeMux I__6010 (
            .O(N__30662),
            .I(n15328_cascade_));
    InMux I__6009 (
            .O(N__30659),
            .I(N__30649));
    InMux I__6008 (
            .O(N__30658),
            .I(N__30649));
    InMux I__6007 (
            .O(N__30657),
            .I(N__30642));
    InMux I__6006 (
            .O(N__30656),
            .I(N__30642));
    InMux I__6005 (
            .O(N__30655),
            .I(N__30637));
    InMux I__6004 (
            .O(N__30654),
            .I(N__30637));
    LocalMux I__6003 (
            .O(N__30649),
            .I(N__30633));
    InMux I__6002 (
            .O(N__30648),
            .I(N__30630));
    InMux I__6001 (
            .O(N__30647),
            .I(N__30627));
    LocalMux I__6000 (
            .O(N__30642),
            .I(N__30622));
    LocalMux I__5999 (
            .O(N__30637),
            .I(N__30622));
    InMux I__5998 (
            .O(N__30636),
            .I(N__30619));
    Span4Mux_h I__5997 (
            .O(N__30633),
            .I(N__30615));
    LocalMux I__5996 (
            .O(N__30630),
            .I(N__30610));
    LocalMux I__5995 (
            .O(N__30627),
            .I(N__30610));
    Span4Mux_v I__5994 (
            .O(N__30622),
            .I(N__30605));
    LocalMux I__5993 (
            .O(N__30619),
            .I(N__30605));
    InMux I__5992 (
            .O(N__30618),
            .I(N__30601));
    Span4Mux_v I__5991 (
            .O(N__30615),
            .I(N__30598));
    Span4Mux_h I__5990 (
            .O(N__30610),
            .I(N__30595));
    Span4Mux_h I__5989 (
            .O(N__30605),
            .I(N__30592));
    InMux I__5988 (
            .O(N__30604),
            .I(N__30589));
    LocalMux I__5987 (
            .O(N__30601),
            .I(acadc_trig));
    Odrv4 I__5986 (
            .O(N__30598),
            .I(acadc_trig));
    Odrv4 I__5985 (
            .O(N__30595),
            .I(acadc_trig));
    Odrv4 I__5984 (
            .O(N__30592),
            .I(acadc_trig));
    LocalMux I__5983 (
            .O(N__30589),
            .I(acadc_trig));
    InMux I__5982 (
            .O(N__30578),
            .I(N__30573));
    InMux I__5981 (
            .O(N__30577),
            .I(N__30570));
    InMux I__5980 (
            .O(N__30576),
            .I(N__30567));
    LocalMux I__5979 (
            .O(N__30573),
            .I(N__30560));
    LocalMux I__5978 (
            .O(N__30570),
            .I(N__30560));
    LocalMux I__5977 (
            .O(N__30567),
            .I(N__30560));
    Span4Mux_v I__5976 (
            .O(N__30560),
            .I(N__30557));
    Span4Mux_v I__5975 (
            .O(N__30557),
            .I(N__30554));
    Odrv4 I__5974 (
            .O(N__30554),
            .I(data_index_6));
    InMux I__5973 (
            .O(N__30551),
            .I(N__30548));
    LocalMux I__5972 (
            .O(N__30548),
            .I(N__30545));
    Odrv12 I__5971 (
            .O(N__30545),
            .I(n8_adj_1221));
    InMux I__5970 (
            .O(N__30542),
            .I(N__30538));
    InMux I__5969 (
            .O(N__30541),
            .I(N__30535));
    LocalMux I__5968 (
            .O(N__30538),
            .I(N__30532));
    LocalMux I__5967 (
            .O(N__30535),
            .I(N__30529));
    Odrv12 I__5966 (
            .O(N__30532),
            .I(n7_adj_1220));
    Odrv4 I__5965 (
            .O(N__30529),
            .I(n7_adj_1220));
    CascadeMux I__5964 (
            .O(N__30524),
            .I(N__30521));
    CascadeBuf I__5963 (
            .O(N__30521),
            .I(N__30518));
    CascadeMux I__5962 (
            .O(N__30518),
            .I(N__30515));
    CascadeBuf I__5961 (
            .O(N__30515),
            .I(N__30512));
    CascadeMux I__5960 (
            .O(N__30512),
            .I(N__30509));
    CascadeBuf I__5959 (
            .O(N__30509),
            .I(N__30506));
    CascadeMux I__5958 (
            .O(N__30506),
            .I(N__30503));
    CascadeBuf I__5957 (
            .O(N__30503),
            .I(N__30500));
    CascadeMux I__5956 (
            .O(N__30500),
            .I(N__30497));
    CascadeBuf I__5955 (
            .O(N__30497),
            .I(N__30494));
    CascadeMux I__5954 (
            .O(N__30494),
            .I(N__30491));
    CascadeBuf I__5953 (
            .O(N__30491),
            .I(N__30488));
    CascadeMux I__5952 (
            .O(N__30488),
            .I(N__30485));
    CascadeBuf I__5951 (
            .O(N__30485),
            .I(N__30482));
    CascadeMux I__5950 (
            .O(N__30482),
            .I(N__30478));
    CascadeMux I__5949 (
            .O(N__30481),
            .I(N__30475));
    CascadeBuf I__5948 (
            .O(N__30478),
            .I(N__30472));
    CascadeBuf I__5947 (
            .O(N__30475),
            .I(N__30469));
    CascadeMux I__5946 (
            .O(N__30472),
            .I(N__30466));
    CascadeMux I__5945 (
            .O(N__30469),
            .I(N__30463));
    CascadeBuf I__5944 (
            .O(N__30466),
            .I(N__30460));
    InMux I__5943 (
            .O(N__30463),
            .I(N__30457));
    CascadeMux I__5942 (
            .O(N__30460),
            .I(N__30454));
    LocalMux I__5941 (
            .O(N__30457),
            .I(N__30451));
    InMux I__5940 (
            .O(N__30454),
            .I(N__30448));
    Span12Mux_h I__5939 (
            .O(N__30451),
            .I(N__30445));
    LocalMux I__5938 (
            .O(N__30448),
            .I(N__30442));
    Span12Mux_v I__5937 (
            .O(N__30445),
            .I(N__30439));
    Span4Mux_h I__5936 (
            .O(N__30442),
            .I(N__30436));
    Odrv12 I__5935 (
            .O(N__30439),
            .I(data_index_9_N_258_7));
    Odrv4 I__5934 (
            .O(N__30436),
            .I(data_index_9_N_258_7));
    InMux I__5933 (
            .O(N__30431),
            .I(N__30428));
    LocalMux I__5932 (
            .O(N__30428),
            .I(N__30425));
    Span4Mux_v I__5931 (
            .O(N__30425),
            .I(N__30421));
    InMux I__5930 (
            .O(N__30424),
            .I(N__30418));
    Span4Mux_v I__5929 (
            .O(N__30421),
            .I(N__30413));
    LocalMux I__5928 (
            .O(N__30418),
            .I(N__30413));
    Odrv4 I__5927 (
            .O(N__30413),
            .I(n7_adj_1222));
    CascadeMux I__5926 (
            .O(N__30410),
            .I(N__30407));
    InMux I__5925 (
            .O(N__30407),
            .I(N__30404));
    LocalMux I__5924 (
            .O(N__30404),
            .I(N__30401));
    Span4Mux_h I__5923 (
            .O(N__30401),
            .I(N__30398));
    Span4Mux_v I__5922 (
            .O(N__30398),
            .I(N__30394));
    CascadeMux I__5921 (
            .O(N__30397),
            .I(N__30391));
    Span4Mux_v I__5920 (
            .O(N__30394),
            .I(N__30388));
    InMux I__5919 (
            .O(N__30391),
            .I(N__30385));
    Odrv4 I__5918 (
            .O(N__30388),
            .I(n8_adj_1223));
    LocalMux I__5917 (
            .O(N__30385),
            .I(n8_adj_1223));
    CascadeMux I__5916 (
            .O(N__30380),
            .I(N__30377));
    CascadeBuf I__5915 (
            .O(N__30377),
            .I(N__30374));
    CascadeMux I__5914 (
            .O(N__30374),
            .I(N__30371));
    CascadeBuf I__5913 (
            .O(N__30371),
            .I(N__30368));
    CascadeMux I__5912 (
            .O(N__30368),
            .I(N__30365));
    CascadeBuf I__5911 (
            .O(N__30365),
            .I(N__30362));
    CascadeMux I__5910 (
            .O(N__30362),
            .I(N__30359));
    CascadeBuf I__5909 (
            .O(N__30359),
            .I(N__30356));
    CascadeMux I__5908 (
            .O(N__30356),
            .I(N__30353));
    CascadeBuf I__5907 (
            .O(N__30353),
            .I(N__30350));
    CascadeMux I__5906 (
            .O(N__30350),
            .I(N__30347));
    CascadeBuf I__5905 (
            .O(N__30347),
            .I(N__30344));
    CascadeMux I__5904 (
            .O(N__30344),
            .I(N__30341));
    CascadeBuf I__5903 (
            .O(N__30341),
            .I(N__30337));
    CascadeMux I__5902 (
            .O(N__30340),
            .I(N__30334));
    CascadeMux I__5901 (
            .O(N__30337),
            .I(N__30331));
    CascadeBuf I__5900 (
            .O(N__30334),
            .I(N__30328));
    CascadeBuf I__5899 (
            .O(N__30331),
            .I(N__30325));
    CascadeMux I__5898 (
            .O(N__30328),
            .I(N__30322));
    CascadeMux I__5897 (
            .O(N__30325),
            .I(N__30319));
    InMux I__5896 (
            .O(N__30322),
            .I(N__30316));
    CascadeBuf I__5895 (
            .O(N__30319),
            .I(N__30313));
    LocalMux I__5894 (
            .O(N__30316),
            .I(N__30310));
    CascadeMux I__5893 (
            .O(N__30313),
            .I(N__30307));
    Span12Mux_s9_h I__5892 (
            .O(N__30310),
            .I(N__30304));
    InMux I__5891 (
            .O(N__30307),
            .I(N__30301));
    Span12Mux_v I__5890 (
            .O(N__30304),
            .I(N__30298));
    LocalMux I__5889 (
            .O(N__30301),
            .I(N__30295));
    Odrv12 I__5888 (
            .O(N__30298),
            .I(data_index_9_N_258_6));
    Odrv12 I__5887 (
            .O(N__30295),
            .I(data_index_9_N_258_6));
    IoInMux I__5886 (
            .O(N__30290),
            .I(N__30287));
    LocalMux I__5885 (
            .O(N__30287),
            .I(N__30284));
    Span4Mux_s3_h I__5884 (
            .O(N__30284),
            .I(N__30281));
    Sp12to4 I__5883 (
            .O(N__30281),
            .I(N__30278));
    Span12Mux_s9_v I__5882 (
            .O(N__30278),
            .I(N__30275));
    Odrv12 I__5881 (
            .O(N__30275),
            .I(ICE_SPI_MISO));
    InMux I__5880 (
            .O(N__30272),
            .I(N__30269));
    LocalMux I__5879 (
            .O(N__30269),
            .I(\comm_spi.n10446 ));
    InMux I__5878 (
            .O(N__30266),
            .I(n14035));
    InMux I__5877 (
            .O(N__30263),
            .I(n14036));
    InMux I__5876 (
            .O(N__30260),
            .I(N__30255));
    InMux I__5875 (
            .O(N__30259),
            .I(N__30252));
    InMux I__5874 (
            .O(N__30258),
            .I(N__30249));
    LocalMux I__5873 (
            .O(N__30255),
            .I(N__30244));
    LocalMux I__5872 (
            .O(N__30252),
            .I(N__30244));
    LocalMux I__5871 (
            .O(N__30249),
            .I(data_index_7));
    Odrv12 I__5870 (
            .O(N__30244),
            .I(data_index_7));
    InMux I__5869 (
            .O(N__30239),
            .I(n14037));
    InMux I__5868 (
            .O(N__30236),
            .I(bfn_14_17_0_));
    InMux I__5867 (
            .O(N__30233),
            .I(N__30228));
    InMux I__5866 (
            .O(N__30232),
            .I(N__30225));
    InMux I__5865 (
            .O(N__30231),
            .I(N__30222));
    LocalMux I__5864 (
            .O(N__30228),
            .I(data_index_3));
    LocalMux I__5863 (
            .O(N__30225),
            .I(data_index_3));
    LocalMux I__5862 (
            .O(N__30222),
            .I(data_index_3));
    CascadeMux I__5861 (
            .O(N__30215),
            .I(N__30209));
    CascadeMux I__5860 (
            .O(N__30214),
            .I(N__30206));
    CascadeMux I__5859 (
            .O(N__30213),
            .I(N__30203));
    InMux I__5858 (
            .O(N__30212),
            .I(N__30200));
    InMux I__5857 (
            .O(N__30209),
            .I(N__30193));
    InMux I__5856 (
            .O(N__30206),
            .I(N__30193));
    InMux I__5855 (
            .O(N__30203),
            .I(N__30193));
    LocalMux I__5854 (
            .O(N__30200),
            .I(N__30190));
    LocalMux I__5853 (
            .O(N__30193),
            .I(N__30187));
    Span4Mux_v I__5852 (
            .O(N__30190),
            .I(N__30182));
    Span4Mux_v I__5851 (
            .O(N__30187),
            .I(N__30179));
    InMux I__5850 (
            .O(N__30186),
            .I(N__30174));
    InMux I__5849 (
            .O(N__30185),
            .I(N__30174));
    Span4Mux_h I__5848 (
            .O(N__30182),
            .I(N__30171));
    Span4Mux_v I__5847 (
            .O(N__30179),
            .I(N__30168));
    LocalMux I__5846 (
            .O(N__30174),
            .I(N__30165));
    Span4Mux_h I__5845 (
            .O(N__30171),
            .I(N__30162));
    Span4Mux_h I__5844 (
            .O(N__30168),
            .I(N__30159));
    Span4Mux_h I__5843 (
            .O(N__30165),
            .I(N__30156));
    Sp12to4 I__5842 (
            .O(N__30162),
            .I(N__30151));
    Sp12to4 I__5841 (
            .O(N__30159),
            .I(N__30151));
    Span4Mux_v I__5840 (
            .O(N__30156),
            .I(N__30148));
    Odrv12 I__5839 (
            .O(N__30151),
            .I(M_DRDY2));
    Odrv4 I__5838 (
            .O(N__30148),
            .I(M_DRDY2));
    InMux I__5837 (
            .O(N__30143),
            .I(N__30140));
    LocalMux I__5836 (
            .O(N__30140),
            .I(N__30136));
    InMux I__5835 (
            .O(N__30139),
            .I(N__30133));
    Span4Mux_v I__5834 (
            .O(N__30136),
            .I(N__30130));
    LocalMux I__5833 (
            .O(N__30133),
            .I(acadc_skipcnt_14));
    Odrv4 I__5832 (
            .O(N__30130),
            .I(acadc_skipcnt_14));
    CascadeMux I__5831 (
            .O(N__30125),
            .I(N__30122));
    InMux I__5830 (
            .O(N__30122),
            .I(N__30118));
    InMux I__5829 (
            .O(N__30121),
            .I(N__30115));
    LocalMux I__5828 (
            .O(N__30118),
            .I(N__30112));
    LocalMux I__5827 (
            .O(N__30115),
            .I(acadc_skipcnt_11));
    Odrv4 I__5826 (
            .O(N__30112),
            .I(acadc_skipcnt_11));
    InMux I__5825 (
            .O(N__30107),
            .I(N__30102));
    InMux I__5824 (
            .O(N__30106),
            .I(N__30097));
    InMux I__5823 (
            .O(N__30105),
            .I(N__30097));
    LocalMux I__5822 (
            .O(N__30102),
            .I(N__30094));
    LocalMux I__5821 (
            .O(N__30097),
            .I(acadc_skipCount_11));
    Odrv12 I__5820 (
            .O(N__30094),
            .I(acadc_skipCount_11));
    CascadeMux I__5819 (
            .O(N__30089),
            .I(n23_adj_1199_cascade_));
    InMux I__5818 (
            .O(N__30086),
            .I(N__30083));
    LocalMux I__5817 (
            .O(N__30083),
            .I(n30));
    InMux I__5816 (
            .O(N__30080),
            .I(N__30077));
    LocalMux I__5815 (
            .O(N__30077),
            .I(N__30073));
    InMux I__5814 (
            .O(N__30076),
            .I(N__30070));
    Span4Mux_h I__5813 (
            .O(N__30073),
            .I(N__30067));
    LocalMux I__5812 (
            .O(N__30070),
            .I(acadc_skipcnt_10));
    Odrv4 I__5811 (
            .O(N__30067),
            .I(acadc_skipcnt_10));
    InMux I__5810 (
            .O(N__30062),
            .I(N__30059));
    LocalMux I__5809 (
            .O(N__30059),
            .I(N__30055));
    CascadeMux I__5808 (
            .O(N__30058),
            .I(N__30052));
    Span4Mux_h I__5807 (
            .O(N__30055),
            .I(N__30049));
    InMux I__5806 (
            .O(N__30052),
            .I(N__30045));
    Span4Mux_v I__5805 (
            .O(N__30049),
            .I(N__30042));
    InMux I__5804 (
            .O(N__30048),
            .I(N__30039));
    LocalMux I__5803 (
            .O(N__30045),
            .I(acadc_skipCount_12));
    Odrv4 I__5802 (
            .O(N__30042),
            .I(acadc_skipCount_12));
    LocalMux I__5801 (
            .O(N__30039),
            .I(acadc_skipCount_12));
    CascadeMux I__5800 (
            .O(N__30032),
            .I(N__30029));
    InMux I__5799 (
            .O(N__30029),
            .I(N__30025));
    InMux I__5798 (
            .O(N__30028),
            .I(N__30022));
    LocalMux I__5797 (
            .O(N__30025),
            .I(N__30019));
    LocalMux I__5796 (
            .O(N__30022),
            .I(acadc_skipcnt_12));
    Odrv4 I__5795 (
            .O(N__30019),
            .I(acadc_skipcnt_12));
    InMux I__5794 (
            .O(N__30014),
            .I(N__30011));
    LocalMux I__5793 (
            .O(N__30011),
            .I(n21));
    CascadeMux I__5792 (
            .O(N__30008),
            .I(N__30005));
    InMux I__5791 (
            .O(N__30005),
            .I(N__30000));
    InMux I__5790 (
            .O(N__30004),
            .I(N__29995));
    InMux I__5789 (
            .O(N__30003),
            .I(N__29995));
    LocalMux I__5788 (
            .O(N__30000),
            .I(N__29992));
    LocalMux I__5787 (
            .O(N__29995),
            .I(data_index_0));
    Odrv4 I__5786 (
            .O(N__29992),
            .I(data_index_0));
    InMux I__5785 (
            .O(N__29987),
            .I(N__29984));
    LocalMux I__5784 (
            .O(N__29984),
            .I(N__29981));
    Odrv4 I__5783 (
            .O(N__29981),
            .I(data_index_9_N_647_0));
    InMux I__5782 (
            .O(N__29978),
            .I(N__29973));
    InMux I__5781 (
            .O(N__29977),
            .I(N__29970));
    InMux I__5780 (
            .O(N__29976),
            .I(N__29967));
    LocalMux I__5779 (
            .O(N__29973),
            .I(data_index_1));
    LocalMux I__5778 (
            .O(N__29970),
            .I(data_index_1));
    LocalMux I__5777 (
            .O(N__29967),
            .I(data_index_1));
    InMux I__5776 (
            .O(N__29960),
            .I(N__29954));
    InMux I__5775 (
            .O(N__29959),
            .I(N__29954));
    LocalMux I__5774 (
            .O(N__29954),
            .I(n7_adj_1232));
    InMux I__5773 (
            .O(N__29951),
            .I(n14031));
    InMux I__5772 (
            .O(N__29948),
            .I(N__29943));
    InMux I__5771 (
            .O(N__29947),
            .I(N__29940));
    InMux I__5770 (
            .O(N__29946),
            .I(N__29937));
    LocalMux I__5769 (
            .O(N__29943),
            .I(N__29932));
    LocalMux I__5768 (
            .O(N__29940),
            .I(N__29932));
    LocalMux I__5767 (
            .O(N__29937),
            .I(data_index_2));
    Odrv4 I__5766 (
            .O(N__29932),
            .I(data_index_2));
    InMux I__5765 (
            .O(N__29927),
            .I(N__29921));
    InMux I__5764 (
            .O(N__29926),
            .I(N__29921));
    LocalMux I__5763 (
            .O(N__29921),
            .I(n7_adj_1230));
    InMux I__5762 (
            .O(N__29918),
            .I(n14032));
    InMux I__5761 (
            .O(N__29915),
            .I(n14033));
    InMux I__5760 (
            .O(N__29912),
            .I(N__29908));
    InMux I__5759 (
            .O(N__29911),
            .I(N__29905));
    LocalMux I__5758 (
            .O(N__29908),
            .I(N__29899));
    LocalMux I__5757 (
            .O(N__29905),
            .I(N__29899));
    InMux I__5756 (
            .O(N__29904),
            .I(N__29896));
    Span4Mux_h I__5755 (
            .O(N__29899),
            .I(N__29893));
    LocalMux I__5754 (
            .O(N__29896),
            .I(data_index_4));
    Odrv4 I__5753 (
            .O(N__29893),
            .I(data_index_4));
    InMux I__5752 (
            .O(N__29888),
            .I(N__29882));
    InMux I__5751 (
            .O(N__29887),
            .I(N__29882));
    LocalMux I__5750 (
            .O(N__29882),
            .I(N__29879));
    Odrv4 I__5749 (
            .O(N__29879),
            .I(n7_adj_1226));
    InMux I__5748 (
            .O(N__29876),
            .I(n14034));
    CascadeMux I__5747 (
            .O(N__29873),
            .I(n7_adj_1177_cascade_));
    InMux I__5746 (
            .O(N__29870),
            .I(N__29867));
    LocalMux I__5745 (
            .O(N__29867),
            .I(n8_adj_1178));
    CascadeMux I__5744 (
            .O(N__29864),
            .I(N__29861));
    CascadeBuf I__5743 (
            .O(N__29861),
            .I(N__29858));
    CascadeMux I__5742 (
            .O(N__29858),
            .I(N__29855));
    CascadeBuf I__5741 (
            .O(N__29855),
            .I(N__29852));
    CascadeMux I__5740 (
            .O(N__29852),
            .I(N__29849));
    CascadeBuf I__5739 (
            .O(N__29849),
            .I(N__29846));
    CascadeMux I__5738 (
            .O(N__29846),
            .I(N__29843));
    CascadeBuf I__5737 (
            .O(N__29843),
            .I(N__29840));
    CascadeMux I__5736 (
            .O(N__29840),
            .I(N__29837));
    CascadeBuf I__5735 (
            .O(N__29837),
            .I(N__29834));
    CascadeMux I__5734 (
            .O(N__29834),
            .I(N__29831));
    CascadeBuf I__5733 (
            .O(N__29831),
            .I(N__29828));
    CascadeMux I__5732 (
            .O(N__29828),
            .I(N__29825));
    CascadeBuf I__5731 (
            .O(N__29825),
            .I(N__29822));
    CascadeMux I__5730 (
            .O(N__29822),
            .I(N__29818));
    CascadeMux I__5729 (
            .O(N__29821),
            .I(N__29815));
    CascadeBuf I__5728 (
            .O(N__29818),
            .I(N__29812));
    CascadeBuf I__5727 (
            .O(N__29815),
            .I(N__29809));
    CascadeMux I__5726 (
            .O(N__29812),
            .I(N__29806));
    CascadeMux I__5725 (
            .O(N__29809),
            .I(N__29803));
    CascadeBuf I__5724 (
            .O(N__29806),
            .I(N__29800));
    InMux I__5723 (
            .O(N__29803),
            .I(N__29797));
    CascadeMux I__5722 (
            .O(N__29800),
            .I(N__29794));
    LocalMux I__5721 (
            .O(N__29797),
            .I(N__29791));
    InMux I__5720 (
            .O(N__29794),
            .I(N__29788));
    Span4Mux_h I__5719 (
            .O(N__29791),
            .I(N__29785));
    LocalMux I__5718 (
            .O(N__29788),
            .I(N__29782));
    Span4Mux_v I__5717 (
            .O(N__29785),
            .I(N__29779));
    Span4Mux_v I__5716 (
            .O(N__29782),
            .I(N__29776));
    Span4Mux_h I__5715 (
            .O(N__29779),
            .I(N__29773));
    Span4Mux_h I__5714 (
            .O(N__29776),
            .I(N__29770));
    Span4Mux_h I__5713 (
            .O(N__29773),
            .I(N__29767));
    Span4Mux_h I__5712 (
            .O(N__29770),
            .I(N__29764));
    Odrv4 I__5711 (
            .O(N__29767),
            .I(data_index_9_N_258_0));
    Odrv4 I__5710 (
            .O(N__29764),
            .I(data_index_9_N_258_0));
    InMux I__5709 (
            .O(N__29759),
            .I(N__29756));
    LocalMux I__5708 (
            .O(N__29756),
            .I(N__29752));
    InMux I__5707 (
            .O(N__29755),
            .I(N__29749));
    Span4Mux_h I__5706 (
            .O(N__29752),
            .I(N__29746));
    LocalMux I__5705 (
            .O(N__29749),
            .I(acadc_skipcnt_0));
    Odrv4 I__5704 (
            .O(N__29746),
            .I(acadc_skipcnt_0));
    CascadeMux I__5703 (
            .O(N__29741),
            .I(N__29738));
    InMux I__5702 (
            .O(N__29738),
            .I(N__29734));
    InMux I__5701 (
            .O(N__29737),
            .I(N__29731));
    LocalMux I__5700 (
            .O(N__29734),
            .I(N__29728));
    LocalMux I__5699 (
            .O(N__29731),
            .I(acadc_skipcnt_6));
    Odrv4 I__5698 (
            .O(N__29728),
            .I(acadc_skipcnt_6));
    InMux I__5697 (
            .O(N__29723),
            .I(N__29720));
    LocalMux I__5696 (
            .O(N__29720),
            .I(N__29717));
    Odrv4 I__5695 (
            .O(N__29717),
            .I(n18_adj_1276));
    CascadeMux I__5694 (
            .O(N__29714),
            .I(n17_adj_1277_cascade_));
    InMux I__5693 (
            .O(N__29711),
            .I(N__29705));
    InMux I__5692 (
            .O(N__29710),
            .I(N__29705));
    LocalMux I__5691 (
            .O(N__29705),
            .I(n31));
    CascadeMux I__5690 (
            .O(N__29702),
            .I(n31_cascade_));
    InMux I__5689 (
            .O(N__29699),
            .I(N__29696));
    LocalMux I__5688 (
            .O(N__29696),
            .I(n15187));
    InMux I__5687 (
            .O(N__29693),
            .I(N__29687));
    InMux I__5686 (
            .O(N__29692),
            .I(N__29687));
    LocalMux I__5685 (
            .O(N__29687),
            .I(n8_adj_1231));
    CascadeMux I__5684 (
            .O(N__29684),
            .I(N__29681));
    CascadeBuf I__5683 (
            .O(N__29681),
            .I(N__29678));
    CascadeMux I__5682 (
            .O(N__29678),
            .I(N__29675));
    CascadeBuf I__5681 (
            .O(N__29675),
            .I(N__29672));
    CascadeMux I__5680 (
            .O(N__29672),
            .I(N__29669));
    CascadeBuf I__5679 (
            .O(N__29669),
            .I(N__29666));
    CascadeMux I__5678 (
            .O(N__29666),
            .I(N__29663));
    CascadeBuf I__5677 (
            .O(N__29663),
            .I(N__29660));
    CascadeMux I__5676 (
            .O(N__29660),
            .I(N__29657));
    CascadeBuf I__5675 (
            .O(N__29657),
            .I(N__29654));
    CascadeMux I__5674 (
            .O(N__29654),
            .I(N__29651));
    CascadeBuf I__5673 (
            .O(N__29651),
            .I(N__29648));
    CascadeMux I__5672 (
            .O(N__29648),
            .I(N__29645));
    CascadeBuf I__5671 (
            .O(N__29645),
            .I(N__29642));
    CascadeMux I__5670 (
            .O(N__29642),
            .I(N__29638));
    CascadeMux I__5669 (
            .O(N__29641),
            .I(N__29635));
    CascadeBuf I__5668 (
            .O(N__29638),
            .I(N__29632));
    CascadeBuf I__5667 (
            .O(N__29635),
            .I(N__29629));
    CascadeMux I__5666 (
            .O(N__29632),
            .I(N__29626));
    CascadeMux I__5665 (
            .O(N__29629),
            .I(N__29623));
    CascadeBuf I__5664 (
            .O(N__29626),
            .I(N__29620));
    InMux I__5663 (
            .O(N__29623),
            .I(N__29617));
    CascadeMux I__5662 (
            .O(N__29620),
            .I(N__29614));
    LocalMux I__5661 (
            .O(N__29617),
            .I(N__29611));
    InMux I__5660 (
            .O(N__29614),
            .I(N__29608));
    Span4Mux_h I__5659 (
            .O(N__29611),
            .I(N__29605));
    LocalMux I__5658 (
            .O(N__29608),
            .I(N__29602));
    Sp12to4 I__5657 (
            .O(N__29605),
            .I(N__29599));
    Span4Mux_v I__5656 (
            .O(N__29602),
            .I(N__29596));
    Span12Mux_v I__5655 (
            .O(N__29599),
            .I(N__29593));
    Span4Mux_h I__5654 (
            .O(N__29596),
            .I(N__29590));
    Odrv12 I__5653 (
            .O(N__29593),
            .I(data_index_9_N_258_2));
    Odrv4 I__5652 (
            .O(N__29590),
            .I(data_index_9_N_258_2));
    IoInMux I__5651 (
            .O(N__29585),
            .I(N__29582));
    LocalMux I__5650 (
            .O(N__29582),
            .I(N__29578));
    InMux I__5649 (
            .O(N__29581),
            .I(N__29575));
    Span4Mux_s0_v I__5648 (
            .O(N__29578),
            .I(N__29572));
    LocalMux I__5647 (
            .O(N__29575),
            .I(N__29569));
    Span4Mux_v I__5646 (
            .O(N__29572),
            .I(N__29566));
    Span4Mux_v I__5645 (
            .O(N__29569),
            .I(N__29562));
    Span4Mux_v I__5644 (
            .O(N__29566),
            .I(N__29559));
    InMux I__5643 (
            .O(N__29565),
            .I(N__29556));
    Span4Mux_h I__5642 (
            .O(N__29562),
            .I(N__29553));
    Odrv4 I__5641 (
            .O(N__29559),
            .I(M_FLT1));
    LocalMux I__5640 (
            .O(N__29556),
            .I(M_FLT1));
    Odrv4 I__5639 (
            .O(N__29553),
            .I(M_FLT1));
    InMux I__5638 (
            .O(N__29546),
            .I(N__29541));
    InMux I__5637 (
            .O(N__29545),
            .I(N__29538));
    InMux I__5636 (
            .O(N__29544),
            .I(N__29535));
    LocalMux I__5635 (
            .O(N__29541),
            .I(N__29532));
    LocalMux I__5634 (
            .O(N__29538),
            .I(N__29529));
    LocalMux I__5633 (
            .O(N__29535),
            .I(buf_dds_14));
    Odrv12 I__5632 (
            .O(N__29532),
            .I(buf_dds_14));
    Odrv4 I__5631 (
            .O(N__29529),
            .I(buf_dds_14));
    InMux I__5630 (
            .O(N__29522),
            .I(N__29519));
    LocalMux I__5629 (
            .O(N__29519),
            .I(N__29516));
    Odrv4 I__5628 (
            .O(N__29516),
            .I(n4219));
    InMux I__5627 (
            .O(N__29513),
            .I(N__29508));
    InMux I__5626 (
            .O(N__29512),
            .I(N__29505));
    InMux I__5625 (
            .O(N__29511),
            .I(N__29502));
    LocalMux I__5624 (
            .O(N__29508),
            .I(N__29499));
    LocalMux I__5623 (
            .O(N__29505),
            .I(N__29496));
    LocalMux I__5622 (
            .O(N__29502),
            .I(req_data_cnt_15));
    Odrv12 I__5621 (
            .O(N__29499),
            .I(req_data_cnt_15));
    Odrv4 I__5620 (
            .O(N__29496),
            .I(req_data_cnt_15));
    InMux I__5619 (
            .O(N__29489),
            .I(N__29485));
    InMux I__5618 (
            .O(N__29488),
            .I(N__29481));
    LocalMux I__5617 (
            .O(N__29485),
            .I(N__29478));
    InMux I__5616 (
            .O(N__29484),
            .I(N__29475));
    LocalMux I__5615 (
            .O(N__29481),
            .I(req_data_cnt_9));
    Odrv4 I__5614 (
            .O(N__29478),
            .I(req_data_cnt_9));
    LocalMux I__5613 (
            .O(N__29475),
            .I(req_data_cnt_9));
    InMux I__5612 (
            .O(N__29468),
            .I(N__29465));
    LocalMux I__5611 (
            .O(N__29465),
            .I(n22));
    CascadeMux I__5610 (
            .O(N__29462),
            .I(n24_adj_1216_cascade_));
    InMux I__5609 (
            .O(N__29459),
            .I(N__29456));
    LocalMux I__5608 (
            .O(N__29456),
            .I(n30_adj_1278));
    CascadeMux I__5607 (
            .O(N__29453),
            .I(n6791_cascade_));
    CascadeMux I__5606 (
            .O(N__29450),
            .I(n8_adj_1178_cascade_));
    InMux I__5605 (
            .O(N__29447),
            .I(N__29444));
    LocalMux I__5604 (
            .O(N__29444),
            .I(n7_adj_1177));
    IoInMux I__5603 (
            .O(N__29441),
            .I(N__29438));
    LocalMux I__5602 (
            .O(N__29438),
            .I(N__29435));
    Span4Mux_s2_v I__5601 (
            .O(N__29435),
            .I(N__29432));
    Span4Mux_h I__5600 (
            .O(N__29432),
            .I(N__29429));
    Sp12to4 I__5599 (
            .O(N__29429),
            .I(N__29425));
    InMux I__5598 (
            .O(N__29428),
            .I(N__29421));
    Span12Mux_v I__5597 (
            .O(N__29425),
            .I(N__29418));
    InMux I__5596 (
            .O(N__29424),
            .I(N__29415));
    LocalMux I__5595 (
            .O(N__29421),
            .I(N__29412));
    Odrv12 I__5594 (
            .O(N__29418),
            .I(M_OSR1));
    LocalMux I__5593 (
            .O(N__29415),
            .I(M_OSR1));
    Odrv4 I__5592 (
            .O(N__29412),
            .I(M_OSR1));
    InMux I__5591 (
            .O(N__29405),
            .I(N__29402));
    LocalMux I__5590 (
            .O(N__29402),
            .I(N__29399));
    Odrv4 I__5589 (
            .O(N__29399),
            .I(n15479));
    CascadeMux I__5588 (
            .O(N__29396),
            .I(N__29393));
    InMux I__5587 (
            .O(N__29393),
            .I(N__29390));
    LocalMux I__5586 (
            .O(N__29390),
            .I(N__29387));
    Span4Mux_h I__5585 (
            .O(N__29387),
            .I(N__29383));
    InMux I__5584 (
            .O(N__29386),
            .I(N__29380));
    Odrv4 I__5583 (
            .O(N__29383),
            .I(cmd_rdadctmp_31_adj_1081));
    LocalMux I__5582 (
            .O(N__29380),
            .I(cmd_rdadctmp_31_adj_1081));
    CascadeMux I__5581 (
            .O(N__29375),
            .I(n8_adj_1221_cascade_));
    CascadeMux I__5580 (
            .O(N__29372),
            .I(N__29369));
    InMux I__5579 (
            .O(N__29369),
            .I(N__29366));
    LocalMux I__5578 (
            .O(N__29366),
            .I(N__29363));
    Odrv4 I__5577 (
            .O(N__29363),
            .I(n4205));
    InMux I__5576 (
            .O(N__29360),
            .I(N__29357));
    LocalMux I__5575 (
            .O(N__29357),
            .I(N__29353));
    InMux I__5574 (
            .O(N__29356),
            .I(N__29350));
    Span4Mux_v I__5573 (
            .O(N__29353),
            .I(N__29347));
    LocalMux I__5572 (
            .O(N__29350),
            .I(buf_device_acadc_7));
    Odrv4 I__5571 (
            .O(N__29347),
            .I(buf_device_acadc_7));
    CascadeMux I__5570 (
            .O(N__29342),
            .I(n4260_cascade_));
    InMux I__5569 (
            .O(N__29339),
            .I(N__29336));
    LocalMux I__5568 (
            .O(N__29336),
            .I(N__29333));
    Span4Mux_h I__5567 (
            .O(N__29333),
            .I(N__29330));
    Odrv4 I__5566 (
            .O(N__29330),
            .I(n15402));
    InMux I__5565 (
            .O(N__29327),
            .I(N__29324));
    LocalMux I__5564 (
            .O(N__29324),
            .I(N__29321));
    Span4Mux_v I__5563 (
            .O(N__29321),
            .I(N__29318));
    Span4Mux_v I__5562 (
            .O(N__29318),
            .I(N__29315));
    Span4Mux_v I__5561 (
            .O(N__29315),
            .I(N__29312));
    Sp12to4 I__5560 (
            .O(N__29312),
            .I(N__29309));
    Span12Mux_h I__5559 (
            .O(N__29309),
            .I(N__29306));
    Odrv12 I__5558 (
            .O(N__29306),
            .I(ICE_CHKCABLE));
    CascadeMux I__5557 (
            .O(N__29303),
            .I(n90_adj_1154_cascade_));
    InMux I__5556 (
            .O(N__29300),
            .I(N__29297));
    LocalMux I__5555 (
            .O(N__29297),
            .I(N__29294));
    Span4Mux_h I__5554 (
            .O(N__29294),
            .I(N__29291));
    Span4Mux_h I__5553 (
            .O(N__29291),
            .I(N__29288));
    Odrv4 I__5552 (
            .O(N__29288),
            .I(n72));
    CascadeMux I__5551 (
            .O(N__29285),
            .I(N__29282));
    InMux I__5550 (
            .O(N__29282),
            .I(N__29279));
    LocalMux I__5549 (
            .O(N__29279),
            .I(\CLOCK_DDS.tmp_buf_10 ));
    InMux I__5548 (
            .O(N__29276),
            .I(N__29273));
    LocalMux I__5547 (
            .O(N__29273),
            .I(\CLOCK_DDS.tmp_buf_11 ));
    CascadeMux I__5546 (
            .O(N__29270),
            .I(N__29267));
    InMux I__5545 (
            .O(N__29267),
            .I(N__29264));
    LocalMux I__5544 (
            .O(N__29264),
            .I(N__29261));
    Odrv4 I__5543 (
            .O(N__29261),
            .I(\CLOCK_DDS.tmp_buf_12 ));
    CascadeMux I__5542 (
            .O(N__29258),
            .I(N__29255));
    InMux I__5541 (
            .O(N__29255),
            .I(N__29252));
    LocalMux I__5540 (
            .O(N__29252),
            .I(\CLOCK_DDS.tmp_buf_13 ));
    InMux I__5539 (
            .O(N__29249),
            .I(N__29246));
    LocalMux I__5538 (
            .O(N__29246),
            .I(\CLOCK_DDS.tmp_buf_14 ));
    InMux I__5537 (
            .O(N__29243),
            .I(N__29240));
    LocalMux I__5536 (
            .O(N__29240),
            .I(N__29236));
    InMux I__5535 (
            .O(N__29239),
            .I(N__29233));
    Span4Mux_v I__5534 (
            .O(N__29236),
            .I(N__29228));
    LocalMux I__5533 (
            .O(N__29233),
            .I(N__29228));
    Span4Mux_h I__5532 (
            .O(N__29228),
            .I(N__29224));
    InMux I__5531 (
            .O(N__29227),
            .I(N__29221));
    Sp12to4 I__5530 (
            .O(N__29224),
            .I(N__29218));
    LocalMux I__5529 (
            .O(N__29221),
            .I(buf_dds_9));
    Odrv12 I__5528 (
            .O(N__29218),
            .I(buf_dds_9));
    CascadeMux I__5527 (
            .O(N__29213),
            .I(N__29210));
    InMux I__5526 (
            .O(N__29210),
            .I(N__29207));
    LocalMux I__5525 (
            .O(N__29207),
            .I(\CLOCK_DDS.tmp_buf_9 ));
    InMux I__5524 (
            .O(N__29204),
            .I(N__29201));
    LocalMux I__5523 (
            .O(N__29201),
            .I(\CLOCK_DDS.tmp_buf_8 ));
    InMux I__5522 (
            .O(N__29198),
            .I(N__29195));
    LocalMux I__5521 (
            .O(N__29195),
            .I(N__29192));
    Span4Mux_h I__5520 (
            .O(N__29192),
            .I(N__29189));
    Span4Mux_v I__5519 (
            .O(N__29189),
            .I(N__29186));
    Odrv4 I__5518 (
            .O(N__29186),
            .I(n15474));
    InMux I__5517 (
            .O(N__29183),
            .I(N__29180));
    LocalMux I__5516 (
            .O(N__29180),
            .I(N__29177));
    Span4Mux_h I__5515 (
            .O(N__29177),
            .I(N__29174));
    Span4Mux_v I__5514 (
            .O(N__29174),
            .I(N__29171));
    Odrv4 I__5513 (
            .O(N__29171),
            .I(n15478));
    InMux I__5512 (
            .O(N__29168),
            .I(N__29165));
    LocalMux I__5511 (
            .O(N__29165),
            .I(N__29162));
    Span4Mux_v I__5510 (
            .O(N__29162),
            .I(N__29159));
    Odrv4 I__5509 (
            .O(N__29159),
            .I(n15680));
    InMux I__5508 (
            .O(N__29156),
            .I(N__29153));
    LocalMux I__5507 (
            .O(N__29153),
            .I(N__29149));
    InMux I__5506 (
            .O(N__29152),
            .I(N__29146));
    Span12Mux_v I__5505 (
            .O(N__29149),
            .I(N__29143));
    LocalMux I__5504 (
            .O(N__29146),
            .I(N__29140));
    Odrv12 I__5503 (
            .O(N__29143),
            .I(\comm_spi.n10449 ));
    Odrv4 I__5502 (
            .O(N__29140),
            .I(\comm_spi.n10449 ));
    InMux I__5501 (
            .O(N__29135),
            .I(N__29132));
    LocalMux I__5500 (
            .O(N__29132),
            .I(N__29129));
    Span4Mux_h I__5499 (
            .O(N__29129),
            .I(N__29125));
    InMux I__5498 (
            .O(N__29128),
            .I(N__29122));
    Odrv4 I__5497 (
            .O(N__29125),
            .I(\comm_spi.n10448 ));
    LocalMux I__5496 (
            .O(N__29122),
            .I(\comm_spi.n10448 ));
    InMux I__5495 (
            .O(N__29117),
            .I(N__29114));
    LocalMux I__5494 (
            .O(N__29114),
            .I(N__29111));
    Span4Mux_h I__5493 (
            .O(N__29111),
            .I(N__29108));
    Span4Mux_h I__5492 (
            .O(N__29108),
            .I(N__29105));
    Odrv4 I__5491 (
            .O(N__29105),
            .I(n15387));
    InMux I__5490 (
            .O(N__29102),
            .I(N__29099));
    LocalMux I__5489 (
            .O(N__29099),
            .I(N__29096));
    Span4Mux_v I__5488 (
            .O(N__29096),
            .I(N__29093));
    Span4Mux_h I__5487 (
            .O(N__29093),
            .I(N__29090));
    Odrv4 I__5486 (
            .O(N__29090),
            .I(n15390));
    InMux I__5485 (
            .O(N__29087),
            .I(N__29084));
    LocalMux I__5484 (
            .O(N__29084),
            .I(N__29081));
    Odrv12 I__5483 (
            .O(N__29081),
            .I(buf_data2_22));
    InMux I__5482 (
            .O(N__29078),
            .I(N__29075));
    LocalMux I__5481 (
            .O(N__29075),
            .I(N__29071));
    CascadeMux I__5480 (
            .O(N__29074),
            .I(N__29068));
    Span4Mux_h I__5479 (
            .O(N__29071),
            .I(N__29065));
    InMux I__5478 (
            .O(N__29068),
            .I(N__29062));
    Span4Mux_h I__5477 (
            .O(N__29065),
            .I(N__29056));
    LocalMux I__5476 (
            .O(N__29062),
            .I(N__29056));
    InMux I__5475 (
            .O(N__29061),
            .I(N__29053));
    Span4Mux_h I__5474 (
            .O(N__29056),
            .I(N__29050));
    LocalMux I__5473 (
            .O(N__29053),
            .I(buf_adcdata4_22));
    Odrv4 I__5472 (
            .O(N__29050),
            .I(buf_adcdata4_22));
    InMux I__5471 (
            .O(N__29045),
            .I(N__29042));
    LocalMux I__5470 (
            .O(N__29042),
            .I(N__29039));
    Span4Mux_v I__5469 (
            .O(N__29039),
            .I(N__29036));
    Span4Mux_h I__5468 (
            .O(N__29036),
            .I(N__29033));
    Odrv4 I__5467 (
            .O(N__29033),
            .I(n4102));
    InMux I__5466 (
            .O(N__29030),
            .I(N__29025));
    InMux I__5465 (
            .O(N__29029),
            .I(N__29022));
    InMux I__5464 (
            .O(N__29028),
            .I(N__29019));
    LocalMux I__5463 (
            .O(N__29025),
            .I(\comm_spi.n16902 ));
    LocalMux I__5462 (
            .O(N__29022),
            .I(\comm_spi.n16902 ));
    LocalMux I__5461 (
            .O(N__29019),
            .I(\comm_spi.n16902 ));
    InMux I__5460 (
            .O(N__29012),
            .I(N__29009));
    LocalMux I__5459 (
            .O(N__29009),
            .I(N__29006));
    Span4Mux_v I__5458 (
            .O(N__29006),
            .I(N__29002));
    InMux I__5457 (
            .O(N__29005),
            .I(N__28999));
    Odrv4 I__5456 (
            .O(N__29002),
            .I(\comm_spi.n10476 ));
    LocalMux I__5455 (
            .O(N__28999),
            .I(\comm_spi.n10476 ));
    InMux I__5454 (
            .O(N__28994),
            .I(N__28991));
    LocalMux I__5453 (
            .O(N__28991),
            .I(N__28988));
    Span4Mux_v I__5452 (
            .O(N__28988),
            .I(N__28985));
    Span4Mux_h I__5451 (
            .O(N__28985),
            .I(N__28981));
    InMux I__5450 (
            .O(N__28984),
            .I(N__28978));
    Odrv4 I__5449 (
            .O(N__28981),
            .I(\comm_spi.n10480 ));
    LocalMux I__5448 (
            .O(N__28978),
            .I(\comm_spi.n10480 ));
    SRMux I__5447 (
            .O(N__28973),
            .I(N__28970));
    LocalMux I__5446 (
            .O(N__28970),
            .I(\comm_spi.data_tx_7__N_816 ));
    InMux I__5445 (
            .O(N__28967),
            .I(N__28964));
    LocalMux I__5444 (
            .O(N__28964),
            .I(N__28960));
    InMux I__5443 (
            .O(N__28963),
            .I(N__28957));
    Span4Mux_v I__5442 (
            .O(N__28960),
            .I(N__28954));
    LocalMux I__5441 (
            .O(N__28957),
            .I(\comm_spi.n10472 ));
    Odrv4 I__5440 (
            .O(N__28954),
            .I(\comm_spi.n10472 ));
    InMux I__5439 (
            .O(N__28949),
            .I(N__28946));
    LocalMux I__5438 (
            .O(N__28946),
            .I(N__28942));
    InMux I__5437 (
            .O(N__28945),
            .I(N__28939));
    Odrv4 I__5436 (
            .O(N__28942),
            .I(\comm_spi.n10471 ));
    LocalMux I__5435 (
            .O(N__28939),
            .I(\comm_spi.n10471 ));
    InMux I__5434 (
            .O(N__28934),
            .I(N__28931));
    LocalMux I__5433 (
            .O(N__28931),
            .I(N__28928));
    Span4Mux_v I__5432 (
            .O(N__28928),
            .I(N__28924));
    InMux I__5431 (
            .O(N__28927),
            .I(N__28921));
    Odrv4 I__5430 (
            .O(N__28924),
            .I(\comm_spi.n10475 ));
    LocalMux I__5429 (
            .O(N__28921),
            .I(\comm_spi.n10475 ));
    SRMux I__5428 (
            .O(N__28916),
            .I(N__28913));
    LocalMux I__5427 (
            .O(N__28913),
            .I(N__28910));
    Odrv4 I__5426 (
            .O(N__28910),
            .I(\comm_spi.data_tx_7__N_807 ));
    InMux I__5425 (
            .O(N__28907),
            .I(N__28904));
    LocalMux I__5424 (
            .O(N__28904),
            .I(N__28901));
    Span4Mux_v I__5423 (
            .O(N__28901),
            .I(N__28898));
    Span4Mux_h I__5422 (
            .O(N__28898),
            .I(N__28893));
    InMux I__5421 (
            .O(N__28897),
            .I(N__28890));
    InMux I__5420 (
            .O(N__28896),
            .I(N__28887));
    Odrv4 I__5419 (
            .O(N__28893),
            .I(\comm_spi.n16896 ));
    LocalMux I__5418 (
            .O(N__28890),
            .I(\comm_spi.n16896 ));
    LocalMux I__5417 (
            .O(N__28887),
            .I(\comm_spi.n16896 ));
    InMux I__5416 (
            .O(N__28880),
            .I(n13972));
    InMux I__5415 (
            .O(N__28877),
            .I(n13973));
    InMux I__5414 (
            .O(N__28874),
            .I(bfn_13_18_0_));
    InMux I__5413 (
            .O(N__28871),
            .I(n13975));
    InMux I__5412 (
            .O(N__28868),
            .I(n13976));
    InMux I__5411 (
            .O(N__28865),
            .I(n13977));
    InMux I__5410 (
            .O(N__28862),
            .I(n13978));
    InMux I__5409 (
            .O(N__28859),
            .I(n13979));
    InMux I__5408 (
            .O(N__28856),
            .I(n13980));
    SRMux I__5407 (
            .O(N__28853),
            .I(N__28850));
    LocalMux I__5406 (
            .O(N__28850),
            .I(N__28845));
    SRMux I__5405 (
            .O(N__28849),
            .I(N__28842));
    SRMux I__5404 (
            .O(N__28848),
            .I(N__28839));
    Span4Mux_v I__5403 (
            .O(N__28845),
            .I(N__28830));
    LocalMux I__5402 (
            .O(N__28842),
            .I(N__28830));
    LocalMux I__5401 (
            .O(N__28839),
            .I(N__28830));
    SRMux I__5400 (
            .O(N__28838),
            .I(N__28827));
    SRMux I__5399 (
            .O(N__28837),
            .I(N__28824));
    Span4Mux_v I__5398 (
            .O(N__28830),
            .I(N__28814));
    LocalMux I__5397 (
            .O(N__28827),
            .I(N__28814));
    LocalMux I__5396 (
            .O(N__28824),
            .I(N__28814));
    SRMux I__5395 (
            .O(N__28823),
            .I(N__28811));
    SRMux I__5394 (
            .O(N__28822),
            .I(N__28808));
    SRMux I__5393 (
            .O(N__28821),
            .I(N__28803));
    Span4Mux_v I__5392 (
            .O(N__28814),
            .I(N__28795));
    LocalMux I__5391 (
            .O(N__28811),
            .I(N__28795));
    LocalMux I__5390 (
            .O(N__28808),
            .I(N__28795));
    SRMux I__5389 (
            .O(N__28807),
            .I(N__28792));
    SRMux I__5388 (
            .O(N__28806),
            .I(N__28789));
    LocalMux I__5387 (
            .O(N__28803),
            .I(N__28786));
    SRMux I__5386 (
            .O(N__28802),
            .I(N__28783));
    Span4Mux_v I__5385 (
            .O(N__28795),
            .I(N__28775));
    LocalMux I__5384 (
            .O(N__28792),
            .I(N__28775));
    LocalMux I__5383 (
            .O(N__28789),
            .I(N__28775));
    Span4Mux_v I__5382 (
            .O(N__28786),
            .I(N__28762));
    LocalMux I__5381 (
            .O(N__28783),
            .I(N__28762));
    IoInMux I__5380 (
            .O(N__28782),
            .I(N__28759));
    Span4Mux_v I__5379 (
            .O(N__28775),
            .I(N__28756));
    SRMux I__5378 (
            .O(N__28774),
            .I(N__28753));
    InMux I__5377 (
            .O(N__28773),
            .I(N__28744));
    InMux I__5376 (
            .O(N__28772),
            .I(N__28744));
    InMux I__5375 (
            .O(N__28771),
            .I(N__28744));
    InMux I__5374 (
            .O(N__28770),
            .I(N__28735));
    InMux I__5373 (
            .O(N__28769),
            .I(N__28735));
    InMux I__5372 (
            .O(N__28768),
            .I(N__28735));
    InMux I__5371 (
            .O(N__28767),
            .I(N__28735));
    Span4Mux_h I__5370 (
            .O(N__28762),
            .I(N__28732));
    LocalMux I__5369 (
            .O(N__28759),
            .I(N__28729));
    Span4Mux_h I__5368 (
            .O(N__28756),
            .I(N__28724));
    LocalMux I__5367 (
            .O(N__28753),
            .I(N__28724));
    InMux I__5366 (
            .O(N__28752),
            .I(N__28721));
    InMux I__5365 (
            .O(N__28751),
            .I(N__28718));
    LocalMux I__5364 (
            .O(N__28744),
            .I(N__28713));
    LocalMux I__5363 (
            .O(N__28735),
            .I(N__28713));
    Span4Mux_h I__5362 (
            .O(N__28732),
            .I(N__28710));
    Span4Mux_s2_v I__5361 (
            .O(N__28729),
            .I(N__28707));
    Span4Mux_h I__5360 (
            .O(N__28724),
            .I(N__28704));
    LocalMux I__5359 (
            .O(N__28721),
            .I(N__28699));
    LocalMux I__5358 (
            .O(N__28718),
            .I(N__28699));
    Span12Mux_v I__5357 (
            .O(N__28713),
            .I(N__28696));
    Span4Mux_v I__5356 (
            .O(N__28710),
            .I(N__28691));
    Span4Mux_v I__5355 (
            .O(N__28707),
            .I(N__28691));
    Span4Mux_h I__5354 (
            .O(N__28704),
            .I(N__28686));
    Span4Mux_v I__5353 (
            .O(N__28699),
            .I(N__28686));
    Odrv12 I__5352 (
            .O(N__28696),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5351 (
            .O(N__28691),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5350 (
            .O(N__28686),
            .I(CONSTANT_ONE_NET));
    InMux I__5349 (
            .O(N__28679),
            .I(N__28675));
    InMux I__5348 (
            .O(N__28678),
            .I(N__28672));
    LocalMux I__5347 (
            .O(N__28675),
            .I(N__28669));
    LocalMux I__5346 (
            .O(N__28672),
            .I(acadc_skipcnt_1));
    Odrv4 I__5345 (
            .O(N__28669),
            .I(acadc_skipcnt_1));
    InMux I__5344 (
            .O(N__28664),
            .I(bfn_13_17_0_));
    InMux I__5343 (
            .O(N__28661),
            .I(n13967));
    InMux I__5342 (
            .O(N__28658),
            .I(n13968));
    CascadeMux I__5341 (
            .O(N__28655),
            .I(N__28652));
    InMux I__5340 (
            .O(N__28652),
            .I(N__28648));
    InMux I__5339 (
            .O(N__28651),
            .I(N__28645));
    LocalMux I__5338 (
            .O(N__28648),
            .I(N__28642));
    LocalMux I__5337 (
            .O(N__28645),
            .I(acadc_skipcnt_4));
    Odrv4 I__5336 (
            .O(N__28642),
            .I(acadc_skipcnt_4));
    InMux I__5335 (
            .O(N__28637),
            .I(n13969));
    InMux I__5334 (
            .O(N__28634),
            .I(n13970));
    InMux I__5333 (
            .O(N__28631),
            .I(n13971));
    InMux I__5332 (
            .O(N__28628),
            .I(N__28625));
    LocalMux I__5331 (
            .O(N__28625),
            .I(N__28622));
    Span12Mux_h I__5330 (
            .O(N__28622),
            .I(N__28619));
    Odrv12 I__5329 (
            .O(N__28619),
            .I(buf_data2_13));
    InMux I__5328 (
            .O(N__28616),
            .I(N__28611));
    InMux I__5327 (
            .O(N__28615),
            .I(N__28608));
    InMux I__5326 (
            .O(N__28614),
            .I(N__28605));
    LocalMux I__5325 (
            .O(N__28611),
            .I(N__28598));
    LocalMux I__5324 (
            .O(N__28608),
            .I(N__28598));
    LocalMux I__5323 (
            .O(N__28605),
            .I(N__28598));
    Odrv12 I__5322 (
            .O(N__28598),
            .I(buf_adcdata4_13));
    InMux I__5321 (
            .O(N__28595),
            .I(N__28592));
    LocalMux I__5320 (
            .O(N__28592),
            .I(N__28589));
    Span4Mux_v I__5319 (
            .O(N__28589),
            .I(N__28586));
    Span4Mux_h I__5318 (
            .O(N__28586),
            .I(N__28583));
    Span4Mux_h I__5317 (
            .O(N__28583),
            .I(N__28580));
    Odrv4 I__5316 (
            .O(N__28580),
            .I(n4059));
    InMux I__5315 (
            .O(N__28577),
            .I(N__28574));
    LocalMux I__5314 (
            .O(N__28574),
            .I(n8_adj_1233));
    CascadeMux I__5313 (
            .O(N__28571),
            .I(n8_adj_1233_cascade_));
    IoInMux I__5312 (
            .O(N__28568),
            .I(N__28565));
    LocalMux I__5311 (
            .O(N__28565),
            .I(N__28562));
    Span4Mux_s3_v I__5310 (
            .O(N__28562),
            .I(N__28559));
    Span4Mux_v I__5309 (
            .O(N__28559),
            .I(N__28555));
    CascadeMux I__5308 (
            .O(N__28558),
            .I(N__28551));
    Span4Mux_v I__5307 (
            .O(N__28555),
            .I(N__28548));
    InMux I__5306 (
            .O(N__28554),
            .I(N__28545));
    InMux I__5305 (
            .O(N__28551),
            .I(N__28542));
    Odrv4 I__5304 (
            .O(N__28548),
            .I(M_FLT0));
    LocalMux I__5303 (
            .O(N__28545),
            .I(M_FLT0));
    LocalMux I__5302 (
            .O(N__28542),
            .I(M_FLT0));
    InMux I__5301 (
            .O(N__28535),
            .I(N__28532));
    LocalMux I__5300 (
            .O(N__28532),
            .I(N__28529));
    Odrv12 I__5299 (
            .O(N__28529),
            .I(n66_adj_1166));
    InMux I__5298 (
            .O(N__28526),
            .I(bfn_13_16_0_));
    InMux I__5297 (
            .O(N__28523),
            .I(N__28519));
    InMux I__5296 (
            .O(N__28522),
            .I(N__28516));
    LocalMux I__5295 (
            .O(N__28519),
            .I(eis_end_N_773));
    LocalMux I__5294 (
            .O(N__28516),
            .I(eis_end_N_773));
    CascadeMux I__5293 (
            .O(N__28511),
            .I(eis_end_N_773_cascade_));
    InMux I__5292 (
            .O(N__28508),
            .I(N__28505));
    LocalMux I__5291 (
            .O(N__28505),
            .I(n15510));
    InMux I__5290 (
            .O(N__28502),
            .I(N__28496));
    InMux I__5289 (
            .O(N__28501),
            .I(N__28496));
    LocalMux I__5288 (
            .O(N__28496),
            .I(n8_adj_1227));
    CascadeMux I__5287 (
            .O(N__28493),
            .I(N__28490));
    InMux I__5286 (
            .O(N__28490),
            .I(N__28484));
    InMux I__5285 (
            .O(N__28489),
            .I(N__28484));
    LocalMux I__5284 (
            .O(N__28484),
            .I(N__28480));
    CascadeMux I__5283 (
            .O(N__28483),
            .I(N__28477));
    Span4Mux_h I__5282 (
            .O(N__28480),
            .I(N__28474));
    InMux I__5281 (
            .O(N__28477),
            .I(N__28471));
    Odrv4 I__5280 (
            .O(N__28474),
            .I(cmd_rdadctmp_24_adj_1088));
    LocalMux I__5279 (
            .O(N__28471),
            .I(cmd_rdadctmp_24_adj_1088));
    CascadeMux I__5278 (
            .O(N__28466),
            .I(N__28463));
    CascadeBuf I__5277 (
            .O(N__28463),
            .I(N__28460));
    CascadeMux I__5276 (
            .O(N__28460),
            .I(N__28457));
    CascadeBuf I__5275 (
            .O(N__28457),
            .I(N__28454));
    CascadeMux I__5274 (
            .O(N__28454),
            .I(N__28451));
    CascadeBuf I__5273 (
            .O(N__28451),
            .I(N__28448));
    CascadeMux I__5272 (
            .O(N__28448),
            .I(N__28445));
    CascadeBuf I__5271 (
            .O(N__28445),
            .I(N__28442));
    CascadeMux I__5270 (
            .O(N__28442),
            .I(N__28439));
    CascadeBuf I__5269 (
            .O(N__28439),
            .I(N__28436));
    CascadeMux I__5268 (
            .O(N__28436),
            .I(N__28433));
    CascadeBuf I__5267 (
            .O(N__28433),
            .I(N__28430));
    CascadeMux I__5266 (
            .O(N__28430),
            .I(N__28427));
    CascadeBuf I__5265 (
            .O(N__28427),
            .I(N__28423));
    CascadeMux I__5264 (
            .O(N__28426),
            .I(N__28420));
    CascadeMux I__5263 (
            .O(N__28423),
            .I(N__28417));
    CascadeBuf I__5262 (
            .O(N__28420),
            .I(N__28414));
    CascadeBuf I__5261 (
            .O(N__28417),
            .I(N__28411));
    CascadeMux I__5260 (
            .O(N__28414),
            .I(N__28408));
    CascadeMux I__5259 (
            .O(N__28411),
            .I(N__28405));
    InMux I__5258 (
            .O(N__28408),
            .I(N__28402));
    CascadeBuf I__5257 (
            .O(N__28405),
            .I(N__28399));
    LocalMux I__5256 (
            .O(N__28402),
            .I(N__28396));
    CascadeMux I__5255 (
            .O(N__28399),
            .I(N__28393));
    Span4Mux_h I__5254 (
            .O(N__28396),
            .I(N__28390));
    InMux I__5253 (
            .O(N__28393),
            .I(N__28387));
    Span4Mux_v I__5252 (
            .O(N__28390),
            .I(N__28384));
    LocalMux I__5251 (
            .O(N__28387),
            .I(N__28381));
    Span4Mux_h I__5250 (
            .O(N__28384),
            .I(N__28378));
    Span4Mux_v I__5249 (
            .O(N__28381),
            .I(N__28375));
    Span4Mux_h I__5248 (
            .O(N__28378),
            .I(N__28372));
    Span4Mux_h I__5247 (
            .O(N__28375),
            .I(N__28369));
    Odrv4 I__5246 (
            .O(N__28372),
            .I(data_index_9_N_258_1));
    Odrv4 I__5245 (
            .O(N__28369),
            .I(data_index_9_N_258_1));
    SRMux I__5244 (
            .O(N__28364),
            .I(N__28360));
    SRMux I__5243 (
            .O(N__28363),
            .I(N__28355));
    LocalMux I__5242 (
            .O(N__28360),
            .I(N__28350));
    SRMux I__5241 (
            .O(N__28359),
            .I(N__28347));
    SRMux I__5240 (
            .O(N__28358),
            .I(N__28341));
    LocalMux I__5239 (
            .O(N__28355),
            .I(N__28337));
    SRMux I__5238 (
            .O(N__28354),
            .I(N__28334));
    SRMux I__5237 (
            .O(N__28353),
            .I(N__28331));
    Span4Mux_v I__5236 (
            .O(N__28350),
            .I(N__28326));
    LocalMux I__5235 (
            .O(N__28347),
            .I(N__28326));
    SRMux I__5234 (
            .O(N__28346),
            .I(N__28323));
    SRMux I__5233 (
            .O(N__28345),
            .I(N__28319));
    SRMux I__5232 (
            .O(N__28344),
            .I(N__28316));
    LocalMux I__5231 (
            .O(N__28341),
            .I(N__28313));
    SRMux I__5230 (
            .O(N__28340),
            .I(N__28310));
    Span4Mux_h I__5229 (
            .O(N__28337),
            .I(N__28305));
    LocalMux I__5228 (
            .O(N__28334),
            .I(N__28305));
    LocalMux I__5227 (
            .O(N__28331),
            .I(N__28302));
    Span4Mux_v I__5226 (
            .O(N__28326),
            .I(N__28297));
    LocalMux I__5225 (
            .O(N__28323),
            .I(N__28297));
    SRMux I__5224 (
            .O(N__28322),
            .I(N__28294));
    LocalMux I__5223 (
            .O(N__28319),
            .I(N__28291));
    LocalMux I__5222 (
            .O(N__28316),
            .I(N__28288));
    Span4Mux_h I__5221 (
            .O(N__28313),
            .I(N__28285));
    LocalMux I__5220 (
            .O(N__28310),
            .I(N__28282));
    Span4Mux_v I__5219 (
            .O(N__28305),
            .I(N__28273));
    Span4Mux_h I__5218 (
            .O(N__28302),
            .I(N__28273));
    Span4Mux_v I__5217 (
            .O(N__28297),
            .I(N__28273));
    LocalMux I__5216 (
            .O(N__28294),
            .I(N__28273));
    Span4Mux_v I__5215 (
            .O(N__28291),
            .I(N__28269));
    Span4Mux_h I__5214 (
            .O(N__28288),
            .I(N__28266));
    Span4Mux_v I__5213 (
            .O(N__28285),
            .I(N__28261));
    Span4Mux_h I__5212 (
            .O(N__28282),
            .I(N__28261));
    Span4Mux_v I__5211 (
            .O(N__28273),
            .I(N__28258));
    SRMux I__5210 (
            .O(N__28272),
            .I(N__28255));
    Span4Mux_h I__5209 (
            .O(N__28269),
            .I(N__28252));
    Span4Mux_v I__5208 (
            .O(N__28266),
            .I(N__28249));
    Span4Mux_v I__5207 (
            .O(N__28261),
            .I(N__28242));
    Span4Mux_h I__5206 (
            .O(N__28258),
            .I(N__28242));
    LocalMux I__5205 (
            .O(N__28255),
            .I(N__28242));
    Span4Mux_h I__5204 (
            .O(N__28252),
            .I(N__28239));
    Span4Mux_h I__5203 (
            .O(N__28249),
            .I(N__28236));
    Sp12to4 I__5202 (
            .O(N__28242),
            .I(N__28233));
    Odrv4 I__5201 (
            .O(N__28239),
            .I(raw_buf1_N_775));
    Odrv4 I__5200 (
            .O(N__28236),
            .I(raw_buf1_N_775));
    Odrv12 I__5199 (
            .O(N__28233),
            .I(raw_buf1_N_775));
    InMux I__5198 (
            .O(N__28226),
            .I(N__28222));
    InMux I__5197 (
            .O(N__28225),
            .I(N__28219));
    LocalMux I__5196 (
            .O(N__28222),
            .I(N__28214));
    LocalMux I__5195 (
            .O(N__28219),
            .I(N__28214));
    Span4Mux_h I__5194 (
            .O(N__28214),
            .I(N__28211));
    Odrv4 I__5193 (
            .O(N__28211),
            .I(n14087));
    CascadeMux I__5192 (
            .O(N__28208),
            .I(n15356_cascade_));
    CascadeMux I__5191 (
            .O(N__28205),
            .I(n15695_cascade_));
    InMux I__5190 (
            .O(N__28202),
            .I(N__28199));
    LocalMux I__5189 (
            .O(N__28199),
            .I(n15696));
    CascadeMux I__5188 (
            .O(N__28196),
            .I(n15700_cascade_));
    InMux I__5187 (
            .O(N__28193),
            .I(N__28190));
    LocalMux I__5186 (
            .O(N__28190),
            .I(n3));
    CEMux I__5185 (
            .O(N__28187),
            .I(N__28184));
    LocalMux I__5184 (
            .O(N__28184),
            .I(n8459));
    CascadeMux I__5183 (
            .O(N__28181),
            .I(N__28178));
    CascadeBuf I__5182 (
            .O(N__28178),
            .I(N__28175));
    CascadeMux I__5181 (
            .O(N__28175),
            .I(N__28172));
    CascadeBuf I__5180 (
            .O(N__28172),
            .I(N__28169));
    CascadeMux I__5179 (
            .O(N__28169),
            .I(N__28166));
    CascadeBuf I__5178 (
            .O(N__28166),
            .I(N__28163));
    CascadeMux I__5177 (
            .O(N__28163),
            .I(N__28160));
    CascadeBuf I__5176 (
            .O(N__28160),
            .I(N__28157));
    CascadeMux I__5175 (
            .O(N__28157),
            .I(N__28154));
    CascadeBuf I__5174 (
            .O(N__28154),
            .I(N__28151));
    CascadeMux I__5173 (
            .O(N__28151),
            .I(N__28148));
    CascadeBuf I__5172 (
            .O(N__28148),
            .I(N__28145));
    CascadeMux I__5171 (
            .O(N__28145),
            .I(N__28142));
    CascadeBuf I__5170 (
            .O(N__28142),
            .I(N__28138));
    CascadeMux I__5169 (
            .O(N__28141),
            .I(N__28135));
    CascadeMux I__5168 (
            .O(N__28138),
            .I(N__28132));
    CascadeBuf I__5167 (
            .O(N__28135),
            .I(N__28129));
    CascadeBuf I__5166 (
            .O(N__28132),
            .I(N__28126));
    CascadeMux I__5165 (
            .O(N__28129),
            .I(N__28123));
    CascadeMux I__5164 (
            .O(N__28126),
            .I(N__28120));
    InMux I__5163 (
            .O(N__28123),
            .I(N__28117));
    CascadeBuf I__5162 (
            .O(N__28120),
            .I(N__28114));
    LocalMux I__5161 (
            .O(N__28117),
            .I(N__28111));
    CascadeMux I__5160 (
            .O(N__28114),
            .I(N__28108));
    Span4Mux_v I__5159 (
            .O(N__28111),
            .I(N__28105));
    InMux I__5158 (
            .O(N__28108),
            .I(N__28102));
    Span4Mux_h I__5157 (
            .O(N__28105),
            .I(N__28099));
    LocalMux I__5156 (
            .O(N__28102),
            .I(N__28096));
    Span4Mux_h I__5155 (
            .O(N__28099),
            .I(N__28093));
    Span12Mux_v I__5154 (
            .O(N__28096),
            .I(N__28090));
    Odrv4 I__5153 (
            .O(N__28093),
            .I(data_index_9_N_258_4));
    Odrv12 I__5152 (
            .O(N__28090),
            .I(data_index_9_N_258_4));
    IoInMux I__5151 (
            .O(N__28085),
            .I(N__28082));
    LocalMux I__5150 (
            .O(N__28082),
            .I(N__28079));
    IoSpan4Mux I__5149 (
            .O(N__28079),
            .I(N__28076));
    Span4Mux_s3_v I__5148 (
            .O(N__28076),
            .I(N__28073));
    Sp12to4 I__5147 (
            .O(N__28073),
            .I(N__28070));
    Span12Mux_s10_v I__5146 (
            .O(N__28070),
            .I(N__28067));
    Span12Mux_h I__5145 (
            .O(N__28067),
            .I(N__28062));
    InMux I__5144 (
            .O(N__28066),
            .I(N__28057));
    InMux I__5143 (
            .O(N__28065),
            .I(N__28057));
    Odrv12 I__5142 (
            .O(N__28062),
            .I(M_OSR0));
    LocalMux I__5141 (
            .O(N__28057),
            .I(M_OSR0));
    InMux I__5140 (
            .O(N__28052),
            .I(N__28049));
    LocalMux I__5139 (
            .O(N__28049),
            .I(N__28046));
    Span4Mux_h I__5138 (
            .O(N__28046),
            .I(N__28043));
    Odrv4 I__5137 (
            .O(N__28043),
            .I(n15555));
    CascadeMux I__5136 (
            .O(N__28040),
            .I(n3_cascade_));
    CascadeMux I__5135 (
            .O(N__28037),
            .I(n10_adj_1242_cascade_));
    InMux I__5134 (
            .O(N__28034),
            .I(N__28031));
    LocalMux I__5133 (
            .O(N__28031),
            .I(n8_adj_1212));
    InMux I__5132 (
            .O(N__28028),
            .I(N__28024));
    InMux I__5131 (
            .O(N__28027),
            .I(N__28021));
    LocalMux I__5130 (
            .O(N__28024),
            .I(eis_end));
    LocalMux I__5129 (
            .O(N__28021),
            .I(eis_end));
    CascadeMux I__5128 (
            .O(N__28016),
            .I(n15171_cascade_));
    InMux I__5127 (
            .O(N__28013),
            .I(N__28010));
    LocalMux I__5126 (
            .O(N__28010),
            .I(N__28007));
    Odrv4 I__5125 (
            .O(N__28007),
            .I(n15475));
    CascadeMux I__5124 (
            .O(N__28004),
            .I(N__28001));
    InMux I__5123 (
            .O(N__28001),
            .I(N__27998));
    LocalMux I__5122 (
            .O(N__27998),
            .I(n15835));
    InMux I__5121 (
            .O(N__27995),
            .I(N__27992));
    LocalMux I__5120 (
            .O(N__27992),
            .I(N__27989));
    Span4Mux_h I__5119 (
            .O(N__27989),
            .I(N__27986));
    Span4Mux_h I__5118 (
            .O(N__27986),
            .I(N__27983));
    Odrv4 I__5117 (
            .O(N__27983),
            .I(n15542));
    InMux I__5116 (
            .O(N__27980),
            .I(N__27977));
    LocalMux I__5115 (
            .O(N__27977),
            .I(N__27974));
    Odrv4 I__5114 (
            .O(N__27974),
            .I(n15679));
    InMux I__5113 (
            .O(N__27971),
            .I(N__27968));
    LocalMux I__5112 (
            .O(N__27968),
            .I(N__27965));
    Span4Mux_v I__5111 (
            .O(N__27965),
            .I(N__27962));
    Odrv4 I__5110 (
            .O(N__27962),
            .I(n15543));
    InMux I__5109 (
            .O(N__27959),
            .I(N__27956));
    LocalMux I__5108 (
            .O(N__27956),
            .I(N__27951));
    InMux I__5107 (
            .O(N__27955),
            .I(N__27948));
    InMux I__5106 (
            .O(N__27954),
            .I(N__27945));
    Span12Mux_s11_h I__5105 (
            .O(N__27951),
            .I(N__27942));
    LocalMux I__5104 (
            .O(N__27948),
            .I(N__27939));
    LocalMux I__5103 (
            .O(N__27945),
            .I(buf_adcdata3_17));
    Odrv12 I__5102 (
            .O(N__27942),
            .I(buf_adcdata3_17));
    Odrv4 I__5101 (
            .O(N__27939),
            .I(buf_adcdata3_17));
    IoInMux I__5100 (
            .O(N__27932),
            .I(N__27929));
    LocalMux I__5099 (
            .O(N__27929),
            .I(N__27926));
    IoSpan4Mux I__5098 (
            .O(N__27926),
            .I(N__27922));
    InMux I__5097 (
            .O(N__27925),
            .I(N__27919));
    Sp12to4 I__5096 (
            .O(N__27922),
            .I(N__27916));
    LocalMux I__5095 (
            .O(N__27919),
            .I(N__27912));
    Span12Mux_v I__5094 (
            .O(N__27916),
            .I(N__27909));
    InMux I__5093 (
            .O(N__27915),
            .I(N__27906));
    Span4Mux_h I__5092 (
            .O(N__27912),
            .I(N__27903));
    Odrv12 I__5091 (
            .O(N__27909),
            .I(M_DCSEL));
    LocalMux I__5090 (
            .O(N__27906),
            .I(M_DCSEL));
    Odrv4 I__5089 (
            .O(N__27903),
            .I(M_DCSEL));
    CascadeMux I__5088 (
            .O(N__27896),
            .I(n90_adj_1023_cascade_));
    InMux I__5087 (
            .O(N__27893),
            .I(N__27890));
    LocalMux I__5086 (
            .O(N__27890),
            .I(n69_adj_1113));
    InMux I__5085 (
            .O(N__27887),
            .I(N__27884));
    LocalMux I__5084 (
            .O(N__27884),
            .I(N__27881));
    Odrv4 I__5083 (
            .O(N__27881),
            .I(n96));
    InMux I__5082 (
            .O(N__27878),
            .I(N__27874));
    InMux I__5081 (
            .O(N__27877),
            .I(N__27871));
    LocalMux I__5080 (
            .O(N__27874),
            .I(buf_device_acadc_4));
    LocalMux I__5079 (
            .O(N__27871),
            .I(buf_device_acadc_4));
    CascadeMux I__5078 (
            .O(N__27866),
            .I(n4814_cascade_));
    CascadeMux I__5077 (
            .O(N__27863),
            .I(N__27857));
    InMux I__5076 (
            .O(N__27862),
            .I(N__27851));
    InMux I__5075 (
            .O(N__27861),
            .I(N__27851));
    InMux I__5074 (
            .O(N__27860),
            .I(N__27848));
    InMux I__5073 (
            .O(N__27857),
            .I(N__27845));
    InMux I__5072 (
            .O(N__27856),
            .I(N__27842));
    LocalMux I__5071 (
            .O(N__27851),
            .I(n5_adj_1235));
    LocalMux I__5070 (
            .O(N__27848),
            .I(n5_adj_1235));
    LocalMux I__5069 (
            .O(N__27845),
            .I(n5_adj_1235));
    LocalMux I__5068 (
            .O(N__27842),
            .I(n5_adj_1235));
    CascadeMux I__5067 (
            .O(N__27833),
            .I(n13475_cascade_));
    CascadeMux I__5066 (
            .O(N__27830),
            .I(n15802_cascade_));
    InMux I__5065 (
            .O(N__27827),
            .I(N__27824));
    LocalMux I__5064 (
            .O(N__27824),
            .I(N__27821));
    Span4Mux_h I__5063 (
            .O(N__27821),
            .I(N__27818));
    Span4Mux_h I__5062 (
            .O(N__27818),
            .I(N__27815));
    Odrv4 I__5061 (
            .O(N__27815),
            .I(n10_adj_1249));
    CascadeMux I__5060 (
            .O(N__27812),
            .I(n15657_cascade_));
    InMux I__5059 (
            .O(N__27809),
            .I(N__27806));
    LocalMux I__5058 (
            .O(N__27806),
            .I(N__27803));
    Span4Mux_h I__5057 (
            .O(N__27803),
            .I(N__27800));
    Span4Mux_h I__5056 (
            .O(N__27800),
            .I(N__27797));
    Odrv4 I__5055 (
            .O(N__27797),
            .I(n13_adj_1042));
    InMux I__5054 (
            .O(N__27794),
            .I(N__27791));
    LocalMux I__5053 (
            .O(N__27791),
            .I(N__27788));
    Span4Mux_h I__5052 (
            .O(N__27788),
            .I(N__27784));
    InMux I__5051 (
            .O(N__27787),
            .I(N__27781));
    Span4Mux_h I__5050 (
            .O(N__27784),
            .I(N__27778));
    LocalMux I__5049 (
            .O(N__27781),
            .I(N__27775));
    Odrv4 I__5048 (
            .O(N__27778),
            .I(\comm_spi.n10479 ));
    Odrv12 I__5047 (
            .O(N__27775),
            .I(\comm_spi.n10479 ));
    SRMux I__5046 (
            .O(N__27770),
            .I(N__27767));
    LocalMux I__5045 (
            .O(N__27767),
            .I(N__27764));
    Span4Mux_v I__5044 (
            .O(N__27764),
            .I(N__27761));
    Odrv4 I__5043 (
            .O(N__27761),
            .I(\comm_spi.data_tx_7__N_806 ));
    InMux I__5042 (
            .O(N__27758),
            .I(N__27755));
    LocalMux I__5041 (
            .O(N__27755),
            .I(N__27752));
    Odrv12 I__5040 (
            .O(N__27752),
            .I(n15576));
    InMux I__5039 (
            .O(N__27749),
            .I(N__27746));
    LocalMux I__5038 (
            .O(N__27746),
            .I(N__27743));
    Span4Mux_v I__5037 (
            .O(N__27743),
            .I(N__27740));
    Odrv4 I__5036 (
            .O(N__27740),
            .I(n15691));
    CascadeMux I__5035 (
            .O(N__27737),
            .I(n15567_cascade_));
    InMux I__5034 (
            .O(N__27734),
            .I(N__27731));
    LocalMux I__5033 (
            .O(N__27731),
            .I(N__27728));
    Span4Mux_h I__5032 (
            .O(N__27728),
            .I(N__27725));
    Odrv4 I__5031 (
            .O(N__27725),
            .I(n7_adj_1255));
    InMux I__5030 (
            .O(N__27722),
            .I(N__27719));
    LocalMux I__5029 (
            .O(N__27719),
            .I(n6));
    CascadeMux I__5028 (
            .O(N__27716),
            .I(n5_adj_1235_cascade_));
    CascadeMux I__5027 (
            .O(N__27713),
            .I(n15535_cascade_));
    CascadeMux I__5026 (
            .O(N__27710),
            .I(n15_cascade_));
    CEMux I__5025 (
            .O(N__27707),
            .I(N__27704));
    LocalMux I__5024 (
            .O(N__27704),
            .I(N__27701));
    Span4Mux_h I__5023 (
            .O(N__27701),
            .I(N__27698));
    Odrv4 I__5022 (
            .O(N__27698),
            .I(n9021));
    InMux I__5021 (
            .O(N__27695),
            .I(N__27692));
    LocalMux I__5020 (
            .O(N__27692),
            .I(n4814));
    InMux I__5019 (
            .O(N__27689),
            .I(N__27680));
    InMux I__5018 (
            .O(N__27688),
            .I(N__27680));
    InMux I__5017 (
            .O(N__27687),
            .I(N__27680));
    LocalMux I__5016 (
            .O(N__27680),
            .I(N__27677));
    Span4Mux_h I__5015 (
            .O(N__27677),
            .I(N__27674));
    Span4Mux_h I__5014 (
            .O(N__27674),
            .I(N__27671));
    Odrv4 I__5013 (
            .O(N__27671),
            .I(comm_tx_buf_6));
    InMux I__5012 (
            .O(N__27668),
            .I(N__27665));
    LocalMux I__5011 (
            .O(N__27665),
            .I(N__27662));
    Span4Mux_v I__5010 (
            .O(N__27662),
            .I(N__27659));
    Span4Mux_h I__5009 (
            .O(N__27659),
            .I(N__27654));
    InMux I__5008 (
            .O(N__27658),
            .I(N__27651));
    InMux I__5007 (
            .O(N__27657),
            .I(N__27648));
    Odrv4 I__5006 (
            .O(N__27654),
            .I(\comm_spi.n16884 ));
    LocalMux I__5005 (
            .O(N__27651),
            .I(\comm_spi.n16884 ));
    LocalMux I__5004 (
            .O(N__27648),
            .I(\comm_spi.n16884 ));
    InMux I__5003 (
            .O(N__27641),
            .I(N__27638));
    LocalMux I__5002 (
            .O(N__27638),
            .I(N__27635));
    Span4Mux_v I__5001 (
            .O(N__27635),
            .I(N__27632));
    Span4Mux_h I__5000 (
            .O(N__27632),
            .I(N__27629));
    Span4Mux_h I__4999 (
            .O(N__27629),
            .I(N__27626));
    Odrv4 I__4998 (
            .O(N__27626),
            .I(buf_data1_23));
    CascadeMux I__4997 (
            .O(N__27623),
            .I(n18_cascade_));
    CascadeMux I__4996 (
            .O(N__27620),
            .I(n15466_cascade_));
    CascadeMux I__4995 (
            .O(N__27617),
            .I(N__27614));
    InMux I__4994 (
            .O(N__27614),
            .I(N__27611));
    LocalMux I__4993 (
            .O(N__27611),
            .I(N__27608));
    Span4Mux_h I__4992 (
            .O(N__27608),
            .I(N__27605));
    Span4Mux_v I__4991 (
            .O(N__27605),
            .I(N__27602));
    Odrv4 I__4990 (
            .O(N__27602),
            .I(n104));
    InMux I__4989 (
            .O(N__27599),
            .I(N__27596));
    LocalMux I__4988 (
            .O(N__27596),
            .I(n56));
    InMux I__4987 (
            .O(N__27593),
            .I(N__27590));
    LocalMux I__4986 (
            .O(N__27590),
            .I(N__27587));
    Span4Mux_h I__4985 (
            .O(N__27587),
            .I(N__27583));
    InMux I__4984 (
            .O(N__27586),
            .I(N__27580));
    Span4Mux_h I__4983 (
            .O(N__27583),
            .I(N__27575));
    LocalMux I__4982 (
            .O(N__27580),
            .I(N__27575));
    Span4Mux_h I__4981 (
            .O(N__27575),
            .I(N__27572));
    Span4Mux_v I__4980 (
            .O(N__27572),
            .I(N__27568));
    InMux I__4979 (
            .O(N__27571),
            .I(N__27565));
    Span4Mux_h I__4978 (
            .O(N__27568),
            .I(N__27562));
    LocalMux I__4977 (
            .O(N__27565),
            .I(buf_adcdata3_1));
    Odrv4 I__4976 (
            .O(N__27562),
            .I(buf_adcdata3_1));
    InMux I__4975 (
            .O(N__27557),
            .I(N__27554));
    LocalMux I__4974 (
            .O(N__27554),
            .I(N__27551));
    Span12Mux_h I__4973 (
            .O(N__27551),
            .I(N__27548));
    Odrv12 I__4972 (
            .O(N__27548),
            .I(buf_data1_1));
    InMux I__4971 (
            .O(N__27545),
            .I(N__27542));
    LocalMux I__4970 (
            .O(N__27542),
            .I(N__27539));
    Span4Mux_h I__4969 (
            .O(N__27539),
            .I(N__27536));
    Span4Mux_h I__4968 (
            .O(N__27536),
            .I(N__27533));
    Odrv4 I__4967 (
            .O(N__27533),
            .I(n4151));
    CascadeMux I__4966 (
            .O(N__27530),
            .I(N__27521));
    CascadeMux I__4965 (
            .O(N__27529),
            .I(N__27518));
    InMux I__4964 (
            .O(N__27528),
            .I(N__27506));
    InMux I__4963 (
            .O(N__27527),
            .I(N__27506));
    InMux I__4962 (
            .O(N__27526),
            .I(N__27503));
    InMux I__4961 (
            .O(N__27525),
            .I(N__27490));
    InMux I__4960 (
            .O(N__27524),
            .I(N__27490));
    InMux I__4959 (
            .O(N__27521),
            .I(N__27490));
    InMux I__4958 (
            .O(N__27518),
            .I(N__27490));
    InMux I__4957 (
            .O(N__27517),
            .I(N__27490));
    InMux I__4956 (
            .O(N__27516),
            .I(N__27490));
    CascadeMux I__4955 (
            .O(N__27515),
            .I(N__27486));
    CascadeMux I__4954 (
            .O(N__27514),
            .I(N__27479));
    CascadeMux I__4953 (
            .O(N__27513),
            .I(N__27476));
    CascadeMux I__4952 (
            .O(N__27512),
            .I(N__27473));
    InMux I__4951 (
            .O(N__27511),
            .I(N__27461));
    LocalMux I__4950 (
            .O(N__27506),
            .I(N__27454));
    LocalMux I__4949 (
            .O(N__27503),
            .I(N__27454));
    LocalMux I__4948 (
            .O(N__27490),
            .I(N__27444));
    InMux I__4947 (
            .O(N__27489),
            .I(N__27441));
    InMux I__4946 (
            .O(N__27486),
            .I(N__27438));
    InMux I__4945 (
            .O(N__27485),
            .I(N__27429));
    InMux I__4944 (
            .O(N__27484),
            .I(N__27429));
    InMux I__4943 (
            .O(N__27483),
            .I(N__27429));
    InMux I__4942 (
            .O(N__27482),
            .I(N__27429));
    InMux I__4941 (
            .O(N__27479),
            .I(N__27416));
    InMux I__4940 (
            .O(N__27476),
            .I(N__27416));
    InMux I__4939 (
            .O(N__27473),
            .I(N__27416));
    InMux I__4938 (
            .O(N__27472),
            .I(N__27416));
    InMux I__4937 (
            .O(N__27471),
            .I(N__27416));
    InMux I__4936 (
            .O(N__27470),
            .I(N__27416));
    CascadeMux I__4935 (
            .O(N__27469),
            .I(N__27412));
    InMux I__4934 (
            .O(N__27468),
            .I(N__27407));
    CascadeMux I__4933 (
            .O(N__27467),
            .I(N__27404));
    InMux I__4932 (
            .O(N__27466),
            .I(N__27400));
    CascadeMux I__4931 (
            .O(N__27465),
            .I(N__27395));
    InMux I__4930 (
            .O(N__27464),
            .I(N__27390));
    LocalMux I__4929 (
            .O(N__27461),
            .I(N__27387));
    InMux I__4928 (
            .O(N__27460),
            .I(N__27384));
    InMux I__4927 (
            .O(N__27459),
            .I(N__27381));
    Span4Mux_h I__4926 (
            .O(N__27454),
            .I(N__27369));
    InMux I__4925 (
            .O(N__27453),
            .I(N__27354));
    InMux I__4924 (
            .O(N__27452),
            .I(N__27354));
    InMux I__4923 (
            .O(N__27451),
            .I(N__27354));
    InMux I__4922 (
            .O(N__27450),
            .I(N__27354));
    InMux I__4921 (
            .O(N__27449),
            .I(N__27354));
    InMux I__4920 (
            .O(N__27448),
            .I(N__27354));
    InMux I__4919 (
            .O(N__27447),
            .I(N__27354));
    Span4Mux_v I__4918 (
            .O(N__27444),
            .I(N__27347));
    LocalMux I__4917 (
            .O(N__27441),
            .I(N__27347));
    LocalMux I__4916 (
            .O(N__27438),
            .I(N__27340));
    LocalMux I__4915 (
            .O(N__27429),
            .I(N__27340));
    LocalMux I__4914 (
            .O(N__27416),
            .I(N__27340));
    InMux I__4913 (
            .O(N__27415),
            .I(N__27337));
    InMux I__4912 (
            .O(N__27412),
            .I(N__27329));
    InMux I__4911 (
            .O(N__27411),
            .I(N__27329));
    InMux I__4910 (
            .O(N__27410),
            .I(N__27329));
    LocalMux I__4909 (
            .O(N__27407),
            .I(N__27326));
    InMux I__4908 (
            .O(N__27404),
            .I(N__27323));
    InMux I__4907 (
            .O(N__27403),
            .I(N__27319));
    LocalMux I__4906 (
            .O(N__27400),
            .I(N__27316));
    InMux I__4905 (
            .O(N__27399),
            .I(N__27305));
    InMux I__4904 (
            .O(N__27398),
            .I(N__27305));
    InMux I__4903 (
            .O(N__27395),
            .I(N__27305));
    InMux I__4902 (
            .O(N__27394),
            .I(N__27305));
    InMux I__4901 (
            .O(N__27393),
            .I(N__27305));
    LocalMux I__4900 (
            .O(N__27390),
            .I(N__27302));
    Span4Mux_v I__4899 (
            .O(N__27387),
            .I(N__27299));
    LocalMux I__4898 (
            .O(N__27384),
            .I(N__27294));
    LocalMux I__4897 (
            .O(N__27381),
            .I(N__27294));
    InMux I__4896 (
            .O(N__27380),
            .I(N__27289));
    InMux I__4895 (
            .O(N__27379),
            .I(N__27289));
    InMux I__4894 (
            .O(N__27378),
            .I(N__27273));
    InMux I__4893 (
            .O(N__27377),
            .I(N__27273));
    InMux I__4892 (
            .O(N__27376),
            .I(N__27273));
    InMux I__4891 (
            .O(N__27375),
            .I(N__27273));
    InMux I__4890 (
            .O(N__27374),
            .I(N__27273));
    InMux I__4889 (
            .O(N__27373),
            .I(N__27273));
    InMux I__4888 (
            .O(N__27372),
            .I(N__27273));
    Span4Mux_v I__4887 (
            .O(N__27369),
            .I(N__27270));
    LocalMux I__4886 (
            .O(N__27354),
            .I(N__27267));
    CascadeMux I__4885 (
            .O(N__27353),
            .I(N__27264));
    InMux I__4884 (
            .O(N__27352),
            .I(N__27261));
    Span4Mux_h I__4883 (
            .O(N__27347),
            .I(N__27258));
    Span4Mux_v I__4882 (
            .O(N__27340),
            .I(N__27253));
    LocalMux I__4881 (
            .O(N__27337),
            .I(N__27253));
    InMux I__4880 (
            .O(N__27336),
            .I(N__27247));
    LocalMux I__4879 (
            .O(N__27329),
            .I(N__27244));
    Span4Mux_h I__4878 (
            .O(N__27326),
            .I(N__27239));
    LocalMux I__4877 (
            .O(N__27323),
            .I(N__27239));
    CascadeMux I__4876 (
            .O(N__27322),
            .I(N__27231));
    LocalMux I__4875 (
            .O(N__27319),
            .I(N__27222));
    Span4Mux_h I__4874 (
            .O(N__27316),
            .I(N__27222));
    LocalMux I__4873 (
            .O(N__27305),
            .I(N__27222));
    Span4Mux_v I__4872 (
            .O(N__27302),
            .I(N__27215));
    Span4Mux_v I__4871 (
            .O(N__27299),
            .I(N__27215));
    Span4Mux_h I__4870 (
            .O(N__27294),
            .I(N__27215));
    LocalMux I__4869 (
            .O(N__27289),
            .I(N__27212));
    InMux I__4868 (
            .O(N__27288),
            .I(N__27209));
    LocalMux I__4867 (
            .O(N__27273),
            .I(N__27202));
    Span4Mux_v I__4866 (
            .O(N__27270),
            .I(N__27202));
    Span4Mux_h I__4865 (
            .O(N__27267),
            .I(N__27202));
    InMux I__4864 (
            .O(N__27264),
            .I(N__27199));
    LocalMux I__4863 (
            .O(N__27261),
            .I(N__27194));
    Sp12to4 I__4862 (
            .O(N__27258),
            .I(N__27194));
    Sp12to4 I__4861 (
            .O(N__27253),
            .I(N__27191));
    InMux I__4860 (
            .O(N__27252),
            .I(N__27188));
    InMux I__4859 (
            .O(N__27251),
            .I(N__27183));
    InMux I__4858 (
            .O(N__27250),
            .I(N__27183));
    LocalMux I__4857 (
            .O(N__27247),
            .I(N__27180));
    Span4Mux_v I__4856 (
            .O(N__27244),
            .I(N__27175));
    Span4Mux_h I__4855 (
            .O(N__27239),
            .I(N__27175));
    InMux I__4854 (
            .O(N__27238),
            .I(N__27172));
    InMux I__4853 (
            .O(N__27237),
            .I(N__27161));
    InMux I__4852 (
            .O(N__27236),
            .I(N__27161));
    InMux I__4851 (
            .O(N__27235),
            .I(N__27161));
    InMux I__4850 (
            .O(N__27234),
            .I(N__27161));
    InMux I__4849 (
            .O(N__27231),
            .I(N__27161));
    InMux I__4848 (
            .O(N__27230),
            .I(N__27156));
    InMux I__4847 (
            .O(N__27229),
            .I(N__27156));
    Span4Mux_v I__4846 (
            .O(N__27222),
            .I(N__27151));
    Span4Mux_h I__4845 (
            .O(N__27215),
            .I(N__27151));
    Span4Mux_h I__4844 (
            .O(N__27212),
            .I(N__27144));
    LocalMux I__4843 (
            .O(N__27209),
            .I(N__27144));
    Span4Mux_h I__4842 (
            .O(N__27202),
            .I(N__27144));
    LocalMux I__4841 (
            .O(N__27199),
            .I(N__27137));
    Span12Mux_v I__4840 (
            .O(N__27194),
            .I(N__27137));
    Span12Mux_h I__4839 (
            .O(N__27191),
            .I(N__27137));
    LocalMux I__4838 (
            .O(N__27188),
            .I(adc_state_0_adj_1117));
    LocalMux I__4837 (
            .O(N__27183),
            .I(adc_state_0_adj_1117));
    Odrv4 I__4836 (
            .O(N__27180),
            .I(adc_state_0_adj_1117));
    Odrv4 I__4835 (
            .O(N__27175),
            .I(adc_state_0_adj_1117));
    LocalMux I__4834 (
            .O(N__27172),
            .I(adc_state_0_adj_1117));
    LocalMux I__4833 (
            .O(N__27161),
            .I(adc_state_0_adj_1117));
    LocalMux I__4832 (
            .O(N__27156),
            .I(adc_state_0_adj_1117));
    Odrv4 I__4831 (
            .O(N__27151),
            .I(adc_state_0_adj_1117));
    Odrv4 I__4830 (
            .O(N__27144),
            .I(adc_state_0_adj_1117));
    Odrv12 I__4829 (
            .O(N__27137),
            .I(adc_state_0_adj_1117));
    InMux I__4828 (
            .O(N__27116),
            .I(N__27106));
    InMux I__4827 (
            .O(N__27115),
            .I(N__27101));
    CascadeMux I__4826 (
            .O(N__27114),
            .I(N__27098));
    InMux I__4825 (
            .O(N__27113),
            .I(N__27092));
    InMux I__4824 (
            .O(N__27112),
            .I(N__27087));
    InMux I__4823 (
            .O(N__27111),
            .I(N__27087));
    InMux I__4822 (
            .O(N__27110),
            .I(N__27082));
    InMux I__4821 (
            .O(N__27109),
            .I(N__27082));
    LocalMux I__4820 (
            .O(N__27106),
            .I(N__27079));
    InMux I__4819 (
            .O(N__27105),
            .I(N__27076));
    InMux I__4818 (
            .O(N__27104),
            .I(N__27073));
    LocalMux I__4817 (
            .O(N__27101),
            .I(N__27070));
    InMux I__4816 (
            .O(N__27098),
            .I(N__27067));
    InMux I__4815 (
            .O(N__27097),
            .I(N__27060));
    InMux I__4814 (
            .O(N__27096),
            .I(N__27060));
    InMux I__4813 (
            .O(N__27095),
            .I(N__27060));
    LocalMux I__4812 (
            .O(N__27092),
            .I(N__27053));
    LocalMux I__4811 (
            .O(N__27087),
            .I(N__27053));
    LocalMux I__4810 (
            .O(N__27082),
            .I(N__27053));
    Span4Mux_v I__4809 (
            .O(N__27079),
            .I(N__27048));
    LocalMux I__4808 (
            .O(N__27076),
            .I(N__27048));
    LocalMux I__4807 (
            .O(N__27073),
            .I(DTRIG_N_957_adj_1150));
    Odrv12 I__4806 (
            .O(N__27070),
            .I(DTRIG_N_957_adj_1150));
    LocalMux I__4805 (
            .O(N__27067),
            .I(DTRIG_N_957_adj_1150));
    LocalMux I__4804 (
            .O(N__27060),
            .I(DTRIG_N_957_adj_1150));
    Odrv4 I__4803 (
            .O(N__27053),
            .I(DTRIG_N_957_adj_1150));
    Odrv4 I__4802 (
            .O(N__27048),
            .I(DTRIG_N_957_adj_1150));
    InMux I__4801 (
            .O(N__27035),
            .I(N__27030));
    InMux I__4800 (
            .O(N__27034),
            .I(N__27027));
    InMux I__4799 (
            .O(N__27033),
            .I(N__27024));
    LocalMux I__4798 (
            .O(N__27030),
            .I(N__27019));
    LocalMux I__4797 (
            .O(N__27027),
            .I(N__27011));
    LocalMux I__4796 (
            .O(N__27024),
            .I(N__27011));
    InMux I__4795 (
            .O(N__27023),
            .I(N__27002));
    InMux I__4794 (
            .O(N__27022),
            .I(N__27002));
    Span4Mux_v I__4793 (
            .O(N__27019),
            .I(N__26999));
    InMux I__4792 (
            .O(N__27018),
            .I(N__26992));
    InMux I__4791 (
            .O(N__27017),
            .I(N__26992));
    InMux I__4790 (
            .O(N__27016),
            .I(N__26992));
    Span4Mux_h I__4789 (
            .O(N__27011),
            .I(N__26989));
    InMux I__4788 (
            .O(N__27010),
            .I(N__26982));
    InMux I__4787 (
            .O(N__27009),
            .I(N__26982));
    InMux I__4786 (
            .O(N__27008),
            .I(N__26982));
    InMux I__4785 (
            .O(N__27007),
            .I(N__26979));
    LocalMux I__4784 (
            .O(N__27002),
            .I(N__26976));
    Odrv4 I__4783 (
            .O(N__26999),
            .I(adc_state_1_adj_1116));
    LocalMux I__4782 (
            .O(N__26992),
            .I(adc_state_1_adj_1116));
    Odrv4 I__4781 (
            .O(N__26989),
            .I(adc_state_1_adj_1116));
    LocalMux I__4780 (
            .O(N__26982),
            .I(adc_state_1_adj_1116));
    LocalMux I__4779 (
            .O(N__26979),
            .I(adc_state_1_adj_1116));
    Odrv4 I__4778 (
            .O(N__26976),
            .I(adc_state_1_adj_1116));
    CEMux I__4777 (
            .O(N__26963),
            .I(N__26959));
    CEMux I__4776 (
            .O(N__26962),
            .I(N__26956));
    LocalMux I__4775 (
            .O(N__26959),
            .I(N__26951));
    LocalMux I__4774 (
            .O(N__26956),
            .I(N__26951));
    Odrv4 I__4773 (
            .O(N__26951),
            .I(\ADC_VAC4.n12 ));
    SRMux I__4772 (
            .O(N__26948),
            .I(N__26945));
    LocalMux I__4771 (
            .O(N__26945),
            .I(N__26942));
    Odrv12 I__4770 (
            .O(N__26942),
            .I(\ADC_VAC4.n14930 ));
    InMux I__4769 (
            .O(N__26939),
            .I(N__26935));
    InMux I__4768 (
            .O(N__26938),
            .I(N__26932));
    LocalMux I__4767 (
            .O(N__26935),
            .I(\comm_spi.n10467 ));
    LocalMux I__4766 (
            .O(N__26932),
            .I(\comm_spi.n10467 ));
    InMux I__4765 (
            .O(N__26927),
            .I(N__26924));
    LocalMux I__4764 (
            .O(N__26924),
            .I(N__26920));
    InMux I__4763 (
            .O(N__26923),
            .I(N__26917));
    Odrv4 I__4762 (
            .O(N__26920),
            .I(\comm_spi.n10468 ));
    LocalMux I__4761 (
            .O(N__26917),
            .I(\comm_spi.n10468 ));
    SRMux I__4760 (
            .O(N__26912),
            .I(N__26909));
    LocalMux I__4759 (
            .O(N__26909),
            .I(N__26906));
    Span4Mux_v I__4758 (
            .O(N__26906),
            .I(N__26903));
    Odrv4 I__4757 (
            .O(N__26903),
            .I(\comm_spi.data_tx_7__N_822 ));
    IoInMux I__4756 (
            .O(N__26900),
            .I(N__26897));
    LocalMux I__4755 (
            .O(N__26897),
            .I(N__26894));
    IoSpan4Mux I__4754 (
            .O(N__26894),
            .I(N__26891));
    Span4Mux_s0_v I__4753 (
            .O(N__26891),
            .I(N__26888));
    Sp12to4 I__4752 (
            .O(N__26888),
            .I(N__26885));
    Span12Mux_h I__4751 (
            .O(N__26885),
            .I(N__26882));
    Odrv12 I__4750 (
            .O(N__26882),
            .I(DDS_CS1));
    InMux I__4749 (
            .O(N__26879),
            .I(N__26870));
    InMux I__4748 (
            .O(N__26878),
            .I(N__26870));
    InMux I__4747 (
            .O(N__26877),
            .I(N__26870));
    LocalMux I__4746 (
            .O(N__26870),
            .I(N__26867));
    Span4Mux_h I__4745 (
            .O(N__26867),
            .I(N__26864));
    Odrv4 I__4744 (
            .O(N__26864),
            .I(comm_tx_buf_7));
    CascadeMux I__4743 (
            .O(N__26861),
            .I(n15156_cascade_));
    InMux I__4742 (
            .O(N__26858),
            .I(N__26829));
    InMux I__4741 (
            .O(N__26857),
            .I(N__26820));
    InMux I__4740 (
            .O(N__26856),
            .I(N__26820));
    InMux I__4739 (
            .O(N__26855),
            .I(N__26820));
    InMux I__4738 (
            .O(N__26854),
            .I(N__26820));
    InMux I__4737 (
            .O(N__26853),
            .I(N__26813));
    InMux I__4736 (
            .O(N__26852),
            .I(N__26813));
    InMux I__4735 (
            .O(N__26851),
            .I(N__26813));
    InMux I__4734 (
            .O(N__26850),
            .I(N__26807));
    InMux I__4733 (
            .O(N__26849),
            .I(N__26804));
    InMux I__4732 (
            .O(N__26848),
            .I(N__26801));
    InMux I__4731 (
            .O(N__26847),
            .I(N__26798));
    InMux I__4730 (
            .O(N__26846),
            .I(N__26794));
    InMux I__4729 (
            .O(N__26845),
            .I(N__26791));
    InMux I__4728 (
            .O(N__26844),
            .I(N__26782));
    InMux I__4727 (
            .O(N__26843),
            .I(N__26782));
    InMux I__4726 (
            .O(N__26842),
            .I(N__26782));
    InMux I__4725 (
            .O(N__26841),
            .I(N__26782));
    InMux I__4724 (
            .O(N__26840),
            .I(N__26775));
    InMux I__4723 (
            .O(N__26839),
            .I(N__26775));
    InMux I__4722 (
            .O(N__26838),
            .I(N__26775));
    InMux I__4721 (
            .O(N__26837),
            .I(N__26762));
    InMux I__4720 (
            .O(N__26836),
            .I(N__26762));
    InMux I__4719 (
            .O(N__26835),
            .I(N__26762));
    InMux I__4718 (
            .O(N__26834),
            .I(N__26762));
    InMux I__4717 (
            .O(N__26833),
            .I(N__26762));
    InMux I__4716 (
            .O(N__26832),
            .I(N__26762));
    LocalMux I__4715 (
            .O(N__26829),
            .I(N__26757));
    LocalMux I__4714 (
            .O(N__26820),
            .I(N__26757));
    LocalMux I__4713 (
            .O(N__26813),
            .I(N__26754));
    InMux I__4712 (
            .O(N__26812),
            .I(N__26746));
    InMux I__4711 (
            .O(N__26811),
            .I(N__26746));
    InMux I__4710 (
            .O(N__26810),
            .I(N__26746));
    LocalMux I__4709 (
            .O(N__26807),
            .I(N__26743));
    LocalMux I__4708 (
            .O(N__26804),
            .I(N__26736));
    LocalMux I__4707 (
            .O(N__26801),
            .I(N__26736));
    LocalMux I__4706 (
            .O(N__26798),
            .I(N__26736));
    InMux I__4705 (
            .O(N__26797),
            .I(N__26733));
    LocalMux I__4704 (
            .O(N__26794),
            .I(N__26722));
    LocalMux I__4703 (
            .O(N__26791),
            .I(N__26722));
    LocalMux I__4702 (
            .O(N__26782),
            .I(N__26722));
    LocalMux I__4701 (
            .O(N__26775),
            .I(N__26722));
    LocalMux I__4700 (
            .O(N__26762),
            .I(N__26722));
    Span4Mux_v I__4699 (
            .O(N__26757),
            .I(N__26719));
    Span4Mux_v I__4698 (
            .O(N__26754),
            .I(N__26716));
    InMux I__4697 (
            .O(N__26753),
            .I(N__26713));
    LocalMux I__4696 (
            .O(N__26746),
            .I(N__26710));
    Span4Mux_h I__4695 (
            .O(N__26743),
            .I(N__26705));
    Span4Mux_v I__4694 (
            .O(N__26736),
            .I(N__26705));
    LocalMux I__4693 (
            .O(N__26733),
            .I(N__26700));
    Span12Mux_v I__4692 (
            .O(N__26722),
            .I(N__26700));
    Span4Mux_h I__4691 (
            .O(N__26719),
            .I(N__26695));
    Span4Mux_v I__4690 (
            .O(N__26716),
            .I(N__26695));
    LocalMux I__4689 (
            .O(N__26713),
            .I(n9694));
    Odrv12 I__4688 (
            .O(N__26710),
            .I(n9694));
    Odrv4 I__4687 (
            .O(N__26705),
            .I(n9694));
    Odrv12 I__4686 (
            .O(N__26700),
            .I(n9694));
    Odrv4 I__4685 (
            .O(N__26695),
            .I(n9694));
    CascadeMux I__4684 (
            .O(N__26684),
            .I(\ADC_VAC4.n15257_cascade_ ));
    CEMux I__4683 (
            .O(N__26681),
            .I(N__26678));
    LocalMux I__4682 (
            .O(N__26678),
            .I(\ADC_VAC4.n15258 ));
    InMux I__4681 (
            .O(N__26675),
            .I(N__26672));
    LocalMux I__4680 (
            .O(N__26672),
            .I(\ADC_VAC4.n15278 ));
    CascadeMux I__4679 (
            .O(N__26669),
            .I(N__26666));
    InMux I__4678 (
            .O(N__26666),
            .I(N__26661));
    CascadeMux I__4677 (
            .O(N__26665),
            .I(N__26658));
    CascadeMux I__4676 (
            .O(N__26664),
            .I(N__26654));
    LocalMux I__4675 (
            .O(N__26661),
            .I(N__26651));
    InMux I__4674 (
            .O(N__26658),
            .I(N__26648));
    InMux I__4673 (
            .O(N__26657),
            .I(N__26643));
    InMux I__4672 (
            .O(N__26654),
            .I(N__26643));
    Span4Mux_h I__4671 (
            .O(N__26651),
            .I(N__26638));
    LocalMux I__4670 (
            .O(N__26648),
            .I(N__26638));
    LocalMux I__4669 (
            .O(N__26643),
            .I(N__26633));
    Span4Mux_v I__4668 (
            .O(N__26638),
            .I(N__26630));
    InMux I__4667 (
            .O(N__26637),
            .I(N__26625));
    InMux I__4666 (
            .O(N__26636),
            .I(N__26625));
    Span12Mux_v I__4665 (
            .O(N__26633),
            .I(N__26620));
    Sp12to4 I__4664 (
            .O(N__26630),
            .I(N__26620));
    LocalMux I__4663 (
            .O(N__26625),
            .I(N__26617));
    Span12Mux_h I__4662 (
            .O(N__26620),
            .I(N__26614));
    Span12Mux_h I__4661 (
            .O(N__26617),
            .I(N__26611));
    Odrv12 I__4660 (
            .O(N__26614),
            .I(M_DRDY4));
    Odrv12 I__4659 (
            .O(N__26611),
            .I(M_DRDY4));
    CascadeMux I__4658 (
            .O(N__26606),
            .I(n14_cascade_));
    InMux I__4657 (
            .O(N__26603),
            .I(N__26600));
    LocalMux I__4656 (
            .O(N__26600),
            .I(N__26597));
    Odrv4 I__4655 (
            .O(N__26597),
            .I(n15156));
    IoInMux I__4654 (
            .O(N__26594),
            .I(N__26591));
    LocalMux I__4653 (
            .O(N__26591),
            .I(N__26588));
    Span4Mux_s1_v I__4652 (
            .O(N__26588),
            .I(N__26585));
    Span4Mux_v I__4651 (
            .O(N__26585),
            .I(N__26582));
    Span4Mux_v I__4650 (
            .O(N__26582),
            .I(N__26578));
    CascadeMux I__4649 (
            .O(N__26581),
            .I(N__26575));
    Sp12to4 I__4648 (
            .O(N__26578),
            .I(N__26572));
    InMux I__4647 (
            .O(N__26575),
            .I(N__26569));
    Odrv12 I__4646 (
            .O(N__26572),
            .I(M_CS4));
    LocalMux I__4645 (
            .O(N__26569),
            .I(M_CS4));
    InMux I__4644 (
            .O(N__26564),
            .I(N__26561));
    LocalMux I__4643 (
            .O(N__26561),
            .I(N__26558));
    Sp12to4 I__4642 (
            .O(N__26558),
            .I(N__26555));
    Odrv12 I__4641 (
            .O(N__26555),
            .I(buf_data2_11));
    InMux I__4640 (
            .O(N__26552),
            .I(N__26549));
    LocalMux I__4639 (
            .O(N__26549),
            .I(N__26545));
    CascadeMux I__4638 (
            .O(N__26548),
            .I(N__26542));
    Span4Mux_v I__4637 (
            .O(N__26545),
            .I(N__26538));
    InMux I__4636 (
            .O(N__26542),
            .I(N__26535));
    InMux I__4635 (
            .O(N__26541),
            .I(N__26532));
    Span4Mux_h I__4634 (
            .O(N__26538),
            .I(N__26529));
    LocalMux I__4633 (
            .O(N__26535),
            .I(N__26526));
    LocalMux I__4632 (
            .O(N__26532),
            .I(N__26519));
    Span4Mux_h I__4631 (
            .O(N__26529),
            .I(N__26519));
    Span4Mux_v I__4630 (
            .O(N__26526),
            .I(N__26519));
    Odrv4 I__4629 (
            .O(N__26519),
            .I(buf_adcdata4_11));
    InMux I__4628 (
            .O(N__26516),
            .I(N__26513));
    LocalMux I__4627 (
            .O(N__26513),
            .I(N__26510));
    Span4Mux_h I__4626 (
            .O(N__26510),
            .I(N__26507));
    Span4Mux_v I__4625 (
            .O(N__26507),
            .I(N__26504));
    Span4Mux_h I__4624 (
            .O(N__26504),
            .I(N__26501));
    Odrv4 I__4623 (
            .O(N__26501),
            .I(n4061));
    InMux I__4622 (
            .O(N__26498),
            .I(N__26495));
    LocalMux I__4621 (
            .O(N__26495),
            .I(\ADC_VAC4.n17 ));
    CascadeMux I__4620 (
            .O(N__26492),
            .I(N__26489));
    InMux I__4619 (
            .O(N__26489),
            .I(N__26485));
    InMux I__4618 (
            .O(N__26488),
            .I(N__26482));
    LocalMux I__4617 (
            .O(N__26485),
            .I(N__26478));
    LocalMux I__4616 (
            .O(N__26482),
            .I(N__26475));
    InMux I__4615 (
            .O(N__26481),
            .I(N__26472));
    Odrv4 I__4614 (
            .O(N__26478),
            .I(cmd_rdadctmp_26_adj_1086));
    Odrv4 I__4613 (
            .O(N__26475),
            .I(cmd_rdadctmp_26_adj_1086));
    LocalMux I__4612 (
            .O(N__26472),
            .I(cmd_rdadctmp_26_adj_1086));
    InMux I__4611 (
            .O(N__26465),
            .I(N__26462));
    LocalMux I__4610 (
            .O(N__26462),
            .I(N__26459));
    Span4Mux_h I__4609 (
            .O(N__26459),
            .I(N__26455));
    InMux I__4608 (
            .O(N__26458),
            .I(N__26452));
    Span4Mux_v I__4607 (
            .O(N__26455),
            .I(N__26448));
    LocalMux I__4606 (
            .O(N__26452),
            .I(N__26445));
    InMux I__4605 (
            .O(N__26451),
            .I(N__26442));
    Span4Mux_h I__4604 (
            .O(N__26448),
            .I(N__26437));
    Span4Mux_v I__4603 (
            .O(N__26445),
            .I(N__26437));
    LocalMux I__4602 (
            .O(N__26442),
            .I(buf_adcdata3_18));
    Odrv4 I__4601 (
            .O(N__26437),
            .I(buf_adcdata3_18));
    InMux I__4600 (
            .O(N__26432),
            .I(N__26429));
    LocalMux I__4599 (
            .O(N__26429),
            .I(N__26426));
    Span4Mux_h I__4598 (
            .O(N__26426),
            .I(N__26423));
    Odrv4 I__4597 (
            .O(N__26423),
            .I(n15811));
    CascadeMux I__4596 (
            .O(N__26420),
            .I(N__26417));
    InMux I__4595 (
            .O(N__26417),
            .I(N__26413));
    InMux I__4594 (
            .O(N__26416),
            .I(N__26410));
    LocalMux I__4593 (
            .O(N__26413),
            .I(N__26405));
    LocalMux I__4592 (
            .O(N__26410),
            .I(N__26405));
    Span4Mux_h I__4591 (
            .O(N__26405),
            .I(N__26401));
    InMux I__4590 (
            .O(N__26404),
            .I(N__26398));
    Odrv4 I__4589 (
            .O(N__26401),
            .I(cmd_rdadctmp_21_adj_1128));
    LocalMux I__4588 (
            .O(N__26398),
            .I(cmd_rdadctmp_21_adj_1128));
    InMux I__4587 (
            .O(N__26393),
            .I(N__26389));
    InMux I__4586 (
            .O(N__26392),
            .I(N__26385));
    LocalMux I__4585 (
            .O(N__26389),
            .I(N__26382));
    CascadeMux I__4584 (
            .O(N__26388),
            .I(N__26379));
    LocalMux I__4583 (
            .O(N__26385),
            .I(N__26376));
    Span4Mux_h I__4582 (
            .O(N__26382),
            .I(N__26373));
    InMux I__4581 (
            .O(N__26379),
            .I(N__26370));
    Odrv4 I__4580 (
            .O(N__26376),
            .I(cmd_rdadctmp_22_adj_1127));
    Odrv4 I__4579 (
            .O(N__26373),
            .I(cmd_rdadctmp_22_adj_1127));
    LocalMux I__4578 (
            .O(N__26370),
            .I(cmd_rdadctmp_22_adj_1127));
    InMux I__4577 (
            .O(N__26363),
            .I(N__26359));
    InMux I__4576 (
            .O(N__26362),
            .I(N__26356));
    LocalMux I__4575 (
            .O(N__26359),
            .I(N__26352));
    LocalMux I__4574 (
            .O(N__26356),
            .I(N__26349));
    InMux I__4573 (
            .O(N__26355),
            .I(N__26346));
    Span12Mux_h I__4572 (
            .O(N__26352),
            .I(N__26343));
    Span4Mux_v I__4571 (
            .O(N__26349),
            .I(N__26340));
    LocalMux I__4570 (
            .O(N__26346),
            .I(buf_adcdata3_16));
    Odrv12 I__4569 (
            .O(N__26343),
            .I(buf_adcdata3_16));
    Odrv4 I__4568 (
            .O(N__26340),
            .I(buf_adcdata3_16));
    InMux I__4567 (
            .O(N__26333),
            .I(N__26330));
    LocalMux I__4566 (
            .O(N__26330),
            .I(n90));
    CascadeMux I__4565 (
            .O(N__26327),
            .I(N__26322));
    InMux I__4564 (
            .O(N__26326),
            .I(N__26319));
    InMux I__4563 (
            .O(N__26325),
            .I(N__26314));
    InMux I__4562 (
            .O(N__26322),
            .I(N__26314));
    LocalMux I__4561 (
            .O(N__26319),
            .I(cmd_rdadctmp_23_adj_1126));
    LocalMux I__4560 (
            .O(N__26314),
            .I(cmd_rdadctmp_23_adj_1126));
    InMux I__4559 (
            .O(N__26309),
            .I(N__26304));
    InMux I__4558 (
            .O(N__26308),
            .I(N__26299));
    InMux I__4557 (
            .O(N__26307),
            .I(N__26299));
    LocalMux I__4556 (
            .O(N__26304),
            .I(cmd_rdadctmp_24_adj_1125));
    LocalMux I__4555 (
            .O(N__26299),
            .I(cmd_rdadctmp_24_adj_1125));
    CascadeMux I__4554 (
            .O(N__26294),
            .I(N__26290));
    CascadeMux I__4553 (
            .O(N__26293),
            .I(N__26286));
    InMux I__4552 (
            .O(N__26290),
            .I(N__26281));
    InMux I__4551 (
            .O(N__26289),
            .I(N__26281));
    InMux I__4550 (
            .O(N__26286),
            .I(N__26278));
    LocalMux I__4549 (
            .O(N__26281),
            .I(N__26275));
    LocalMux I__4548 (
            .O(N__26278),
            .I(N__26272));
    Odrv4 I__4547 (
            .O(N__26275),
            .I(cmd_rdadctmp_25_adj_1124));
    Odrv4 I__4546 (
            .O(N__26272),
            .I(cmd_rdadctmp_25_adj_1124));
    IoInMux I__4545 (
            .O(N__26267),
            .I(N__26264));
    LocalMux I__4544 (
            .O(N__26264),
            .I(N__26261));
    Span4Mux_s1_v I__4543 (
            .O(N__26261),
            .I(N__26258));
    Sp12to4 I__4542 (
            .O(N__26258),
            .I(N__26254));
    InMux I__4541 (
            .O(N__26257),
            .I(N__26250));
    Span12Mux_h I__4540 (
            .O(N__26254),
            .I(N__26247));
    CascadeMux I__4539 (
            .O(N__26253),
            .I(N__26244));
    LocalMux I__4538 (
            .O(N__26250),
            .I(N__26241));
    Span12Mux_v I__4537 (
            .O(N__26247),
            .I(N__26238));
    InMux I__4536 (
            .O(N__26244),
            .I(N__26235));
    Span4Mux_h I__4535 (
            .O(N__26241),
            .I(N__26232));
    Odrv12 I__4534 (
            .O(N__26238),
            .I(M_POW));
    LocalMux I__4533 (
            .O(N__26235),
            .I(M_POW));
    Odrv4 I__4532 (
            .O(N__26232),
            .I(M_POW));
    InMux I__4531 (
            .O(N__26225),
            .I(N__26222));
    LocalMux I__4530 (
            .O(N__26222),
            .I(N__26219));
    Span4Mux_v I__4529 (
            .O(N__26219),
            .I(N__26216));
    Span4Mux_h I__4528 (
            .O(N__26216),
            .I(N__26213));
    Span4Mux_h I__4527 (
            .O(N__26213),
            .I(N__26208));
    InMux I__4526 (
            .O(N__26212),
            .I(N__26205));
    InMux I__4525 (
            .O(N__26211),
            .I(N__26202));
    Span4Mux_h I__4524 (
            .O(N__26208),
            .I(N__26199));
    LocalMux I__4523 (
            .O(N__26205),
            .I(buf_adcdata3_19));
    LocalMux I__4522 (
            .O(N__26202),
            .I(buf_adcdata3_19));
    Odrv4 I__4521 (
            .O(N__26199),
            .I(buf_adcdata3_19));
    InMux I__4520 (
            .O(N__26192),
            .I(N__26189));
    LocalMux I__4519 (
            .O(N__26189),
            .I(n87));
    InMux I__4518 (
            .O(N__26186),
            .I(N__26172));
    InMux I__4517 (
            .O(N__26185),
            .I(N__26172));
    InMux I__4516 (
            .O(N__26184),
            .I(N__26167));
    InMux I__4515 (
            .O(N__26183),
            .I(N__26167));
    InMux I__4514 (
            .O(N__26182),
            .I(N__26164));
    InMux I__4513 (
            .O(N__26181),
            .I(N__26154));
    InMux I__4512 (
            .O(N__26180),
            .I(N__26149));
    InMux I__4511 (
            .O(N__26179),
            .I(N__26149));
    InMux I__4510 (
            .O(N__26178),
            .I(N__26144));
    InMux I__4509 (
            .O(N__26177),
            .I(N__26144));
    LocalMux I__4508 (
            .O(N__26172),
            .I(N__26139));
    LocalMux I__4507 (
            .O(N__26167),
            .I(N__26139));
    LocalMux I__4506 (
            .O(N__26164),
            .I(N__26136));
    InMux I__4505 (
            .O(N__26163),
            .I(N__26131));
    InMux I__4504 (
            .O(N__26162),
            .I(N__26131));
    InMux I__4503 (
            .O(N__26161),
            .I(N__26128));
    InMux I__4502 (
            .O(N__26160),
            .I(N__26117));
    InMux I__4501 (
            .O(N__26159),
            .I(N__26117));
    InMux I__4500 (
            .O(N__26158),
            .I(N__26117));
    InMux I__4499 (
            .O(N__26157),
            .I(N__26117));
    LocalMux I__4498 (
            .O(N__26154),
            .I(N__26110));
    LocalMux I__4497 (
            .O(N__26149),
            .I(N__26105));
    LocalMux I__4496 (
            .O(N__26144),
            .I(N__26105));
    Span4Mux_v I__4495 (
            .O(N__26139),
            .I(N__26096));
    Span4Mux_h I__4494 (
            .O(N__26136),
            .I(N__26096));
    LocalMux I__4493 (
            .O(N__26131),
            .I(N__26096));
    LocalMux I__4492 (
            .O(N__26128),
            .I(N__26096));
    InMux I__4491 (
            .O(N__26127),
            .I(N__26093));
    InMux I__4490 (
            .O(N__26126),
            .I(N__26090));
    LocalMux I__4489 (
            .O(N__26117),
            .I(N__26085));
    InMux I__4488 (
            .O(N__26116),
            .I(N__26076));
    InMux I__4487 (
            .O(N__26115),
            .I(N__26076));
    InMux I__4486 (
            .O(N__26114),
            .I(N__26076));
    InMux I__4485 (
            .O(N__26113),
            .I(N__26076));
    Span4Mux_h I__4484 (
            .O(N__26110),
            .I(N__26066));
    Span4Mux_h I__4483 (
            .O(N__26105),
            .I(N__26063));
    Span4Mux_h I__4482 (
            .O(N__26096),
            .I(N__26058));
    LocalMux I__4481 (
            .O(N__26093),
            .I(N__26058));
    LocalMux I__4480 (
            .O(N__26090),
            .I(N__26055));
    InMux I__4479 (
            .O(N__26089),
            .I(N__26050));
    InMux I__4478 (
            .O(N__26088),
            .I(N__26050));
    Span4Mux_h I__4477 (
            .O(N__26085),
            .I(N__26045));
    LocalMux I__4476 (
            .O(N__26076),
            .I(N__26045));
    InMux I__4475 (
            .O(N__26075),
            .I(N__26030));
    InMux I__4474 (
            .O(N__26074),
            .I(N__26030));
    InMux I__4473 (
            .O(N__26073),
            .I(N__26030));
    InMux I__4472 (
            .O(N__26072),
            .I(N__26030));
    InMux I__4471 (
            .O(N__26071),
            .I(N__26030));
    InMux I__4470 (
            .O(N__26070),
            .I(N__26030));
    InMux I__4469 (
            .O(N__26069),
            .I(N__26030));
    Odrv4 I__4468 (
            .O(N__26066),
            .I(n8272));
    Odrv4 I__4467 (
            .O(N__26063),
            .I(n8272));
    Odrv4 I__4466 (
            .O(N__26058),
            .I(n8272));
    Odrv4 I__4465 (
            .O(N__26055),
            .I(n8272));
    LocalMux I__4464 (
            .O(N__26050),
            .I(n8272));
    Odrv4 I__4463 (
            .O(N__26045),
            .I(n8272));
    LocalMux I__4462 (
            .O(N__26030),
            .I(n8272));
    CascadeMux I__4461 (
            .O(N__26015),
            .I(n4_adj_1264_cascade_));
    InMux I__4460 (
            .O(N__26012),
            .I(N__26009));
    LocalMux I__4459 (
            .O(N__26009),
            .I(N__26006));
    Odrv12 I__4458 (
            .O(N__26006),
            .I(n8055));
    CascadeMux I__4457 (
            .O(N__26003),
            .I(N__25999));
    InMux I__4456 (
            .O(N__26002),
            .I(N__25996));
    InMux I__4455 (
            .O(N__25999),
            .I(N__25992));
    LocalMux I__4454 (
            .O(N__25996),
            .I(N__25989));
    CascadeMux I__4453 (
            .O(N__25995),
            .I(N__25986));
    LocalMux I__4452 (
            .O(N__25992),
            .I(N__25983));
    Span4Mux_v I__4451 (
            .O(N__25989),
            .I(N__25980));
    InMux I__4450 (
            .O(N__25986),
            .I(N__25977));
    Span12Mux_v I__4449 (
            .O(N__25983),
            .I(N__25972));
    Sp12to4 I__4448 (
            .O(N__25980),
            .I(N__25972));
    LocalMux I__4447 (
            .O(N__25977),
            .I(buf_adcdata4_15));
    Odrv12 I__4446 (
            .O(N__25972),
            .I(buf_adcdata4_15));
    CascadeMux I__4445 (
            .O(N__25967),
            .I(N__25963));
    InMux I__4444 (
            .O(N__25966),
            .I(N__25957));
    InMux I__4443 (
            .O(N__25963),
            .I(N__25952));
    InMux I__4442 (
            .O(N__25962),
            .I(N__25952));
    InMux I__4441 (
            .O(N__25961),
            .I(N__25949));
    InMux I__4440 (
            .O(N__25960),
            .I(N__25946));
    LocalMux I__4439 (
            .O(N__25957),
            .I(N__25932));
    LocalMux I__4438 (
            .O(N__25952),
            .I(N__25932));
    LocalMux I__4437 (
            .O(N__25949),
            .I(N__25927));
    LocalMux I__4436 (
            .O(N__25946),
            .I(N__25927));
    InMux I__4435 (
            .O(N__25945),
            .I(N__25917));
    InMux I__4434 (
            .O(N__25944),
            .I(N__25910));
    InMux I__4433 (
            .O(N__25943),
            .I(N__25910));
    InMux I__4432 (
            .O(N__25942),
            .I(N__25910));
    InMux I__4431 (
            .O(N__25941),
            .I(N__25905));
    InMux I__4430 (
            .O(N__25940),
            .I(N__25905));
    InMux I__4429 (
            .O(N__25939),
            .I(N__25898));
    InMux I__4428 (
            .O(N__25938),
            .I(N__25898));
    InMux I__4427 (
            .O(N__25937),
            .I(N__25898));
    Span4Mux_v I__4426 (
            .O(N__25932),
            .I(N__25894));
    Span4Mux_h I__4425 (
            .O(N__25927),
            .I(N__25891));
    InMux I__4424 (
            .O(N__25926),
            .I(N__25884));
    InMux I__4423 (
            .O(N__25925),
            .I(N__25884));
    InMux I__4422 (
            .O(N__25924),
            .I(N__25884));
    InMux I__4421 (
            .O(N__25923),
            .I(N__25875));
    InMux I__4420 (
            .O(N__25922),
            .I(N__25875));
    InMux I__4419 (
            .O(N__25921),
            .I(N__25875));
    InMux I__4418 (
            .O(N__25920),
            .I(N__25872));
    LocalMux I__4417 (
            .O(N__25917),
            .I(N__25869));
    LocalMux I__4416 (
            .O(N__25910),
            .I(N__25866));
    LocalMux I__4415 (
            .O(N__25905),
            .I(N__25861));
    LocalMux I__4414 (
            .O(N__25898),
            .I(N__25861));
    InMux I__4413 (
            .O(N__25897),
            .I(N__25858));
    Span4Mux_h I__4412 (
            .O(N__25894),
            .I(N__25853));
    Span4Mux_v I__4411 (
            .O(N__25891),
            .I(N__25853));
    LocalMux I__4410 (
            .O(N__25884),
            .I(N__25850));
    InMux I__4409 (
            .O(N__25883),
            .I(N__25847));
    InMux I__4408 (
            .O(N__25882),
            .I(N__25844));
    LocalMux I__4407 (
            .O(N__25875),
            .I(N__25841));
    LocalMux I__4406 (
            .O(N__25872),
            .I(N__25836));
    Span4Mux_v I__4405 (
            .O(N__25869),
            .I(N__25836));
    Span4Mux_v I__4404 (
            .O(N__25866),
            .I(N__25833));
    Span4Mux_v I__4403 (
            .O(N__25861),
            .I(N__25830));
    LocalMux I__4402 (
            .O(N__25858),
            .I(N__25825));
    Span4Mux_v I__4401 (
            .O(N__25853),
            .I(N__25825));
    Span4Mux_v I__4400 (
            .O(N__25850),
            .I(N__25822));
    LocalMux I__4399 (
            .O(N__25847),
            .I(N__25811));
    LocalMux I__4398 (
            .O(N__25844),
            .I(N__25811));
    Span4Mux_h I__4397 (
            .O(N__25841),
            .I(N__25811));
    Span4Mux_h I__4396 (
            .O(N__25836),
            .I(N__25811));
    Span4Mux_v I__4395 (
            .O(N__25833),
            .I(N__25811));
    Span4Mux_h I__4394 (
            .O(N__25830),
            .I(N__25806));
    Span4Mux_v I__4393 (
            .O(N__25825),
            .I(N__25806));
    Odrv4 I__4392 (
            .O(N__25822),
            .I(n15144));
    Odrv4 I__4391 (
            .O(N__25811),
            .I(n15144));
    Odrv4 I__4390 (
            .O(N__25806),
            .I(n15144));
    CascadeMux I__4389 (
            .O(N__25799),
            .I(N__25795));
    InMux I__4388 (
            .O(N__25798),
            .I(N__25792));
    InMux I__4387 (
            .O(N__25795),
            .I(N__25789));
    LocalMux I__4386 (
            .O(N__25792),
            .I(N__25786));
    LocalMux I__4385 (
            .O(N__25789),
            .I(N__25783));
    Span4Mux_h I__4384 (
            .O(N__25786),
            .I(N__25780));
    Span4Mux_v I__4383 (
            .O(N__25783),
            .I(N__25776));
    Span4Mux_h I__4382 (
            .O(N__25780),
            .I(N__25773));
    InMux I__4381 (
            .O(N__25779),
            .I(N__25770));
    Span4Mux_h I__4380 (
            .O(N__25776),
            .I(N__25767));
    Span4Mux_h I__4379 (
            .O(N__25773),
            .I(N__25764));
    LocalMux I__4378 (
            .O(N__25770),
            .I(buf_adcdata4_17));
    Odrv4 I__4377 (
            .O(N__25767),
            .I(buf_adcdata4_17));
    Odrv4 I__4376 (
            .O(N__25764),
            .I(buf_adcdata4_17));
    InMux I__4375 (
            .O(N__25757),
            .I(N__25754));
    LocalMux I__4374 (
            .O(N__25754),
            .I(n71));
    CascadeMux I__4373 (
            .O(N__25751),
            .I(N__25748));
    InMux I__4372 (
            .O(N__25748),
            .I(N__25745));
    LocalMux I__4371 (
            .O(N__25745),
            .I(N__25742));
    Span4Mux_v I__4370 (
            .O(N__25742),
            .I(N__25737));
    InMux I__4369 (
            .O(N__25741),
            .I(N__25734));
    CascadeMux I__4368 (
            .O(N__25740),
            .I(N__25731));
    Span4Mux_h I__4367 (
            .O(N__25737),
            .I(N__25728));
    LocalMux I__4366 (
            .O(N__25734),
            .I(N__25725));
    InMux I__4365 (
            .O(N__25731),
            .I(N__25722));
    Odrv4 I__4364 (
            .O(N__25728),
            .I(cmd_rdadctmp_26_adj_1123));
    Odrv4 I__4363 (
            .O(N__25725),
            .I(cmd_rdadctmp_26_adj_1123));
    LocalMux I__4362 (
            .O(N__25722),
            .I(cmd_rdadctmp_26_adj_1123));
    CascadeMux I__4361 (
            .O(N__25715),
            .I(N__25712));
    InMux I__4360 (
            .O(N__25712),
            .I(N__25709));
    LocalMux I__4359 (
            .O(N__25709),
            .I(N__25704));
    CascadeMux I__4358 (
            .O(N__25708),
            .I(N__25701));
    CascadeMux I__4357 (
            .O(N__25707),
            .I(N__25698));
    Span4Mux_v I__4356 (
            .O(N__25704),
            .I(N__25695));
    InMux I__4355 (
            .O(N__25701),
            .I(N__25690));
    InMux I__4354 (
            .O(N__25698),
            .I(N__25690));
    Odrv4 I__4353 (
            .O(N__25695),
            .I(cmd_rdadctmp_27_adj_1085));
    LocalMux I__4352 (
            .O(N__25690),
            .I(cmd_rdadctmp_27_adj_1085));
    InMux I__4351 (
            .O(N__25685),
            .I(N__25682));
    LocalMux I__4350 (
            .O(N__25682),
            .I(N__25679));
    Span4Mux_v I__4349 (
            .O(N__25679),
            .I(N__25676));
    Sp12to4 I__4348 (
            .O(N__25676),
            .I(N__25673));
    Span12Mux_h I__4347 (
            .O(N__25673),
            .I(N__25670));
    Span12Mux_v I__4346 (
            .O(N__25670),
            .I(N__25665));
    InMux I__4345 (
            .O(N__25669),
            .I(N__25660));
    InMux I__4344 (
            .O(N__25668),
            .I(N__25660));
    Odrv12 I__4343 (
            .O(N__25665),
            .I(buf_adcdata3_23));
    LocalMux I__4342 (
            .O(N__25660),
            .I(buf_adcdata3_23));
    CascadeMux I__4341 (
            .O(N__25655),
            .I(N__25652));
    InMux I__4340 (
            .O(N__25652),
            .I(N__25648));
    CascadeMux I__4339 (
            .O(N__25651),
            .I(N__25644));
    LocalMux I__4338 (
            .O(N__25648),
            .I(N__25641));
    InMux I__4337 (
            .O(N__25647),
            .I(N__25638));
    InMux I__4336 (
            .O(N__25644),
            .I(N__25635));
    Span4Mux_v I__4335 (
            .O(N__25641),
            .I(N__25632));
    LocalMux I__4334 (
            .O(N__25638),
            .I(cmd_rdadctmp_27_adj_1122));
    LocalMux I__4333 (
            .O(N__25635),
            .I(cmd_rdadctmp_27_adj_1122));
    Odrv4 I__4332 (
            .O(N__25632),
            .I(cmd_rdadctmp_27_adj_1122));
    CascadeMux I__4331 (
            .O(N__25625),
            .I(N__25621));
    InMux I__4330 (
            .O(N__25624),
            .I(N__25618));
    InMux I__4329 (
            .O(N__25621),
            .I(N__25615));
    LocalMux I__4328 (
            .O(N__25618),
            .I(N__25612));
    LocalMux I__4327 (
            .O(N__25615),
            .I(N__25609));
    Span4Mux_v I__4326 (
            .O(N__25612),
            .I(N__25606));
    Span4Mux_v I__4325 (
            .O(N__25609),
            .I(N__25602));
    Span4Mux_v I__4324 (
            .O(N__25606),
            .I(N__25599));
    InMux I__4323 (
            .O(N__25605),
            .I(N__25596));
    Span4Mux_v I__4322 (
            .O(N__25602),
            .I(N__25593));
    Span4Mux_h I__4321 (
            .O(N__25599),
            .I(N__25588));
    LocalMux I__4320 (
            .O(N__25596),
            .I(N__25588));
    Odrv4 I__4319 (
            .O(N__25593),
            .I(cmd_rdadctmp_28_adj_1121));
    Odrv4 I__4318 (
            .O(N__25588),
            .I(cmd_rdadctmp_28_adj_1121));
    InMux I__4317 (
            .O(N__25583),
            .I(N__25576));
    InMux I__4316 (
            .O(N__25582),
            .I(N__25576));
    InMux I__4315 (
            .O(N__25581),
            .I(N__25573));
    LocalMux I__4314 (
            .O(N__25576),
            .I(N__25568));
    LocalMux I__4313 (
            .O(N__25573),
            .I(N__25565));
    CascadeMux I__4312 (
            .O(N__25572),
            .I(N__25562));
    CascadeMux I__4311 (
            .O(N__25571),
            .I(N__25559));
    Span4Mux_v I__4310 (
            .O(N__25568),
            .I(N__25555));
    Span4Mux_h I__4309 (
            .O(N__25565),
            .I(N__25552));
    InMux I__4308 (
            .O(N__25562),
            .I(N__25545));
    InMux I__4307 (
            .O(N__25559),
            .I(N__25545));
    InMux I__4306 (
            .O(N__25558),
            .I(N__25545));
    Span4Mux_h I__4305 (
            .O(N__25555),
            .I(N__25542));
    Span4Mux_h I__4304 (
            .O(N__25552),
            .I(N__25539));
    LocalMux I__4303 (
            .O(N__25545),
            .I(n15221));
    Odrv4 I__4302 (
            .O(N__25542),
            .I(n15221));
    Odrv4 I__4301 (
            .O(N__25539),
            .I(n15221));
    CascadeMux I__4300 (
            .O(N__25532),
            .I(n17_cascade_));
    CascadeMux I__4299 (
            .O(N__25529),
            .I(n8702_cascade_));
    InMux I__4298 (
            .O(N__25526),
            .I(N__25520));
    InMux I__4297 (
            .O(N__25525),
            .I(N__25520));
    LocalMux I__4296 (
            .O(N__25520),
            .I(bit_cnt_3));
    InMux I__4295 (
            .O(N__25517),
            .I(N__25508));
    InMux I__4294 (
            .O(N__25516),
            .I(N__25508));
    InMux I__4293 (
            .O(N__25515),
            .I(N__25508));
    LocalMux I__4292 (
            .O(N__25508),
            .I(bit_cnt_2));
    CascadeMux I__4291 (
            .O(N__25505),
            .I(N__25501));
    CascadeMux I__4290 (
            .O(N__25504),
            .I(N__25496));
    InMux I__4289 (
            .O(N__25501),
            .I(N__25490));
    InMux I__4288 (
            .O(N__25500),
            .I(N__25490));
    InMux I__4287 (
            .O(N__25499),
            .I(N__25485));
    InMux I__4286 (
            .O(N__25496),
            .I(N__25485));
    InMux I__4285 (
            .O(N__25495),
            .I(N__25482));
    LocalMux I__4284 (
            .O(N__25490),
            .I(N__25477));
    LocalMux I__4283 (
            .O(N__25485),
            .I(N__25477));
    LocalMux I__4282 (
            .O(N__25482),
            .I(N__25472));
    Span4Mux_v I__4281 (
            .O(N__25477),
            .I(N__25472));
    Odrv4 I__4280 (
            .O(N__25472),
            .I(bit_cnt_0));
    CascadeMux I__4279 (
            .O(N__25469),
            .I(n16524_cascade_));
    CascadeMux I__4278 (
            .O(N__25466),
            .I(n16527_cascade_));
    CascadeMux I__4277 (
            .O(N__25463),
            .I(n15565_cascade_));
    CascadeMux I__4276 (
            .O(N__25460),
            .I(n13_adj_1257_cascade_));
    CEMux I__4275 (
            .O(N__25457),
            .I(N__25454));
    LocalMux I__4274 (
            .O(N__25454),
            .I(N__25451));
    Span4Mux_v I__4273 (
            .O(N__25451),
            .I(N__25445));
    CEMux I__4272 (
            .O(N__25450),
            .I(N__25442));
    CEMux I__4271 (
            .O(N__25449),
            .I(N__25439));
    InMux I__4270 (
            .O(N__25448),
            .I(N__25436));
    Span4Mux_h I__4269 (
            .O(N__25445),
            .I(N__25427));
    LocalMux I__4268 (
            .O(N__25442),
            .I(N__25427));
    LocalMux I__4267 (
            .O(N__25439),
            .I(N__25427));
    LocalMux I__4266 (
            .O(N__25436),
            .I(N__25427));
    Span4Mux_h I__4265 (
            .O(N__25427),
            .I(N__25424));
    Odrv4 I__4264 (
            .O(N__25424),
            .I(n8823));
    InMux I__4263 (
            .O(N__25421),
            .I(N__25418));
    LocalMux I__4262 (
            .O(N__25418),
            .I(N__25414));
    InMux I__4261 (
            .O(N__25417),
            .I(N__25411));
    Odrv4 I__4260 (
            .O(N__25414),
            .I(n41));
    LocalMux I__4259 (
            .O(N__25411),
            .I(n41));
    InMux I__4258 (
            .O(N__25406),
            .I(N__25403));
    LocalMux I__4257 (
            .O(N__25403),
            .I(n13457));
    InMux I__4256 (
            .O(N__25400),
            .I(N__25394));
    InMux I__4255 (
            .O(N__25399),
            .I(N__25394));
    LocalMux I__4254 (
            .O(N__25394),
            .I(n13458));
    InMux I__4253 (
            .O(N__25391),
            .I(N__25388));
    LocalMux I__4252 (
            .O(N__25388),
            .I(N__25385));
    Span4Mux_v I__4251 (
            .O(N__25385),
            .I(N__25382));
    Span4Mux_h I__4250 (
            .O(N__25382),
            .I(N__25379));
    Span4Mux_h I__4249 (
            .O(N__25379),
            .I(N__25376));
    Span4Mux_v I__4248 (
            .O(N__25376),
            .I(N__25373));
    Odrv4 I__4247 (
            .O(N__25373),
            .I(buf_data4_13));
    InMux I__4246 (
            .O(N__25370),
            .I(N__25367));
    LocalMux I__4245 (
            .O(N__25367),
            .I(N__25364));
    Span4Mux_h I__4244 (
            .O(N__25364),
            .I(N__25361));
    Odrv4 I__4243 (
            .O(N__25361),
            .I(comm_buf_10_5));
    CEMux I__4242 (
            .O(N__25358),
            .I(N__25352));
    CEMux I__4241 (
            .O(N__25357),
            .I(N__25349));
    CEMux I__4240 (
            .O(N__25356),
            .I(N__25346));
    CEMux I__4239 (
            .O(N__25355),
            .I(N__25343));
    LocalMux I__4238 (
            .O(N__25352),
            .I(N__25340));
    LocalMux I__4237 (
            .O(N__25349),
            .I(N__25337));
    LocalMux I__4236 (
            .O(N__25346),
            .I(N__25334));
    LocalMux I__4235 (
            .O(N__25343),
            .I(N__25331));
    Span4Mux_v I__4234 (
            .O(N__25340),
            .I(N__25326));
    Span4Mux_v I__4233 (
            .O(N__25337),
            .I(N__25326));
    Odrv4 I__4232 (
            .O(N__25334),
            .I(n9045));
    Odrv12 I__4231 (
            .O(N__25331),
            .I(n9045));
    Odrv4 I__4230 (
            .O(N__25326),
            .I(n9045));
    SRMux I__4229 (
            .O(N__25319),
            .I(N__25314));
    SRMux I__4228 (
            .O(N__25318),
            .I(N__25310));
    SRMux I__4227 (
            .O(N__25317),
            .I(N__25307));
    LocalMux I__4226 (
            .O(N__25314),
            .I(N__25304));
    SRMux I__4225 (
            .O(N__25313),
            .I(N__25301));
    LocalMux I__4224 (
            .O(N__25310),
            .I(N__25298));
    LocalMux I__4223 (
            .O(N__25307),
            .I(N__25295));
    Span4Mux_h I__4222 (
            .O(N__25304),
            .I(N__25292));
    LocalMux I__4221 (
            .O(N__25301),
            .I(N__25289));
    Span4Mux_v I__4220 (
            .O(N__25298),
            .I(N__25284));
    Span4Mux_v I__4219 (
            .O(N__25295),
            .I(N__25284));
    Odrv4 I__4218 (
            .O(N__25292),
            .I(n10646));
    Odrv12 I__4217 (
            .O(N__25289),
            .I(n10646));
    Odrv4 I__4216 (
            .O(N__25284),
            .I(n10646));
    CascadeMux I__4215 (
            .O(N__25277),
            .I(n11_adj_1279_cascade_));
    CEMux I__4214 (
            .O(N__25274),
            .I(N__25271));
    LocalMux I__4213 (
            .O(N__25271),
            .I(N__25262));
    CEMux I__4212 (
            .O(N__25270),
            .I(N__25259));
    CEMux I__4211 (
            .O(N__25269),
            .I(N__25256));
    CEMux I__4210 (
            .O(N__25268),
            .I(N__25253));
    CEMux I__4209 (
            .O(N__25267),
            .I(N__25250));
    CEMux I__4208 (
            .O(N__25266),
            .I(N__25247));
    CEMux I__4207 (
            .O(N__25265),
            .I(N__25244));
    Span4Mux_v I__4206 (
            .O(N__25262),
            .I(N__25239));
    LocalMux I__4205 (
            .O(N__25259),
            .I(N__25239));
    LocalMux I__4204 (
            .O(N__25256),
            .I(N__25234));
    LocalMux I__4203 (
            .O(N__25253),
            .I(N__25234));
    LocalMux I__4202 (
            .O(N__25250),
            .I(N__25231));
    LocalMux I__4201 (
            .O(N__25247),
            .I(N__25228));
    LocalMux I__4200 (
            .O(N__25244),
            .I(N__25225));
    Span4Mux_h I__4199 (
            .O(N__25239),
            .I(N__25221));
    Span4Mux_v I__4198 (
            .O(N__25234),
            .I(N__25218));
    Span4Mux_v I__4197 (
            .O(N__25231),
            .I(N__25213));
    Span4Mux_h I__4196 (
            .O(N__25228),
            .I(N__25213));
    Span4Mux_h I__4195 (
            .O(N__25225),
            .I(N__25210));
    InMux I__4194 (
            .O(N__25224),
            .I(N__25207));
    Odrv4 I__4193 (
            .O(N__25221),
            .I(n8654));
    Odrv4 I__4192 (
            .O(N__25218),
            .I(n8654));
    Odrv4 I__4191 (
            .O(N__25213),
            .I(n8654));
    Odrv4 I__4190 (
            .O(N__25210),
            .I(n8654));
    LocalMux I__4189 (
            .O(N__25207),
            .I(n8654));
    CascadeMux I__4188 (
            .O(N__25196),
            .I(N__25193));
    InMux I__4187 (
            .O(N__25193),
            .I(N__25189));
    InMux I__4186 (
            .O(N__25192),
            .I(N__25186));
    LocalMux I__4185 (
            .O(N__25189),
            .I(N__25183));
    LocalMux I__4184 (
            .O(N__25186),
            .I(N__25180));
    Odrv4 I__4183 (
            .O(N__25183),
            .I(n5));
    Odrv12 I__4182 (
            .O(N__25180),
            .I(n5));
    CEMux I__4181 (
            .O(N__25175),
            .I(N__25172));
    LocalMux I__4180 (
            .O(N__25172),
            .I(N__25169));
    Odrv12 I__4179 (
            .O(N__25169),
            .I(n8763));
    InMux I__4178 (
            .O(N__25166),
            .I(N__25162));
    InMux I__4177 (
            .O(N__25165),
            .I(N__25159));
    LocalMux I__4176 (
            .O(N__25162),
            .I(n13470));
    LocalMux I__4175 (
            .O(N__25159),
            .I(n13470));
    InMux I__4174 (
            .O(N__25154),
            .I(N__25151));
    LocalMux I__4173 (
            .O(N__25151),
            .I(n13497));
    CascadeMux I__4172 (
            .O(N__25148),
            .I(n13497_cascade_));
    CascadeMux I__4171 (
            .O(N__25145),
            .I(n9045_cascade_));
    CascadeMux I__4170 (
            .O(N__25142),
            .I(N__25139));
    InMux I__4169 (
            .O(N__25139),
            .I(N__25136));
    LocalMux I__4168 (
            .O(N__25136),
            .I(N__25133));
    Span4Mux_h I__4167 (
            .O(N__25133),
            .I(N__25130));
    Odrv4 I__4166 (
            .O(N__25130),
            .I(comm_buf_11_6));
    InMux I__4165 (
            .O(N__25127),
            .I(N__25124));
    LocalMux I__4164 (
            .O(N__25124),
            .I(N__25121));
    Span4Mux_h I__4163 (
            .O(N__25121),
            .I(N__25118));
    Odrv4 I__4162 (
            .O(N__25118),
            .I(n16488));
    CascadeMux I__4161 (
            .O(N__25115),
            .I(N__25112));
    InMux I__4160 (
            .O(N__25112),
            .I(N__25109));
    LocalMux I__4159 (
            .O(N__25109),
            .I(N__25106));
    Span4Mux_v I__4158 (
            .O(N__25106),
            .I(N__25103));
    Span4Mux_h I__4157 (
            .O(N__25103),
            .I(N__25100));
    Span4Mux_h I__4156 (
            .O(N__25100),
            .I(N__25097));
    Odrv4 I__4155 (
            .O(N__25097),
            .I(buf_data4_14));
    InMux I__4154 (
            .O(N__25094),
            .I(N__25091));
    LocalMux I__4153 (
            .O(N__25091),
            .I(comm_buf_10_6));
    CascadeMux I__4152 (
            .O(N__25088),
            .I(n13457_cascade_));
    CascadeMux I__4151 (
            .O(N__25085),
            .I(n15161_cascade_));
    CEMux I__4150 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__4149 (
            .O(N__25079),
            .I(N__25076));
    Span4Mux_h I__4148 (
            .O(N__25076),
            .I(N__25073));
    Odrv4 I__4147 (
            .O(N__25073),
            .I(n8997));
    CascadeMux I__4146 (
            .O(N__25070),
            .I(n8997_cascade_));
    SRMux I__4145 (
            .O(N__25067),
            .I(N__25064));
    LocalMux I__4144 (
            .O(N__25064),
            .I(n10632));
    InMux I__4143 (
            .O(N__25061),
            .I(N__25058));
    LocalMux I__4142 (
            .O(N__25058),
            .I(N__25055));
    Span4Mux_v I__4141 (
            .O(N__25055),
            .I(N__25052));
    Span4Mux_h I__4140 (
            .O(N__25052),
            .I(N__25049));
    Span4Mux_h I__4139 (
            .O(N__25049),
            .I(N__25046));
    Odrv4 I__4138 (
            .O(N__25046),
            .I(buf_data4_16));
    InMux I__4137 (
            .O(N__25043),
            .I(N__25040));
    LocalMux I__4136 (
            .O(N__25040),
            .I(N__25037));
    Span4Mux_h I__4135 (
            .O(N__25037),
            .I(N__25034));
    Odrv4 I__4134 (
            .O(N__25034),
            .I(comm_buf_9_0));
    CEMux I__4133 (
            .O(N__25031),
            .I(N__25026));
    CEMux I__4132 (
            .O(N__25030),
            .I(N__25023));
    InMux I__4131 (
            .O(N__25029),
            .I(N__25020));
    LocalMux I__4130 (
            .O(N__25026),
            .I(n9027));
    LocalMux I__4129 (
            .O(N__25023),
            .I(n9027));
    LocalMux I__4128 (
            .O(N__25020),
            .I(n9027));
    SRMux I__4127 (
            .O(N__25013),
            .I(N__25009));
    SRMux I__4126 (
            .O(N__25012),
            .I(N__25006));
    LocalMux I__4125 (
            .O(N__25009),
            .I(N__25003));
    LocalMux I__4124 (
            .O(N__25006),
            .I(N__24998));
    Span4Mux_h I__4123 (
            .O(N__25003),
            .I(N__24998));
    Odrv4 I__4122 (
            .O(N__24998),
            .I(n10639));
    CascadeMux I__4121 (
            .O(N__24995),
            .I(N__24992));
    InMux I__4120 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__4119 (
            .O(N__24989),
            .I(N__24986));
    Span4Mux_h I__4118 (
            .O(N__24986),
            .I(N__24983));
    Odrv4 I__4117 (
            .O(N__24983),
            .I(comm_buf_11_1));
    InMux I__4116 (
            .O(N__24980),
            .I(N__24977));
    LocalMux I__4115 (
            .O(N__24977),
            .I(N__24974));
    Span4Mux_v I__4114 (
            .O(N__24974),
            .I(N__24971));
    Span4Mux_h I__4113 (
            .O(N__24971),
            .I(N__24968));
    Odrv4 I__4112 (
            .O(N__24968),
            .I(n16422));
    InMux I__4111 (
            .O(N__24965),
            .I(N__24962));
    LocalMux I__4110 (
            .O(N__24962),
            .I(N__24959));
    Span4Mux_h I__4109 (
            .O(N__24959),
            .I(N__24956));
    Span4Mux_v I__4108 (
            .O(N__24956),
            .I(N__24953));
    Span4Mux_v I__4107 (
            .O(N__24953),
            .I(N__24950));
    Span4Mux_h I__4106 (
            .O(N__24950),
            .I(N__24947));
    Span4Mux_h I__4105 (
            .O(N__24947),
            .I(N__24944));
    Odrv4 I__4104 (
            .O(N__24944),
            .I(buf_data4_9));
    InMux I__4103 (
            .O(N__24941),
            .I(N__24938));
    LocalMux I__4102 (
            .O(N__24938),
            .I(comm_buf_10_1));
    InMux I__4101 (
            .O(N__24935),
            .I(N__24929));
    InMux I__4100 (
            .O(N__24934),
            .I(N__24929));
    LocalMux I__4099 (
            .O(N__24929),
            .I(N__24925));
    InMux I__4098 (
            .O(N__24928),
            .I(N__24922));
    Span4Mux_h I__4097 (
            .O(N__24925),
            .I(N__24919));
    LocalMux I__4096 (
            .O(N__24922),
            .I(N__24916));
    Span4Mux_v I__4095 (
            .O(N__24919),
            .I(N__24913));
    Span12Mux_v I__4094 (
            .O(N__24916),
            .I(N__24910));
    Odrv4 I__4093 (
            .O(N__24913),
            .I(comm_tx_buf_2));
    Odrv12 I__4092 (
            .O(N__24910),
            .I(comm_tx_buf_2));
    SRMux I__4091 (
            .O(N__24905),
            .I(N__24902));
    LocalMux I__4090 (
            .O(N__24902),
            .I(N__24899));
    Span4Mux_h I__4089 (
            .O(N__24899),
            .I(N__24896));
    Sp12to4 I__4088 (
            .O(N__24896),
            .I(N__24893));
    Odrv12 I__4087 (
            .O(N__24893),
            .I(\comm_spi.data_tx_7__N_810 ));
    InMux I__4086 (
            .O(N__24890),
            .I(N__24886));
    InMux I__4085 (
            .O(N__24889),
            .I(N__24883));
    LocalMux I__4084 (
            .O(N__24886),
            .I(\comm_spi.n16905 ));
    LocalMux I__4083 (
            .O(N__24883),
            .I(\comm_spi.n16905 ));
    InMux I__4082 (
            .O(N__24878),
            .I(N__24875));
    LocalMux I__4081 (
            .O(N__24875),
            .I(N__24872));
    Span4Mux_v I__4080 (
            .O(N__24872),
            .I(N__24868));
    InMux I__4079 (
            .O(N__24871),
            .I(N__24865));
    Span4Mux_h I__4078 (
            .O(N__24868),
            .I(N__24862));
    LocalMux I__4077 (
            .O(N__24865),
            .I(N__24859));
    Odrv4 I__4076 (
            .O(N__24862),
            .I(\comm_spi.n10463 ));
    Odrv4 I__4075 (
            .O(N__24859),
            .I(\comm_spi.n10463 ));
    InMux I__4074 (
            .O(N__24854),
            .I(N__24850));
    InMux I__4073 (
            .O(N__24853),
            .I(N__24847));
    LocalMux I__4072 (
            .O(N__24850),
            .I(\comm_spi.n10464 ));
    LocalMux I__4071 (
            .O(N__24847),
            .I(\comm_spi.n10464 ));
    InMux I__4070 (
            .O(N__24842),
            .I(N__24839));
    LocalMux I__4069 (
            .O(N__24839),
            .I(N__24836));
    Span4Mux_v I__4068 (
            .O(N__24836),
            .I(N__24833));
    Span4Mux_h I__4067 (
            .O(N__24833),
            .I(N__24830));
    Span4Mux_h I__4066 (
            .O(N__24830),
            .I(N__24827));
    Odrv4 I__4065 (
            .O(N__24827),
            .I(buf_data4_21));
    InMux I__4064 (
            .O(N__24824),
            .I(N__24821));
    LocalMux I__4063 (
            .O(N__24821),
            .I(N__24818));
    Span4Mux_h I__4062 (
            .O(N__24818),
            .I(N__24815));
    Odrv4 I__4061 (
            .O(N__24815),
            .I(comm_buf_9_5));
    InMux I__4060 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__4059 (
            .O(N__24809),
            .I(N__24806));
    Span4Mux_h I__4058 (
            .O(N__24806),
            .I(N__24803));
    Span4Mux_h I__4057 (
            .O(N__24803),
            .I(N__24800));
    Span4Mux_v I__4056 (
            .O(N__24800),
            .I(N__24797));
    Odrv4 I__4055 (
            .O(N__24797),
            .I(buf_data4_22));
    CascadeMux I__4054 (
            .O(N__24794),
            .I(N__24791));
    InMux I__4053 (
            .O(N__24791),
            .I(N__24788));
    LocalMux I__4052 (
            .O(N__24788),
            .I(N__24785));
    Odrv12 I__4051 (
            .O(N__24785),
            .I(comm_buf_9_6));
    InMux I__4050 (
            .O(N__24782),
            .I(N__24779));
    LocalMux I__4049 (
            .O(N__24779),
            .I(N__24776));
    Span4Mux_v I__4048 (
            .O(N__24776),
            .I(N__24773));
    Span4Mux_h I__4047 (
            .O(N__24773),
            .I(N__24770));
    Span4Mux_h I__4046 (
            .O(N__24770),
            .I(N__24767));
    Odrv4 I__4045 (
            .O(N__24767),
            .I(buf_data4_23));
    InMux I__4044 (
            .O(N__24764),
            .I(N__24761));
    LocalMux I__4043 (
            .O(N__24761),
            .I(N__24758));
    Odrv12 I__4042 (
            .O(N__24758),
            .I(comm_buf_9_7));
    InMux I__4041 (
            .O(N__24755),
            .I(N__24752));
    LocalMux I__4040 (
            .O(N__24752),
            .I(N__24749));
    Span4Mux_h I__4039 (
            .O(N__24749),
            .I(N__24746));
    Span4Mux_h I__4038 (
            .O(N__24746),
            .I(N__24743));
    Span4Mux_h I__4037 (
            .O(N__24743),
            .I(N__24740));
    Odrv4 I__4036 (
            .O(N__24740),
            .I(buf_data4_18));
    InMux I__4035 (
            .O(N__24737),
            .I(N__24734));
    LocalMux I__4034 (
            .O(N__24734),
            .I(N__24731));
    Span4Mux_h I__4033 (
            .O(N__24731),
            .I(N__24728));
    Odrv4 I__4032 (
            .O(N__24728),
            .I(comm_buf_9_2));
    InMux I__4031 (
            .O(N__24725),
            .I(N__24722));
    LocalMux I__4030 (
            .O(N__24722),
            .I(N__24719));
    Span4Mux_v I__4029 (
            .O(N__24719),
            .I(N__24716));
    Span4Mux_h I__4028 (
            .O(N__24716),
            .I(N__24713));
    Span4Mux_h I__4027 (
            .O(N__24713),
            .I(N__24710));
    Odrv4 I__4026 (
            .O(N__24710),
            .I(buf_data4_17));
    CascadeMux I__4025 (
            .O(N__24707),
            .I(N__24704));
    InMux I__4024 (
            .O(N__24704),
            .I(N__24701));
    LocalMux I__4023 (
            .O(N__24701),
            .I(N__24698));
    Span4Mux_v I__4022 (
            .O(N__24698),
            .I(N__24695));
    Odrv4 I__4021 (
            .O(N__24695),
            .I(comm_buf_9_1));
    CascadeMux I__4020 (
            .O(N__24692),
            .I(N__24688));
    InMux I__4019 (
            .O(N__24691),
            .I(N__24685));
    InMux I__4018 (
            .O(N__24688),
            .I(N__24682));
    LocalMux I__4017 (
            .O(N__24685),
            .I(\ADC_VAC4.bit_cnt_5 ));
    LocalMux I__4016 (
            .O(N__24682),
            .I(\ADC_VAC4.bit_cnt_5 ));
    InMux I__4015 (
            .O(N__24677),
            .I(N__24674));
    LocalMux I__4014 (
            .O(N__24674),
            .I(\ADC_VAC4.n15354 ));
    CascadeMux I__4013 (
            .O(N__24671),
            .I(\ADC_VAC4.n15619_cascade_ ));
    CEMux I__4012 (
            .O(N__24668),
            .I(N__24665));
    LocalMux I__4011 (
            .O(N__24665),
            .I(\ADC_VAC4.n9631 ));
    CascadeMux I__4010 (
            .O(N__24662),
            .I(\ADC_VAC4.n9631_cascade_ ));
    SRMux I__4009 (
            .O(N__24659),
            .I(N__24656));
    LocalMux I__4008 (
            .O(N__24656),
            .I(\ADC_VAC4.n10783 ));
    InMux I__4007 (
            .O(N__24653),
            .I(N__24649));
    CascadeMux I__4006 (
            .O(N__24652),
            .I(N__24646));
    LocalMux I__4005 (
            .O(N__24649),
            .I(N__24643));
    InMux I__4004 (
            .O(N__24646),
            .I(N__24640));
    Span4Mux_v I__4003 (
            .O(N__24643),
            .I(N__24636));
    LocalMux I__4002 (
            .O(N__24640),
            .I(N__24633));
    InMux I__4001 (
            .O(N__24639),
            .I(N__24630));
    Sp12to4 I__4000 (
            .O(N__24636),
            .I(N__24627));
    Span4Mux_h I__3999 (
            .O(N__24633),
            .I(N__24624));
    LocalMux I__3998 (
            .O(N__24630),
            .I(buf_adcdata4_20));
    Odrv12 I__3997 (
            .O(N__24627),
            .I(buf_adcdata4_20));
    Odrv4 I__3996 (
            .O(N__24624),
            .I(buf_adcdata4_20));
    CascadeMux I__3995 (
            .O(N__24617),
            .I(\comm_spi.n16905_cascade_ ));
    SRMux I__3994 (
            .O(N__24614),
            .I(N__24611));
    LocalMux I__3993 (
            .O(N__24611),
            .I(N__24608));
    Span4Mux_v I__3992 (
            .O(N__24608),
            .I(N__24605));
    Odrv4 I__3991 (
            .O(N__24605),
            .I(\comm_spi.data_tx_7__N_809 ));
    InMux I__3990 (
            .O(N__24602),
            .I(N__24599));
    LocalMux I__3989 (
            .O(N__24599),
            .I(N__24596));
    Span4Mux_v I__3988 (
            .O(N__24596),
            .I(N__24592));
    CascadeMux I__3987 (
            .O(N__24595),
            .I(N__24589));
    Span4Mux_h I__3986 (
            .O(N__24592),
            .I(N__24586));
    InMux I__3985 (
            .O(N__24589),
            .I(N__24583));
    Span4Mux_h I__3984 (
            .O(N__24586),
            .I(N__24580));
    LocalMux I__3983 (
            .O(N__24583),
            .I(buf_adcdata1_9));
    Odrv4 I__3982 (
            .O(N__24580),
            .I(buf_adcdata1_9));
    CascadeMux I__3981 (
            .O(N__24575),
            .I(N__24570));
    InMux I__3980 (
            .O(N__24574),
            .I(N__24565));
    InMux I__3979 (
            .O(N__24573),
            .I(N__24565));
    InMux I__3978 (
            .O(N__24570),
            .I(N__24562));
    LocalMux I__3977 (
            .O(N__24565),
            .I(cmd_rdadctmp_17));
    LocalMux I__3976 (
            .O(N__24562),
            .I(cmd_rdadctmp_17));
    CascadeMux I__3975 (
            .O(N__24557),
            .I(N__24553));
    InMux I__3974 (
            .O(N__24556),
            .I(N__24547));
    InMux I__3973 (
            .O(N__24553),
            .I(N__24547));
    InMux I__3972 (
            .O(N__24552),
            .I(N__24544));
    LocalMux I__3971 (
            .O(N__24547),
            .I(cmd_rdadctmp_19));
    LocalMux I__3970 (
            .O(N__24544),
            .I(cmd_rdadctmp_19));
    InMux I__3969 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__3968 (
            .O(N__24536),
            .I(N__24533));
    Span4Mux_v I__3967 (
            .O(N__24533),
            .I(N__24529));
    CascadeMux I__3966 (
            .O(N__24532),
            .I(N__24526));
    Span4Mux_h I__3965 (
            .O(N__24529),
            .I(N__24523));
    InMux I__3964 (
            .O(N__24526),
            .I(N__24520));
    Span4Mux_h I__3963 (
            .O(N__24523),
            .I(N__24517));
    LocalMux I__3962 (
            .O(N__24520),
            .I(buf_adcdata1_11));
    Odrv4 I__3961 (
            .O(N__24517),
            .I(buf_adcdata1_11));
    InMux I__3960 (
            .O(N__24512),
            .I(N__24508));
    InMux I__3959 (
            .O(N__24511),
            .I(N__24505));
    LocalMux I__3958 (
            .O(N__24508),
            .I(N__24502));
    LocalMux I__3957 (
            .O(N__24505),
            .I(N__24498));
    Span4Mux_h I__3956 (
            .O(N__24502),
            .I(N__24495));
    InMux I__3955 (
            .O(N__24501),
            .I(N__24492));
    Span12Mux_s10_v I__3954 (
            .O(N__24498),
            .I(N__24489));
    Span4Mux_v I__3953 (
            .O(N__24495),
            .I(N__24486));
    LocalMux I__3952 (
            .O(N__24492),
            .I(buf_adcdata3_8));
    Odrv12 I__3951 (
            .O(N__24489),
            .I(buf_adcdata3_8));
    Odrv4 I__3950 (
            .O(N__24486),
            .I(buf_adcdata3_8));
    InMux I__3949 (
            .O(N__24479),
            .I(N__24475));
    InMux I__3948 (
            .O(N__24478),
            .I(N__24472));
    LocalMux I__3947 (
            .O(N__24475),
            .I(\ADC_VAC4.bit_cnt_4 ));
    LocalMux I__3946 (
            .O(N__24472),
            .I(\ADC_VAC4.bit_cnt_4 ));
    InMux I__3945 (
            .O(N__24467),
            .I(N__24463));
    InMux I__3944 (
            .O(N__24466),
            .I(N__24460));
    LocalMux I__3943 (
            .O(N__24463),
            .I(\ADC_VAC4.bit_cnt_3 ));
    LocalMux I__3942 (
            .O(N__24460),
            .I(\ADC_VAC4.bit_cnt_3 ));
    CascadeMux I__3941 (
            .O(N__24455),
            .I(N__24451));
    InMux I__3940 (
            .O(N__24454),
            .I(N__24448));
    InMux I__3939 (
            .O(N__24451),
            .I(N__24445));
    LocalMux I__3938 (
            .O(N__24448),
            .I(\ADC_VAC4.bit_cnt_1 ));
    LocalMux I__3937 (
            .O(N__24445),
            .I(\ADC_VAC4.bit_cnt_1 ));
    InMux I__3936 (
            .O(N__24440),
            .I(N__24436));
    InMux I__3935 (
            .O(N__24439),
            .I(N__24433));
    LocalMux I__3934 (
            .O(N__24436),
            .I(\ADC_VAC4.bit_cnt_2 ));
    LocalMux I__3933 (
            .O(N__24433),
            .I(\ADC_VAC4.bit_cnt_2 ));
    InMux I__3932 (
            .O(N__24428),
            .I(N__24424));
    InMux I__3931 (
            .O(N__24427),
            .I(N__24421));
    LocalMux I__3930 (
            .O(N__24424),
            .I(N__24418));
    LocalMux I__3929 (
            .O(N__24421),
            .I(\ADC_VAC4.bit_cnt_6 ));
    Odrv4 I__3928 (
            .O(N__24418),
            .I(\ADC_VAC4.bit_cnt_6 ));
    InMux I__3927 (
            .O(N__24413),
            .I(N__24409));
    InMux I__3926 (
            .O(N__24412),
            .I(N__24406));
    LocalMux I__3925 (
            .O(N__24409),
            .I(\ADC_VAC4.bit_cnt_0 ));
    LocalMux I__3924 (
            .O(N__24406),
            .I(\ADC_VAC4.bit_cnt_0 ));
    CascadeMux I__3923 (
            .O(N__24401),
            .I(\ADC_VAC4.n15330_cascade_ ));
    InMux I__3922 (
            .O(N__24398),
            .I(N__24394));
    InMux I__3921 (
            .O(N__24397),
            .I(N__24391));
    LocalMux I__3920 (
            .O(N__24394),
            .I(\ADC_VAC4.bit_cnt_7 ));
    LocalMux I__3919 (
            .O(N__24391),
            .I(\ADC_VAC4.bit_cnt_7 ));
    InMux I__3918 (
            .O(N__24386),
            .I(N__24383));
    LocalMux I__3917 (
            .O(N__24383),
            .I(N__24380));
    Odrv4 I__3916 (
            .O(N__24380),
            .I(n69));
    CascadeMux I__3915 (
            .O(N__24377),
            .I(N__24373));
    CascadeMux I__3914 (
            .O(N__24376),
            .I(N__24370));
    InMux I__3913 (
            .O(N__24373),
            .I(N__24365));
    InMux I__3912 (
            .O(N__24370),
            .I(N__24365));
    LocalMux I__3911 (
            .O(N__24365),
            .I(buf_control_0));
    InMux I__3910 (
            .O(N__24362),
            .I(N__24359));
    LocalMux I__3909 (
            .O(N__24359),
            .I(N__24356));
    Span12Mux_h I__3908 (
            .O(N__24356),
            .I(N__24353));
    Odrv12 I__3907 (
            .O(N__24353),
            .I(buf_data2_8));
    InMux I__3906 (
            .O(N__24350),
            .I(N__24347));
    LocalMux I__3905 (
            .O(N__24347),
            .I(N__24343));
    CascadeMux I__3904 (
            .O(N__24346),
            .I(N__24340));
    Span4Mux_h I__3903 (
            .O(N__24343),
            .I(N__24337));
    InMux I__3902 (
            .O(N__24340),
            .I(N__24333));
    Span4Mux_h I__3901 (
            .O(N__24337),
            .I(N__24330));
    CascadeMux I__3900 (
            .O(N__24336),
            .I(N__24327));
    LocalMux I__3899 (
            .O(N__24333),
            .I(N__24324));
    Sp12to4 I__3898 (
            .O(N__24330),
            .I(N__24321));
    InMux I__3897 (
            .O(N__24327),
            .I(N__24318));
    Span4Mux_h I__3896 (
            .O(N__24324),
            .I(N__24315));
    Span12Mux_v I__3895 (
            .O(N__24321),
            .I(N__24312));
    LocalMux I__3894 (
            .O(N__24318),
            .I(buf_adcdata4_8));
    Odrv4 I__3893 (
            .O(N__24315),
            .I(buf_adcdata4_8));
    Odrv12 I__3892 (
            .O(N__24312),
            .I(buf_adcdata4_8));
    InMux I__3891 (
            .O(N__24305),
            .I(N__24302));
    LocalMux I__3890 (
            .O(N__24302),
            .I(N__24299));
    Span4Mux_v I__3889 (
            .O(N__24299),
            .I(N__24296));
    Span4Mux_h I__3888 (
            .O(N__24296),
            .I(N__24293));
    Odrv4 I__3887 (
            .O(N__24293),
            .I(n4064));
    CascadeMux I__3886 (
            .O(N__24290),
            .I(N__24287));
    InMux I__3885 (
            .O(N__24287),
            .I(N__24283));
    CascadeMux I__3884 (
            .O(N__24286),
            .I(N__24280));
    LocalMux I__3883 (
            .O(N__24283),
            .I(N__24277));
    InMux I__3882 (
            .O(N__24280),
            .I(N__24274));
    Odrv12 I__3881 (
            .O(N__24277),
            .I(cmd_rdadctmp_5_adj_1107));
    LocalMux I__3880 (
            .O(N__24274),
            .I(cmd_rdadctmp_5_adj_1107));
    InMux I__3879 (
            .O(N__24269),
            .I(N__24266));
    LocalMux I__3878 (
            .O(N__24266),
            .I(N__24263));
    Span4Mux_h I__3877 (
            .O(N__24263),
            .I(N__24259));
    InMux I__3876 (
            .O(N__24262),
            .I(N__24256));
    Odrv4 I__3875 (
            .O(N__24259),
            .I(cmd_rdadctmp_6_adj_1106));
    LocalMux I__3874 (
            .O(N__24256),
            .I(cmd_rdadctmp_6_adj_1106));
    CascadeMux I__3873 (
            .O(N__24251),
            .I(N__24248));
    InMux I__3872 (
            .O(N__24248),
            .I(N__24245));
    LocalMux I__3871 (
            .O(N__24245),
            .I(N__24241));
    InMux I__3870 (
            .O(N__24244),
            .I(N__24238));
    Span4Mux_h I__3869 (
            .O(N__24241),
            .I(N__24234));
    LocalMux I__3868 (
            .O(N__24238),
            .I(N__24231));
    InMux I__3867 (
            .O(N__24237),
            .I(N__24228));
    Odrv4 I__3866 (
            .O(N__24234),
            .I(cmd_rdadctmp_28_adj_1084));
    Odrv4 I__3865 (
            .O(N__24231),
            .I(cmd_rdadctmp_28_adj_1084));
    LocalMux I__3864 (
            .O(N__24228),
            .I(cmd_rdadctmp_28_adj_1084));
    CascadeMux I__3863 (
            .O(N__24221),
            .I(n16503_cascade_));
    InMux I__3862 (
            .O(N__24218),
            .I(N__24215));
    LocalMux I__3861 (
            .O(N__24215),
            .I(n4_adj_1280));
    CascadeMux I__3860 (
            .O(N__24212),
            .I(n8047_cascade_));
    SRMux I__3859 (
            .O(N__24209),
            .I(N__24206));
    LocalMux I__3858 (
            .O(N__24206),
            .I(N__24202));
    SRMux I__3857 (
            .O(N__24205),
            .I(N__24199));
    Span4Mux_h I__3856 (
            .O(N__24202),
            .I(N__24194));
    LocalMux I__3855 (
            .O(N__24199),
            .I(N__24194));
    Span4Mux_h I__3854 (
            .O(N__24194),
            .I(N__24189));
    SRMux I__3853 (
            .O(N__24193),
            .I(N__24183));
    SRMux I__3852 (
            .O(N__24192),
            .I(N__24180));
    Span4Mux_h I__3851 (
            .O(N__24189),
            .I(N__24177));
    SRMux I__3850 (
            .O(N__24188),
            .I(N__24174));
    SRMux I__3849 (
            .O(N__24187),
            .I(N__24171));
    SRMux I__3848 (
            .O(N__24186),
            .I(N__24168));
    LocalMux I__3847 (
            .O(N__24183),
            .I(n10576));
    LocalMux I__3846 (
            .O(N__24180),
            .I(n10576));
    Odrv4 I__3845 (
            .O(N__24177),
            .I(n10576));
    LocalMux I__3844 (
            .O(N__24174),
            .I(n10576));
    LocalMux I__3843 (
            .O(N__24171),
            .I(n10576));
    LocalMux I__3842 (
            .O(N__24168),
            .I(n10576));
    InMux I__3841 (
            .O(N__24155),
            .I(N__24151));
    CascadeMux I__3840 (
            .O(N__24154),
            .I(N__24148));
    LocalMux I__3839 (
            .O(N__24151),
            .I(N__24145));
    InMux I__3838 (
            .O(N__24148),
            .I(N__24141));
    Span4Mux_h I__3837 (
            .O(N__24145),
            .I(N__24138));
    InMux I__3836 (
            .O(N__24144),
            .I(N__24135));
    LocalMux I__3835 (
            .O(N__24141),
            .I(cmd_rdadctmp_9));
    Odrv4 I__3834 (
            .O(N__24138),
            .I(cmd_rdadctmp_9));
    LocalMux I__3833 (
            .O(N__24135),
            .I(cmd_rdadctmp_9));
    CascadeMux I__3832 (
            .O(N__24128),
            .I(N__24124));
    CascadeMux I__3831 (
            .O(N__24127),
            .I(N__24121));
    InMux I__3830 (
            .O(N__24124),
            .I(N__24116));
    InMux I__3829 (
            .O(N__24121),
            .I(N__24116));
    LocalMux I__3828 (
            .O(N__24116),
            .I(buf_control_3));
    InMux I__3827 (
            .O(N__24113),
            .I(N__24110));
    LocalMux I__3826 (
            .O(N__24110),
            .I(n69_adj_1029));
    InMux I__3825 (
            .O(N__24107),
            .I(N__24104));
    LocalMux I__3824 (
            .O(N__24104),
            .I(N__24100));
    CascadeMux I__3823 (
            .O(N__24103),
            .I(N__24097));
    Span4Mux_v I__3822 (
            .O(N__24100),
            .I(N__24093));
    InMux I__3821 (
            .O(N__24097),
            .I(N__24090));
    InMux I__3820 (
            .O(N__24096),
            .I(N__24087));
    Sp12to4 I__3819 (
            .O(N__24093),
            .I(N__24084));
    LocalMux I__3818 (
            .O(N__24090),
            .I(N__24081));
    LocalMux I__3817 (
            .O(N__24087),
            .I(buf_adcdata4_14));
    Odrv12 I__3816 (
            .O(N__24084),
            .I(buf_adcdata4_14));
    Odrv4 I__3815 (
            .O(N__24081),
            .I(buf_adcdata4_14));
    InMux I__3814 (
            .O(N__24074),
            .I(N__24070));
    InMux I__3813 (
            .O(N__24073),
            .I(N__24067));
    LocalMux I__3812 (
            .O(N__24070),
            .I(N__24064));
    LocalMux I__3811 (
            .O(N__24067),
            .I(N__24061));
    Span4Mux_h I__3810 (
            .O(N__24064),
            .I(N__24057));
    Span12Mux_v I__3809 (
            .O(N__24061),
            .I(N__24054));
    InMux I__3808 (
            .O(N__24060),
            .I(N__24051));
    Span4Mux_v I__3807 (
            .O(N__24057),
            .I(N__24048));
    Span12Mux_h I__3806 (
            .O(N__24054),
            .I(N__24045));
    LocalMux I__3805 (
            .O(N__24051),
            .I(buf_adcdata3_20));
    Odrv4 I__3804 (
            .O(N__24048),
            .I(buf_adcdata3_20));
    Odrv12 I__3803 (
            .O(N__24045),
            .I(buf_adcdata3_20));
    InMux I__3802 (
            .O(N__24038),
            .I(N__24035));
    LocalMux I__3801 (
            .O(N__24035),
            .I(N__24032));
    Span4Mux_v I__3800 (
            .O(N__24032),
            .I(N__24029));
    Odrv4 I__3799 (
            .O(N__24029),
            .I(n61));
    CascadeMux I__3798 (
            .O(N__24026),
            .I(N__24022));
    InMux I__3797 (
            .O(N__24025),
            .I(N__24017));
    InMux I__3796 (
            .O(N__24022),
            .I(N__24017));
    LocalMux I__3795 (
            .O(N__24017),
            .I(buf_control_4));
    CascadeMux I__3794 (
            .O(N__24014),
            .I(N__24011));
    InMux I__3793 (
            .O(N__24011),
            .I(N__24002));
    InMux I__3792 (
            .O(N__24010),
            .I(N__24002));
    InMux I__3791 (
            .O(N__24009),
            .I(N__24002));
    LocalMux I__3790 (
            .O(N__24002),
            .I(cmd_rdadctmp_25_adj_1087));
    CascadeMux I__3789 (
            .O(N__23999),
            .I(N__23996));
    InMux I__3788 (
            .O(N__23996),
            .I(N__23993));
    LocalMux I__3787 (
            .O(N__23993),
            .I(N__23989));
    InMux I__3786 (
            .O(N__23992),
            .I(N__23986));
    Odrv12 I__3785 (
            .O(N__23989),
            .I(cmd_rdadctmp_7_adj_1105));
    LocalMux I__3784 (
            .O(N__23986),
            .I(cmd_rdadctmp_7_adj_1105));
    CascadeMux I__3783 (
            .O(N__23981),
            .I(n16500_cascade_));
    InMux I__3782 (
            .O(N__23978),
            .I(N__23975));
    LocalMux I__3781 (
            .O(N__23975),
            .I(N__23972));
    Span4Mux_h I__3780 (
            .O(N__23972),
            .I(N__23969));
    Sp12to4 I__3779 (
            .O(N__23969),
            .I(N__23966));
    Span12Mux_v I__3778 (
            .O(N__23966),
            .I(N__23963));
    Odrv12 I__3777 (
            .O(N__23963),
            .I(buf_data4_12));
    CascadeMux I__3776 (
            .O(N__23960),
            .I(N__23957));
    InMux I__3775 (
            .O(N__23957),
            .I(N__23954));
    LocalMux I__3774 (
            .O(N__23954),
            .I(comm_buf_10_4));
    InMux I__3773 (
            .O(N__23951),
            .I(N__23948));
    LocalMux I__3772 (
            .O(N__23948),
            .I(N__23945));
    Span4Mux_h I__3771 (
            .O(N__23945),
            .I(N__23942));
    Span4Mux_h I__3770 (
            .O(N__23942),
            .I(N__23939));
    Span4Mux_h I__3769 (
            .O(N__23939),
            .I(N__23936));
    Span4Mux_h I__3768 (
            .O(N__23936),
            .I(N__23933));
    Odrv4 I__3767 (
            .O(N__23933),
            .I(buf_data4_15));
    InMux I__3766 (
            .O(N__23930),
            .I(N__23927));
    LocalMux I__3765 (
            .O(N__23927),
            .I(N__23924));
    Span4Mux_v I__3764 (
            .O(N__23924),
            .I(N__23921));
    Sp12to4 I__3763 (
            .O(N__23921),
            .I(N__23918));
    Odrv12 I__3762 (
            .O(N__23918),
            .I(comm_buf_10_7));
    InMux I__3761 (
            .O(N__23915),
            .I(N__23912));
    LocalMux I__3760 (
            .O(N__23912),
            .I(N__23909));
    Span4Mux_v I__3759 (
            .O(N__23909),
            .I(N__23906));
    Sp12to4 I__3758 (
            .O(N__23906),
            .I(N__23903));
    Span12Mux_h I__3757 (
            .O(N__23903),
            .I(N__23900));
    Span12Mux_v I__3756 (
            .O(N__23900),
            .I(N__23897));
    Odrv12 I__3755 (
            .O(N__23897),
            .I(buf_data4_8));
    InMux I__3754 (
            .O(N__23894),
            .I(N__23891));
    LocalMux I__3753 (
            .O(N__23891),
            .I(N__23888));
    Span4Mux_v I__3752 (
            .O(N__23888),
            .I(N__23885));
    Odrv4 I__3751 (
            .O(N__23885),
            .I(comm_buf_10_0));
    CascadeMux I__3750 (
            .O(N__23882),
            .I(n16434_cascade_));
    CascadeMux I__3749 (
            .O(N__23879),
            .I(n16437_cascade_));
    InMux I__3748 (
            .O(N__23876),
            .I(N__23873));
    LocalMux I__3747 (
            .O(N__23873),
            .I(n109));
    CascadeMux I__3746 (
            .O(N__23870),
            .I(n8054_cascade_));
    InMux I__3745 (
            .O(N__23867),
            .I(N__23864));
    LocalMux I__3744 (
            .O(N__23864),
            .I(N__23861));
    Odrv12 I__3743 (
            .O(N__23861),
            .I(n59));
    CascadeMux I__3742 (
            .O(N__23858),
            .I(n8907_cascade_));
    CEMux I__3741 (
            .O(N__23855),
            .I(N__23852));
    LocalMux I__3740 (
            .O(N__23852),
            .I(n8943));
    CascadeMux I__3739 (
            .O(N__23849),
            .I(n8943_cascade_));
    SRMux I__3738 (
            .O(N__23846),
            .I(N__23843));
    LocalMux I__3737 (
            .O(N__23843),
            .I(N__23840));
    Odrv12 I__3736 (
            .O(N__23840),
            .I(n10625));
    CEMux I__3735 (
            .O(N__23837),
            .I(N__23834));
    LocalMux I__3734 (
            .O(N__23834),
            .I(N__23831));
    Span4Mux_h I__3733 (
            .O(N__23831),
            .I(N__23828));
    Odrv4 I__3732 (
            .O(N__23828),
            .I(n9123));
    CascadeMux I__3731 (
            .O(N__23825),
            .I(n9123_cascade_));
    SRMux I__3730 (
            .O(N__23822),
            .I(N__23819));
    LocalMux I__3729 (
            .O(N__23819),
            .I(n10653));
    InMux I__3728 (
            .O(N__23816),
            .I(N__23813));
    LocalMux I__3727 (
            .O(N__23813),
            .I(N__23810));
    Sp12to4 I__3726 (
            .O(N__23810),
            .I(N__23807));
    Span12Mux_v I__3725 (
            .O(N__23807),
            .I(N__23804));
    Odrv12 I__3724 (
            .O(N__23804),
            .I(buf_data3_16));
    InMux I__3723 (
            .O(N__23801),
            .I(N__23798));
    LocalMux I__3722 (
            .O(N__23798),
            .I(N__23795));
    Span4Mux_v I__3721 (
            .O(N__23795),
            .I(N__23792));
    Odrv4 I__3720 (
            .O(N__23792),
            .I(comm_buf_6_0));
    InMux I__3719 (
            .O(N__23789),
            .I(N__23786));
    LocalMux I__3718 (
            .O(N__23786),
            .I(N__23783));
    Sp12to4 I__3717 (
            .O(N__23783),
            .I(N__23780));
    Span12Mux_v I__3716 (
            .O(N__23780),
            .I(N__23777));
    Odrv12 I__3715 (
            .O(N__23777),
            .I(buf_data3_17));
    InMux I__3714 (
            .O(N__23774),
            .I(N__23771));
    LocalMux I__3713 (
            .O(N__23771),
            .I(N__23768));
    Span4Mux_h I__3712 (
            .O(N__23768),
            .I(N__23765));
    Odrv4 I__3711 (
            .O(N__23765),
            .I(comm_buf_6_1));
    CEMux I__3710 (
            .O(N__23762),
            .I(N__23758));
    CEMux I__3709 (
            .O(N__23761),
            .I(N__23755));
    LocalMux I__3708 (
            .O(N__23758),
            .I(N__23752));
    LocalMux I__3707 (
            .O(N__23755),
            .I(N__23749));
    Odrv12 I__3706 (
            .O(N__23752),
            .I(n8907));
    Odrv4 I__3705 (
            .O(N__23749),
            .I(n8907));
    SRMux I__3704 (
            .O(N__23744),
            .I(N__23740));
    SRMux I__3703 (
            .O(N__23743),
            .I(N__23737));
    LocalMux I__3702 (
            .O(N__23740),
            .I(N__23734));
    LocalMux I__3701 (
            .O(N__23737),
            .I(N__23731));
    Span4Mux_h I__3700 (
            .O(N__23734),
            .I(N__23728));
    Odrv12 I__3699 (
            .O(N__23731),
            .I(n10618));
    Odrv4 I__3698 (
            .O(N__23728),
            .I(n10618));
    InMux I__3697 (
            .O(N__23723),
            .I(N__23720));
    LocalMux I__3696 (
            .O(N__23720),
            .I(N__23717));
    Span4Mux_h I__3695 (
            .O(N__23717),
            .I(N__23714));
    Sp12to4 I__3694 (
            .O(N__23714),
            .I(N__23711));
    Span12Mux_v I__3693 (
            .O(N__23711),
            .I(N__23708));
    Odrv12 I__3692 (
            .O(N__23708),
            .I(buf_data4_10));
    InMux I__3691 (
            .O(N__23705),
            .I(N__23702));
    LocalMux I__3690 (
            .O(N__23702),
            .I(N__23699));
    Span4Mux_h I__3689 (
            .O(N__23699),
            .I(N__23696));
    Odrv4 I__3688 (
            .O(N__23696),
            .I(comm_buf_10_2));
    InMux I__3687 (
            .O(N__23693),
            .I(N__23690));
    LocalMux I__3686 (
            .O(N__23690),
            .I(N__23687));
    Span4Mux_h I__3685 (
            .O(N__23687),
            .I(N__23684));
    Span4Mux_v I__3684 (
            .O(N__23684),
            .I(N__23681));
    Span4Mux_h I__3683 (
            .O(N__23681),
            .I(N__23678));
    Span4Mux_h I__3682 (
            .O(N__23678),
            .I(N__23675));
    Odrv4 I__3681 (
            .O(N__23675),
            .I(buf_data4_11));
    InMux I__3680 (
            .O(N__23672),
            .I(N__23669));
    LocalMux I__3679 (
            .O(N__23669),
            .I(N__23666));
    Span4Mux_h I__3678 (
            .O(N__23666),
            .I(N__23663));
    Odrv4 I__3677 (
            .O(N__23663),
            .I(comm_buf_10_3));
    InMux I__3676 (
            .O(N__23660),
            .I(N__23657));
    LocalMux I__3675 (
            .O(N__23657),
            .I(N__23654));
    Span4Mux_v I__3674 (
            .O(N__23654),
            .I(N__23651));
    Sp12to4 I__3673 (
            .O(N__23651),
            .I(N__23648));
    Odrv12 I__3672 (
            .O(N__23648),
            .I(buf_data3_1));
    InMux I__3671 (
            .O(N__23645),
            .I(N__23642));
    LocalMux I__3670 (
            .O(N__23642),
            .I(N__23639));
    Span4Mux_v I__3669 (
            .O(N__23639),
            .I(N__23636));
    Odrv4 I__3668 (
            .O(N__23636),
            .I(comm_buf_8_1));
    InMux I__3667 (
            .O(N__23633),
            .I(N__23630));
    LocalMux I__3666 (
            .O(N__23630),
            .I(N__23627));
    Span4Mux_v I__3665 (
            .O(N__23627),
            .I(N__23624));
    Span4Mux_h I__3664 (
            .O(N__23624),
            .I(N__23621));
    Span4Mux_h I__3663 (
            .O(N__23621),
            .I(N__23618));
    Odrv4 I__3662 (
            .O(N__23618),
            .I(buf_data3_0));
    InMux I__3661 (
            .O(N__23615),
            .I(N__23612));
    LocalMux I__3660 (
            .O(N__23612),
            .I(N__23609));
    Span4Mux_h I__3659 (
            .O(N__23609),
            .I(N__23606));
    Odrv4 I__3658 (
            .O(N__23606),
            .I(comm_buf_8_0));
    InMux I__3657 (
            .O(N__23603),
            .I(N__23600));
    LocalMux I__3656 (
            .O(N__23600),
            .I(N__23597));
    Sp12to4 I__3655 (
            .O(N__23597),
            .I(N__23594));
    Span12Mux_v I__3654 (
            .O(N__23594),
            .I(N__23591));
    Odrv12 I__3653 (
            .O(N__23591),
            .I(buf_data3_23));
    InMux I__3652 (
            .O(N__23588),
            .I(N__23585));
    LocalMux I__3651 (
            .O(N__23585),
            .I(comm_buf_6_7));
    InMux I__3650 (
            .O(N__23582),
            .I(N__23579));
    LocalMux I__3649 (
            .O(N__23579),
            .I(N__23576));
    Sp12to4 I__3648 (
            .O(N__23576),
            .I(N__23573));
    Span12Mux_v I__3647 (
            .O(N__23573),
            .I(N__23570));
    Odrv12 I__3646 (
            .O(N__23570),
            .I(buf_data3_22));
    InMux I__3645 (
            .O(N__23567),
            .I(N__23564));
    LocalMux I__3644 (
            .O(N__23564),
            .I(N__23561));
    Span4Mux_v I__3643 (
            .O(N__23561),
            .I(N__23558));
    Span4Mux_h I__3642 (
            .O(N__23558),
            .I(N__23555));
    Odrv4 I__3641 (
            .O(N__23555),
            .I(comm_buf_6_6));
    InMux I__3640 (
            .O(N__23552),
            .I(N__23549));
    LocalMux I__3639 (
            .O(N__23549),
            .I(N__23546));
    Span4Mux_v I__3638 (
            .O(N__23546),
            .I(N__23543));
    Sp12to4 I__3637 (
            .O(N__23543),
            .I(N__23540));
    Odrv12 I__3636 (
            .O(N__23540),
            .I(buf_data3_21));
    InMux I__3635 (
            .O(N__23537),
            .I(N__23534));
    LocalMux I__3634 (
            .O(N__23534),
            .I(N__23531));
    Span12Mux_h I__3633 (
            .O(N__23531),
            .I(N__23528));
    Odrv12 I__3632 (
            .O(N__23528),
            .I(comm_buf_6_5));
    InMux I__3631 (
            .O(N__23525),
            .I(N__23522));
    LocalMux I__3630 (
            .O(N__23522),
            .I(N__23519));
    Sp12to4 I__3629 (
            .O(N__23519),
            .I(N__23516));
    Span12Mux_v I__3628 (
            .O(N__23516),
            .I(N__23513));
    Odrv12 I__3627 (
            .O(N__23513),
            .I(buf_data3_20));
    InMux I__3626 (
            .O(N__23510),
            .I(N__23507));
    LocalMux I__3625 (
            .O(N__23507),
            .I(N__23504));
    Odrv4 I__3624 (
            .O(N__23504),
            .I(comm_buf_6_4));
    InMux I__3623 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__3622 (
            .O(N__23498),
            .I(N__23495));
    Span4Mux_v I__3621 (
            .O(N__23495),
            .I(N__23492));
    Sp12to4 I__3620 (
            .O(N__23492),
            .I(N__23489));
    Odrv12 I__3619 (
            .O(N__23489),
            .I(buf_data3_19));
    InMux I__3618 (
            .O(N__23486),
            .I(N__23483));
    LocalMux I__3617 (
            .O(N__23483),
            .I(N__23480));
    Span4Mux_h I__3616 (
            .O(N__23480),
            .I(N__23477));
    Odrv4 I__3615 (
            .O(N__23477),
            .I(comm_buf_6_3));
    InMux I__3614 (
            .O(N__23474),
            .I(N__23471));
    LocalMux I__3613 (
            .O(N__23471),
            .I(N__23468));
    Span4Mux_v I__3612 (
            .O(N__23468),
            .I(N__23465));
    Span4Mux_h I__3611 (
            .O(N__23465),
            .I(N__23462));
    Span4Mux_h I__3610 (
            .O(N__23462),
            .I(N__23459));
    Span4Mux_h I__3609 (
            .O(N__23459),
            .I(N__23456));
    Odrv4 I__3608 (
            .O(N__23456),
            .I(buf_data3_18));
    InMux I__3607 (
            .O(N__23453),
            .I(N__23450));
    LocalMux I__3606 (
            .O(N__23450),
            .I(N__23447));
    Span4Mux_v I__3605 (
            .O(N__23447),
            .I(N__23444));
    Span4Mux_h I__3604 (
            .O(N__23444),
            .I(N__23441));
    Odrv4 I__3603 (
            .O(N__23441),
            .I(comm_buf_6_2));
    CascadeMux I__3602 (
            .O(N__23438),
            .I(N__23435));
    InMux I__3601 (
            .O(N__23435),
            .I(N__23431));
    CascadeMux I__3600 (
            .O(N__23434),
            .I(N__23427));
    LocalMux I__3599 (
            .O(N__23431),
            .I(N__23424));
    InMux I__3598 (
            .O(N__23430),
            .I(N__23419));
    InMux I__3597 (
            .O(N__23427),
            .I(N__23419));
    Odrv4 I__3596 (
            .O(N__23424),
            .I(cmd_rdadctmp_30_adj_1119));
    LocalMux I__3595 (
            .O(N__23419),
            .I(cmd_rdadctmp_30_adj_1119));
    InMux I__3594 (
            .O(N__23414),
            .I(N__23408));
    InMux I__3593 (
            .O(N__23413),
            .I(N__23408));
    LocalMux I__3592 (
            .O(N__23408),
            .I(cmd_rdadctmp_31_adj_1118));
    InMux I__3591 (
            .O(N__23405),
            .I(N__23402));
    LocalMux I__3590 (
            .O(N__23402),
            .I(N__23399));
    Span4Mux_v I__3589 (
            .O(N__23399),
            .I(N__23396));
    Sp12to4 I__3588 (
            .O(N__23396),
            .I(N__23393));
    Odrv12 I__3587 (
            .O(N__23393),
            .I(buf_data3_7));
    InMux I__3586 (
            .O(N__23390),
            .I(N__23387));
    LocalMux I__3585 (
            .O(N__23387),
            .I(N__23384));
    Odrv4 I__3584 (
            .O(N__23384),
            .I(comm_buf_8_7));
    InMux I__3583 (
            .O(N__23381),
            .I(N__23378));
    LocalMux I__3582 (
            .O(N__23378),
            .I(N__23375));
    Span4Mux_h I__3581 (
            .O(N__23375),
            .I(N__23372));
    Odrv4 I__3580 (
            .O(N__23372),
            .I(buf_data3_6));
    InMux I__3579 (
            .O(N__23369),
            .I(N__23366));
    LocalMux I__3578 (
            .O(N__23366),
            .I(N__23363));
    Span4Mux_h I__3577 (
            .O(N__23363),
            .I(N__23360));
    Odrv4 I__3576 (
            .O(N__23360),
            .I(comm_buf_8_6));
    InMux I__3575 (
            .O(N__23357),
            .I(N__23354));
    LocalMux I__3574 (
            .O(N__23354),
            .I(N__23351));
    Span4Mux_h I__3573 (
            .O(N__23351),
            .I(N__23348));
    Span4Mux_h I__3572 (
            .O(N__23348),
            .I(N__23345));
    Odrv4 I__3571 (
            .O(N__23345),
            .I(buf_data3_5));
    InMux I__3570 (
            .O(N__23342),
            .I(N__23339));
    LocalMux I__3569 (
            .O(N__23339),
            .I(N__23336));
    Odrv4 I__3568 (
            .O(N__23336),
            .I(comm_buf_8_5));
    InMux I__3567 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__3566 (
            .O(N__23330),
            .I(N__23327));
    Span4Mux_h I__3565 (
            .O(N__23327),
            .I(N__23324));
    Span4Mux_h I__3564 (
            .O(N__23324),
            .I(N__23321));
    Odrv4 I__3563 (
            .O(N__23321),
            .I(buf_data3_4));
    InMux I__3562 (
            .O(N__23318),
            .I(N__23315));
    LocalMux I__3561 (
            .O(N__23315),
            .I(N__23312));
    Span4Mux_v I__3560 (
            .O(N__23312),
            .I(N__23309));
    Odrv4 I__3559 (
            .O(N__23309),
            .I(comm_buf_8_4));
    InMux I__3558 (
            .O(N__23306),
            .I(N__23303));
    LocalMux I__3557 (
            .O(N__23303),
            .I(N__23300));
    Span4Mux_v I__3556 (
            .O(N__23300),
            .I(N__23297));
    Span4Mux_h I__3555 (
            .O(N__23297),
            .I(N__23294));
    Span4Mux_h I__3554 (
            .O(N__23294),
            .I(N__23291));
    Odrv4 I__3553 (
            .O(N__23291),
            .I(buf_data3_3));
    InMux I__3552 (
            .O(N__23288),
            .I(N__23285));
    LocalMux I__3551 (
            .O(N__23285),
            .I(N__23282));
    Span4Mux_v I__3550 (
            .O(N__23282),
            .I(N__23279));
    Span4Mux_h I__3549 (
            .O(N__23279),
            .I(N__23276));
    Odrv4 I__3548 (
            .O(N__23276),
            .I(comm_buf_8_3));
    InMux I__3547 (
            .O(N__23273),
            .I(N__23270));
    LocalMux I__3546 (
            .O(N__23270),
            .I(N__23267));
    Span12Mux_h I__3545 (
            .O(N__23267),
            .I(N__23264));
    Odrv12 I__3544 (
            .O(N__23264),
            .I(buf_data3_2));
    CascadeMux I__3543 (
            .O(N__23261),
            .I(N__23258));
    InMux I__3542 (
            .O(N__23258),
            .I(N__23255));
    LocalMux I__3541 (
            .O(N__23255),
            .I(N__23252));
    Span4Mux_h I__3540 (
            .O(N__23252),
            .I(N__23249));
    Odrv4 I__3539 (
            .O(N__23249),
            .I(comm_buf_8_2));
    InMux I__3538 (
            .O(N__23246),
            .I(\ADC_VAC4.n14007 ));
    InMux I__3537 (
            .O(N__23243),
            .I(\ADC_VAC4.n14008 ));
    InMux I__3536 (
            .O(N__23240),
            .I(N__23237));
    LocalMux I__3535 (
            .O(N__23237),
            .I(N__23232));
    InMux I__3534 (
            .O(N__23236),
            .I(N__23229));
    InMux I__3533 (
            .O(N__23235),
            .I(N__23226));
    Odrv4 I__3532 (
            .O(N__23232),
            .I(\comm_spi.n16908 ));
    LocalMux I__3531 (
            .O(N__23229),
            .I(\comm_spi.n16908 ));
    LocalMux I__3530 (
            .O(N__23226),
            .I(\comm_spi.n16908 ));
    InMux I__3529 (
            .O(N__23219),
            .I(N__23216));
    LocalMux I__3528 (
            .O(N__23216),
            .I(N__23212));
    InMux I__3527 (
            .O(N__23215),
            .I(N__23209));
    Odrv4 I__3526 (
            .O(N__23212),
            .I(\comm_spi.n10459 ));
    LocalMux I__3525 (
            .O(N__23209),
            .I(\comm_spi.n10459 ));
    InMux I__3524 (
            .O(N__23204),
            .I(N__23201));
    LocalMux I__3523 (
            .O(N__23201),
            .I(N__23197));
    InMux I__3522 (
            .O(N__23200),
            .I(N__23194));
    Span4Mux_h I__3521 (
            .O(N__23197),
            .I(N__23189));
    LocalMux I__3520 (
            .O(N__23194),
            .I(N__23189));
    Odrv4 I__3519 (
            .O(N__23189),
            .I(\comm_spi.n10460 ));
    SRMux I__3518 (
            .O(N__23186),
            .I(N__23183));
    LocalMux I__3517 (
            .O(N__23183),
            .I(N__23180));
    Odrv12 I__3516 (
            .O(N__23180),
            .I(\comm_spi.data_tx_7__N_828 ));
    CascadeMux I__3515 (
            .O(N__23177),
            .I(N__23174));
    InMux I__3514 (
            .O(N__23174),
            .I(N__23170));
    InMux I__3513 (
            .O(N__23173),
            .I(N__23167));
    LocalMux I__3512 (
            .O(N__23170),
            .I(N__23163));
    LocalMux I__3511 (
            .O(N__23167),
            .I(N__23160));
    InMux I__3510 (
            .O(N__23166),
            .I(N__23157));
    Span4Mux_h I__3509 (
            .O(N__23163),
            .I(N__23154));
    Span12Mux_h I__3508 (
            .O(N__23160),
            .I(N__23151));
    LocalMux I__3507 (
            .O(N__23157),
            .I(buf_adcdata4_21));
    Odrv4 I__3506 (
            .O(N__23154),
            .I(buf_adcdata4_21));
    Odrv12 I__3505 (
            .O(N__23151),
            .I(buf_adcdata4_21));
    CascadeMux I__3504 (
            .O(N__23144),
            .I(N__23141));
    InMux I__3503 (
            .O(N__23141),
            .I(N__23132));
    InMux I__3502 (
            .O(N__23140),
            .I(N__23132));
    InMux I__3501 (
            .O(N__23139),
            .I(N__23132));
    LocalMux I__3500 (
            .O(N__23132),
            .I(cmd_rdadctmp_29_adj_1120));
    CascadeMux I__3499 (
            .O(N__23129),
            .I(N__23125));
    InMux I__3498 (
            .O(N__23128),
            .I(N__23118));
    InMux I__3497 (
            .O(N__23125),
            .I(N__23118));
    CascadeMux I__3496 (
            .O(N__23124),
            .I(N__23115));
    InMux I__3495 (
            .O(N__23123),
            .I(N__23112));
    LocalMux I__3494 (
            .O(N__23118),
            .I(N__23108));
    InMux I__3493 (
            .O(N__23115),
            .I(N__23105));
    LocalMux I__3492 (
            .O(N__23112),
            .I(N__23102));
    InMux I__3491 (
            .O(N__23111),
            .I(N__23099));
    Span4Mux_v I__3490 (
            .O(N__23108),
            .I(N__23094));
    LocalMux I__3489 (
            .O(N__23105),
            .I(N__23094));
    Span4Mux_v I__3488 (
            .O(N__23102),
            .I(N__23091));
    LocalMux I__3487 (
            .O(N__23099),
            .I(N__23088));
    Span4Mux_v I__3486 (
            .O(N__23094),
            .I(N__23085));
    Span4Mux_v I__3485 (
            .O(N__23091),
            .I(N__23080));
    Span4Mux_v I__3484 (
            .O(N__23088),
            .I(N__23080));
    Sp12to4 I__3483 (
            .O(N__23085),
            .I(N__23075));
    Sp12to4 I__3482 (
            .O(N__23080),
            .I(N__23075));
    Span12Mux_h I__3481 (
            .O(N__23075),
            .I(N__23072));
    Odrv12 I__3480 (
            .O(N__23072),
            .I(M_DRDY3));
    CascadeMux I__3479 (
            .O(N__23069),
            .I(N__23063));
    InMux I__3478 (
            .O(N__23068),
            .I(N__23059));
    InMux I__3477 (
            .O(N__23067),
            .I(N__23050));
    InMux I__3476 (
            .O(N__23066),
            .I(N__23050));
    InMux I__3475 (
            .O(N__23063),
            .I(N__23050));
    InMux I__3474 (
            .O(N__23062),
            .I(N__23046));
    LocalMux I__3473 (
            .O(N__23059),
            .I(N__23043));
    InMux I__3472 (
            .O(N__23058),
            .I(N__23036));
    InMux I__3471 (
            .O(N__23057),
            .I(N__23033));
    LocalMux I__3470 (
            .O(N__23050),
            .I(N__23030));
    InMux I__3469 (
            .O(N__23049),
            .I(N__23027));
    LocalMux I__3468 (
            .O(N__23046),
            .I(N__23024));
    Span4Mux_h I__3467 (
            .O(N__23043),
            .I(N__23021));
    InMux I__3466 (
            .O(N__23042),
            .I(N__23018));
    InMux I__3465 (
            .O(N__23041),
            .I(N__23011));
    InMux I__3464 (
            .O(N__23040),
            .I(N__23011));
    InMux I__3463 (
            .O(N__23039),
            .I(N__23011));
    LocalMux I__3462 (
            .O(N__23036),
            .I(N__23004));
    LocalMux I__3461 (
            .O(N__23033),
            .I(N__23004));
    Span4Mux_h I__3460 (
            .O(N__23030),
            .I(N__23004));
    LocalMux I__3459 (
            .O(N__23027),
            .I(adc_state_1_adj_1079));
    Odrv4 I__3458 (
            .O(N__23024),
            .I(adc_state_1_adj_1079));
    Odrv4 I__3457 (
            .O(N__23021),
            .I(adc_state_1_adj_1079));
    LocalMux I__3456 (
            .O(N__23018),
            .I(adc_state_1_adj_1079));
    LocalMux I__3455 (
            .O(N__23011),
            .I(adc_state_1_adj_1079));
    Odrv4 I__3454 (
            .O(N__23004),
            .I(adc_state_1_adj_1079));
    CEMux I__3453 (
            .O(N__22991),
            .I(N__22988));
    LocalMux I__3452 (
            .O(N__22988),
            .I(\ADC_VAC3.n9514 ));
    InMux I__3451 (
            .O(N__22985),
            .I(N__22973));
    InMux I__3450 (
            .O(N__22984),
            .I(N__22973));
    InMux I__3449 (
            .O(N__22983),
            .I(N__22966));
    InMux I__3448 (
            .O(N__22982),
            .I(N__22966));
    InMux I__3447 (
            .O(N__22981),
            .I(N__22966));
    CascadeMux I__3446 (
            .O(N__22980),
            .I(N__22963));
    InMux I__3445 (
            .O(N__22979),
            .I(N__22960));
    InMux I__3444 (
            .O(N__22978),
            .I(N__22957));
    LocalMux I__3443 (
            .O(N__22973),
            .I(N__22948));
    LocalMux I__3442 (
            .O(N__22966),
            .I(N__22948));
    InMux I__3441 (
            .O(N__22963),
            .I(N__22945));
    LocalMux I__3440 (
            .O(N__22960),
            .I(N__22940));
    LocalMux I__3439 (
            .O(N__22957),
            .I(N__22940));
    InMux I__3438 (
            .O(N__22956),
            .I(N__22937));
    InMux I__3437 (
            .O(N__22955),
            .I(N__22930));
    InMux I__3436 (
            .O(N__22954),
            .I(N__22930));
    InMux I__3435 (
            .O(N__22953),
            .I(N__22930));
    Span4Mux_v I__3434 (
            .O(N__22948),
            .I(N__22927));
    LocalMux I__3433 (
            .O(N__22945),
            .I(DTRIG_N_957_adj_1114));
    Odrv4 I__3432 (
            .O(N__22940),
            .I(DTRIG_N_957_adj_1114));
    LocalMux I__3431 (
            .O(N__22937),
            .I(DTRIG_N_957_adj_1114));
    LocalMux I__3430 (
            .O(N__22930),
            .I(DTRIG_N_957_adj_1114));
    Odrv4 I__3429 (
            .O(N__22927),
            .I(DTRIG_N_957_adj_1114));
    CascadeMux I__3428 (
            .O(N__22916),
            .I(\ADC_VAC3.n9514_cascade_ ));
    SRMux I__3427 (
            .O(N__22913),
            .I(N__22910));
    LocalMux I__3426 (
            .O(N__22910),
            .I(N__22907));
    Span4Mux_h I__3425 (
            .O(N__22907),
            .I(N__22904));
    Odrv4 I__3424 (
            .O(N__22904),
            .I(\ADC_VAC3.n10744 ));
    InMux I__3423 (
            .O(N__22901),
            .I(bfn_10_17_0_));
    InMux I__3422 (
            .O(N__22898),
            .I(\ADC_VAC4.n14002 ));
    InMux I__3421 (
            .O(N__22895),
            .I(\ADC_VAC4.n14003 ));
    InMux I__3420 (
            .O(N__22892),
            .I(\ADC_VAC4.n14004 ));
    InMux I__3419 (
            .O(N__22889),
            .I(\ADC_VAC4.n14005 ));
    InMux I__3418 (
            .O(N__22886),
            .I(\ADC_VAC4.n14006 ));
    InMux I__3417 (
            .O(N__22883),
            .I(N__22879));
    InMux I__3416 (
            .O(N__22882),
            .I(N__22876));
    LocalMux I__3415 (
            .O(N__22879),
            .I(\ADC_VAC3.bit_cnt_0 ));
    LocalMux I__3414 (
            .O(N__22876),
            .I(\ADC_VAC3.bit_cnt_0 ));
    InMux I__3413 (
            .O(N__22871),
            .I(bfn_10_15_0_));
    CascadeMux I__3412 (
            .O(N__22868),
            .I(N__22864));
    InMux I__3411 (
            .O(N__22867),
            .I(N__22861));
    InMux I__3410 (
            .O(N__22864),
            .I(N__22858));
    LocalMux I__3409 (
            .O(N__22861),
            .I(\ADC_VAC3.bit_cnt_1 ));
    LocalMux I__3408 (
            .O(N__22858),
            .I(\ADC_VAC3.bit_cnt_1 ));
    InMux I__3407 (
            .O(N__22853),
            .I(\ADC_VAC3.n13995 ));
    InMux I__3406 (
            .O(N__22850),
            .I(N__22846));
    InMux I__3405 (
            .O(N__22849),
            .I(N__22843));
    LocalMux I__3404 (
            .O(N__22846),
            .I(\ADC_VAC3.bit_cnt_2 ));
    LocalMux I__3403 (
            .O(N__22843),
            .I(\ADC_VAC3.bit_cnt_2 ));
    InMux I__3402 (
            .O(N__22838),
            .I(\ADC_VAC3.n13996 ));
    InMux I__3401 (
            .O(N__22835),
            .I(N__22831));
    InMux I__3400 (
            .O(N__22834),
            .I(N__22828));
    LocalMux I__3399 (
            .O(N__22831),
            .I(\ADC_VAC3.bit_cnt_3 ));
    LocalMux I__3398 (
            .O(N__22828),
            .I(\ADC_VAC3.bit_cnt_3 ));
    InMux I__3397 (
            .O(N__22823),
            .I(\ADC_VAC3.n13997 ));
    InMux I__3396 (
            .O(N__22820),
            .I(N__22816));
    InMux I__3395 (
            .O(N__22819),
            .I(N__22813));
    LocalMux I__3394 (
            .O(N__22816),
            .I(\ADC_VAC3.bit_cnt_4 ));
    LocalMux I__3393 (
            .O(N__22813),
            .I(\ADC_VAC3.bit_cnt_4 ));
    InMux I__3392 (
            .O(N__22808),
            .I(\ADC_VAC3.n13998 ));
    InMux I__3391 (
            .O(N__22805),
            .I(N__22801));
    InMux I__3390 (
            .O(N__22804),
            .I(N__22798));
    LocalMux I__3389 (
            .O(N__22801),
            .I(\ADC_VAC3.bit_cnt_5 ));
    LocalMux I__3388 (
            .O(N__22798),
            .I(\ADC_VAC3.bit_cnt_5 ));
    InMux I__3387 (
            .O(N__22793),
            .I(\ADC_VAC3.n13999 ));
    InMux I__3386 (
            .O(N__22790),
            .I(N__22786));
    InMux I__3385 (
            .O(N__22789),
            .I(N__22783));
    LocalMux I__3384 (
            .O(N__22786),
            .I(\ADC_VAC3.bit_cnt_6 ));
    LocalMux I__3383 (
            .O(N__22783),
            .I(\ADC_VAC3.bit_cnt_6 ));
    InMux I__3382 (
            .O(N__22778),
            .I(\ADC_VAC3.n14000 ));
    InMux I__3381 (
            .O(N__22775),
            .I(\ADC_VAC3.n14001 ));
    InMux I__3380 (
            .O(N__22772),
            .I(N__22768));
    InMux I__3379 (
            .O(N__22771),
            .I(N__22765));
    LocalMux I__3378 (
            .O(N__22768),
            .I(\ADC_VAC3.bit_cnt_7 ));
    LocalMux I__3377 (
            .O(N__22765),
            .I(\ADC_VAC3.bit_cnt_7 ));
    CascadeMux I__3376 (
            .O(N__22760),
            .I(N__22757));
    InMux I__3375 (
            .O(N__22757),
            .I(N__22754));
    LocalMux I__3374 (
            .O(N__22754),
            .I(N__22750));
    CascadeMux I__3373 (
            .O(N__22753),
            .I(N__22747));
    Span4Mux_v I__3372 (
            .O(N__22750),
            .I(N__22744));
    InMux I__3371 (
            .O(N__22747),
            .I(N__22741));
    Odrv4 I__3370 (
            .O(N__22744),
            .I(cmd_rdadctmp_31));
    LocalMux I__3369 (
            .O(N__22741),
            .I(cmd_rdadctmp_31));
    InMux I__3368 (
            .O(N__22736),
            .I(N__22733));
    LocalMux I__3367 (
            .O(N__22733),
            .I(N__22730));
    Span12Mux_h I__3366 (
            .O(N__22730),
            .I(N__22726));
    InMux I__3365 (
            .O(N__22729),
            .I(N__22723));
    Span12Mux_v I__3364 (
            .O(N__22726),
            .I(N__22720));
    LocalMux I__3363 (
            .O(N__22723),
            .I(buf_adcdata1_23));
    Odrv12 I__3362 (
            .O(N__22720),
            .I(buf_adcdata1_23));
    InMux I__3361 (
            .O(N__22715),
            .I(N__22712));
    LocalMux I__3360 (
            .O(N__22712),
            .I(N__22707));
    CascadeMux I__3359 (
            .O(N__22711),
            .I(N__22704));
    CascadeMux I__3358 (
            .O(N__22710),
            .I(N__22701));
    Span4Mux_h I__3357 (
            .O(N__22707),
            .I(N__22698));
    InMux I__3356 (
            .O(N__22704),
            .I(N__22693));
    InMux I__3355 (
            .O(N__22701),
            .I(N__22693));
    Odrv4 I__3354 (
            .O(N__22698),
            .I(cmd_rdadctmp_23));
    LocalMux I__3353 (
            .O(N__22693),
            .I(cmd_rdadctmp_23));
    InMux I__3352 (
            .O(N__22688),
            .I(N__22685));
    LocalMux I__3351 (
            .O(N__22685),
            .I(N__22681));
    InMux I__3350 (
            .O(N__22684),
            .I(N__22678));
    Span12Mux_s7_h I__3349 (
            .O(N__22681),
            .I(N__22675));
    LocalMux I__3348 (
            .O(N__22678),
            .I(buf_adcdata1_15));
    Odrv12 I__3347 (
            .O(N__22675),
            .I(buf_adcdata1_15));
    CascadeMux I__3346 (
            .O(N__22670),
            .I(N__22667));
    InMux I__3345 (
            .O(N__22667),
            .I(N__22663));
    CascadeMux I__3344 (
            .O(N__22666),
            .I(N__22660));
    LocalMux I__3343 (
            .O(N__22663),
            .I(N__22657));
    InMux I__3342 (
            .O(N__22660),
            .I(N__22653));
    Span4Mux_h I__3341 (
            .O(N__22657),
            .I(N__22650));
    InMux I__3340 (
            .O(N__22656),
            .I(N__22647));
    LocalMux I__3339 (
            .O(N__22653),
            .I(cmd_rdadctmp_20_adj_1129));
    Odrv4 I__3338 (
            .O(N__22650),
            .I(cmd_rdadctmp_20_adj_1129));
    LocalMux I__3337 (
            .O(N__22647),
            .I(cmd_rdadctmp_20_adj_1129));
    InMux I__3336 (
            .O(N__22640),
            .I(N__22636));
    InMux I__3335 (
            .O(N__22639),
            .I(N__22633));
    LocalMux I__3334 (
            .O(N__22636),
            .I(\ADC_VAC2.bit_cnt_4 ));
    LocalMux I__3333 (
            .O(N__22633),
            .I(\ADC_VAC2.bit_cnt_4 ));
    InMux I__3332 (
            .O(N__22628),
            .I(N__22624));
    InMux I__3331 (
            .O(N__22627),
            .I(N__22621));
    LocalMux I__3330 (
            .O(N__22624),
            .I(\ADC_VAC2.bit_cnt_3 ));
    LocalMux I__3329 (
            .O(N__22621),
            .I(\ADC_VAC2.bit_cnt_3 ));
    CascadeMux I__3328 (
            .O(N__22616),
            .I(N__22612));
    InMux I__3327 (
            .O(N__22615),
            .I(N__22609));
    InMux I__3326 (
            .O(N__22612),
            .I(N__22606));
    LocalMux I__3325 (
            .O(N__22609),
            .I(\ADC_VAC2.bit_cnt_5 ));
    LocalMux I__3324 (
            .O(N__22606),
            .I(\ADC_VAC2.bit_cnt_5 ));
    InMux I__3323 (
            .O(N__22601),
            .I(N__22597));
    InMux I__3322 (
            .O(N__22600),
            .I(N__22594));
    LocalMux I__3321 (
            .O(N__22597),
            .I(\ADC_VAC2.bit_cnt_2 ));
    LocalMux I__3320 (
            .O(N__22594),
            .I(\ADC_VAC2.bit_cnt_2 ));
    InMux I__3319 (
            .O(N__22589),
            .I(N__22586));
    LocalMux I__3318 (
            .O(N__22586),
            .I(\ADC_VAC2.n15596 ));
    CascadeMux I__3317 (
            .O(N__22583),
            .I(\ADC_VAC3.n15334_cascade_ ));
    CascadeMux I__3316 (
            .O(N__22580),
            .I(\ADC_VAC3.n15358_cascade_ ));
    CascadeMux I__3315 (
            .O(N__22577),
            .I(\ADC_VAC3.n15602_cascade_ ));
    CEMux I__3314 (
            .O(N__22574),
            .I(N__22571));
    LocalMux I__3313 (
            .O(N__22571),
            .I(N__22568));
    Span4Mux_v I__3312 (
            .O(N__22568),
            .I(N__22565));
    Span4Mux_h I__3311 (
            .O(N__22565),
            .I(N__22562));
    Odrv4 I__3310 (
            .O(N__22562),
            .I(\ADC_VAC3.n15260 ));
    InMux I__3309 (
            .O(N__22559),
            .I(N__22556));
    LocalMux I__3308 (
            .O(N__22556),
            .I(\ADC_VAC3.n15259 ));
    InMux I__3307 (
            .O(N__22553),
            .I(N__22550));
    LocalMux I__3306 (
            .O(N__22550),
            .I(N__22547));
    Span4Mux_h I__3305 (
            .O(N__22547),
            .I(N__22544));
    Odrv4 I__3304 (
            .O(N__22544),
            .I(\ADC_VAC3.n17 ));
    InMux I__3303 (
            .O(N__22541),
            .I(N__22538));
    LocalMux I__3302 (
            .O(N__22538),
            .I(N__22535));
    Odrv4 I__3301 (
            .O(N__22535),
            .I(n8089));
    CascadeMux I__3300 (
            .O(N__22532),
            .I(N__22529));
    InMux I__3299 (
            .O(N__22529),
            .I(N__22526));
    LocalMux I__3298 (
            .O(N__22526),
            .I(N__22523));
    Odrv4 I__3297 (
            .O(N__22523),
            .I(n96_adj_1159));
    CascadeMux I__3296 (
            .O(N__22520),
            .I(n130_adj_1156_cascade_));
    InMux I__3295 (
            .O(N__22517),
            .I(N__22514));
    LocalMux I__3294 (
            .O(N__22514),
            .I(n15587));
    CascadeMux I__3293 (
            .O(N__22511),
            .I(n8051_cascade_));
    CascadeMux I__3292 (
            .O(N__22508),
            .I(N__22505));
    InMux I__3291 (
            .O(N__22505),
            .I(N__22502));
    LocalMux I__3290 (
            .O(N__22502),
            .I(N__22497));
    CascadeMux I__3289 (
            .O(N__22501),
            .I(N__22494));
    CascadeMux I__3288 (
            .O(N__22500),
            .I(N__22491));
    Span4Mux_h I__3287 (
            .O(N__22497),
            .I(N__22488));
    InMux I__3286 (
            .O(N__22494),
            .I(N__22483));
    InMux I__3285 (
            .O(N__22491),
            .I(N__22483));
    Odrv4 I__3284 (
            .O(N__22488),
            .I(cmd_rdadctmp_19_adj_1130));
    LocalMux I__3283 (
            .O(N__22483),
            .I(cmd_rdadctmp_19_adj_1130));
    CascadeMux I__3282 (
            .O(N__22478),
            .I(N__22473));
    CascadeMux I__3281 (
            .O(N__22477),
            .I(N__22470));
    InMux I__3280 (
            .O(N__22476),
            .I(N__22467));
    InMux I__3279 (
            .O(N__22473),
            .I(N__22464));
    InMux I__3278 (
            .O(N__22470),
            .I(N__22461));
    LocalMux I__3277 (
            .O(N__22467),
            .I(N__22456));
    LocalMux I__3276 (
            .O(N__22464),
            .I(N__22456));
    LocalMux I__3275 (
            .O(N__22461),
            .I(cmd_rdadctmp_8));
    Odrv12 I__3274 (
            .O(N__22456),
            .I(cmd_rdadctmp_8));
    InMux I__3273 (
            .O(N__22451),
            .I(N__22448));
    LocalMux I__3272 (
            .O(N__22448),
            .I(N__22445));
    Sp12to4 I__3271 (
            .O(N__22445),
            .I(N__22441));
    InMux I__3270 (
            .O(N__22444),
            .I(N__22438));
    Span12Mux_v I__3269 (
            .O(N__22441),
            .I(N__22435));
    LocalMux I__3268 (
            .O(N__22438),
            .I(buf_adcdata1_0));
    Odrv12 I__3267 (
            .O(N__22435),
            .I(buf_adcdata1_0));
    CascadeMux I__3266 (
            .O(N__22430),
            .I(n76_cascade_));
    CascadeMux I__3265 (
            .O(N__22427),
            .I(n4_adj_1195_cascade_));
    InMux I__3264 (
            .O(N__22424),
            .I(N__22421));
    LocalMux I__3263 (
            .O(N__22421),
            .I(n15632));
    InMux I__3262 (
            .O(N__22418),
            .I(N__22415));
    LocalMux I__3261 (
            .O(N__22415),
            .I(n15589));
    CascadeMux I__3260 (
            .O(N__22412),
            .I(n87_adj_1165_cascade_));
    CascadeMux I__3259 (
            .O(N__22409),
            .I(n69_adj_1161_cascade_));
    InMux I__3258 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__3257 (
            .O(N__22403),
            .I(n130));
    InMux I__3256 (
            .O(N__22400),
            .I(N__22397));
    LocalMux I__3255 (
            .O(N__22397),
            .I(n8050));
    SRMux I__3254 (
            .O(N__22394),
            .I(N__22389));
    SRMux I__3253 (
            .O(N__22393),
            .I(N__22386));
    SRMux I__3252 (
            .O(N__22392),
            .I(N__22380));
    LocalMux I__3251 (
            .O(N__22389),
            .I(N__22377));
    LocalMux I__3250 (
            .O(N__22386),
            .I(N__22374));
    SRMux I__3249 (
            .O(N__22385),
            .I(N__22371));
    SRMux I__3248 (
            .O(N__22384),
            .I(N__22367));
    SRMux I__3247 (
            .O(N__22383),
            .I(N__22364));
    LocalMux I__3246 (
            .O(N__22380),
            .I(N__22361));
    Span4Mux_h I__3245 (
            .O(N__22377),
            .I(N__22358));
    Span4Mux_h I__3244 (
            .O(N__22374),
            .I(N__22355));
    LocalMux I__3243 (
            .O(N__22371),
            .I(N__22352));
    SRMux I__3242 (
            .O(N__22370),
            .I(N__22349));
    LocalMux I__3241 (
            .O(N__22367),
            .I(N__22343));
    LocalMux I__3240 (
            .O(N__22364),
            .I(N__22343));
    Span4Mux_h I__3239 (
            .O(N__22361),
            .I(N__22340));
    Span4Mux_v I__3238 (
            .O(N__22358),
            .I(N__22331));
    Span4Mux_v I__3237 (
            .O(N__22355),
            .I(N__22331));
    Span4Mux_h I__3236 (
            .O(N__22352),
            .I(N__22331));
    LocalMux I__3235 (
            .O(N__22349),
            .I(N__22331));
    SRMux I__3234 (
            .O(N__22348),
            .I(N__22328));
    Span4Mux_h I__3233 (
            .O(N__22343),
            .I(N__22325));
    Span4Mux_h I__3232 (
            .O(N__22340),
            .I(N__22322));
    Span4Mux_v I__3231 (
            .O(N__22331),
            .I(N__22319));
    LocalMux I__3230 (
            .O(N__22328),
            .I(N__22316));
    Odrv4 I__3229 (
            .O(N__22325),
            .I(n10660));
    Odrv4 I__3228 (
            .O(N__22322),
            .I(n10660));
    Odrv4 I__3227 (
            .O(N__22319),
            .I(n10660));
    Odrv12 I__3226 (
            .O(N__22316),
            .I(n10660));
    InMux I__3225 (
            .O(N__22307),
            .I(N__22304));
    LocalMux I__3224 (
            .O(N__22304),
            .I(comm_buf_7_4));
    InMux I__3223 (
            .O(N__22301),
            .I(N__22298));
    LocalMux I__3222 (
            .O(N__22298),
            .I(N__22295));
    Odrv4 I__3221 (
            .O(N__22295),
            .I(comm_buf_11_4));
    InMux I__3220 (
            .O(N__22292),
            .I(N__22289));
    LocalMux I__3219 (
            .O(N__22289),
            .I(comm_buf_9_4));
    CascadeMux I__3218 (
            .O(N__22286),
            .I(n16452_cascade_));
    InMux I__3217 (
            .O(N__22283),
            .I(N__22280));
    LocalMux I__3216 (
            .O(N__22280),
            .I(n16455));
    InMux I__3215 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__3214 (
            .O(N__22274),
            .I(N__22271));
    Span4Mux_v I__3213 (
            .O(N__22271),
            .I(N__22268));
    Span4Mux_h I__3212 (
            .O(N__22268),
            .I(N__22265));
    Odrv4 I__3211 (
            .O(N__22265),
            .I(comm_buf_5_4));
    InMux I__3210 (
            .O(N__22262),
            .I(N__22259));
    LocalMux I__3209 (
            .O(N__22259),
            .I(N__22256));
    Odrv4 I__3208 (
            .O(N__22256),
            .I(comm_buf_4_4));
    InMux I__3207 (
            .O(N__22253),
            .I(N__22250));
    LocalMux I__3206 (
            .O(N__22250),
            .I(n15400));
    CascadeMux I__3205 (
            .O(N__22247),
            .I(n15399_cascade_));
    InMux I__3204 (
            .O(N__22244),
            .I(N__22241));
    LocalMux I__3203 (
            .O(N__22241),
            .I(n16476));
    CascadeMux I__3202 (
            .O(N__22238),
            .I(n15633_cascade_));
    CascadeMux I__3201 (
            .O(N__22235),
            .I(n16458_cascade_));
    CascadeMux I__3200 (
            .O(N__22232),
            .I(n16461_cascade_));
    InMux I__3199 (
            .O(N__22229),
            .I(N__22226));
    LocalMux I__3198 (
            .O(N__22226),
            .I(N__22223));
    Span12Mux_h I__3197 (
            .O(N__22223),
            .I(N__22220));
    Odrv12 I__3196 (
            .O(N__22220),
            .I(comm_buf_7_6));
    InMux I__3195 (
            .O(N__22217),
            .I(N__22214));
    LocalMux I__3194 (
            .O(N__22214),
            .I(N__22211));
    Span12Mux_h I__3193 (
            .O(N__22211),
            .I(N__22208));
    Odrv12 I__3192 (
            .O(N__22208),
            .I(buf_data3_13));
    CascadeMux I__3191 (
            .O(N__22205),
            .I(N__22202));
    InMux I__3190 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__3189 (
            .O(N__22199),
            .I(N__22196));
    Span4Mux_h I__3188 (
            .O(N__22196),
            .I(N__22193));
    Odrv4 I__3187 (
            .O(N__22193),
            .I(comm_buf_7_5));
    InMux I__3186 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__3185 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_h I__3184 (
            .O(N__22184),
            .I(N__22181));
    Span4Mux_v I__3183 (
            .O(N__22181),
            .I(N__22178));
    Span4Mux_h I__3182 (
            .O(N__22178),
            .I(N__22175));
    Span4Mux_h I__3181 (
            .O(N__22175),
            .I(N__22172));
    Odrv4 I__3180 (
            .O(N__22172),
            .I(buf_data3_12));
    InMux I__3179 (
            .O(N__22169),
            .I(N__22166));
    LocalMux I__3178 (
            .O(N__22166),
            .I(N__22163));
    Span4Mux_h I__3177 (
            .O(N__22163),
            .I(N__22160));
    Sp12to4 I__3176 (
            .O(N__22160),
            .I(N__22157));
    Span12Mux_v I__3175 (
            .O(N__22157),
            .I(N__22154));
    Odrv12 I__3174 (
            .O(N__22154),
            .I(buf_data3_11));
    InMux I__3173 (
            .O(N__22151),
            .I(N__22148));
    LocalMux I__3172 (
            .O(N__22148),
            .I(N__22145));
    Odrv4 I__3171 (
            .O(N__22145),
            .I(comm_buf_7_3));
    InMux I__3170 (
            .O(N__22142),
            .I(N__22139));
    LocalMux I__3169 (
            .O(N__22139),
            .I(N__22136));
    Span4Mux_v I__3168 (
            .O(N__22136),
            .I(N__22133));
    Sp12to4 I__3167 (
            .O(N__22133),
            .I(N__22130));
    Span12Mux_h I__3166 (
            .O(N__22130),
            .I(N__22127));
    Span12Mux_v I__3165 (
            .O(N__22127),
            .I(N__22124));
    Odrv12 I__3164 (
            .O(N__22124),
            .I(buf_data3_10));
    InMux I__3163 (
            .O(N__22121),
            .I(N__22118));
    LocalMux I__3162 (
            .O(N__22118),
            .I(N__22115));
    Odrv12 I__3161 (
            .O(N__22115),
            .I(comm_buf_7_2));
    InMux I__3160 (
            .O(N__22112),
            .I(N__22109));
    LocalMux I__3159 (
            .O(N__22109),
            .I(N__22106));
    Span4Mux_h I__3158 (
            .O(N__22106),
            .I(N__22103));
    Sp12to4 I__3157 (
            .O(N__22103),
            .I(N__22100));
    Span12Mux_v I__3156 (
            .O(N__22100),
            .I(N__22097));
    Span12Mux_h I__3155 (
            .O(N__22097),
            .I(N__22094));
    Odrv12 I__3154 (
            .O(N__22094),
            .I(buf_data3_9));
    CascadeMux I__3153 (
            .O(N__22091),
            .I(N__22088));
    InMux I__3152 (
            .O(N__22088),
            .I(N__22085));
    LocalMux I__3151 (
            .O(N__22085),
            .I(N__22082));
    Span4Mux_h I__3150 (
            .O(N__22082),
            .I(N__22079));
    Odrv4 I__3149 (
            .O(N__22079),
            .I(comm_buf_7_1));
    InMux I__3148 (
            .O(N__22076),
            .I(N__22073));
    LocalMux I__3147 (
            .O(N__22073),
            .I(N__22070));
    Span4Mux_v I__3146 (
            .O(N__22070),
            .I(N__22067));
    Span4Mux_h I__3145 (
            .O(N__22067),
            .I(N__22064));
    Odrv4 I__3144 (
            .O(N__22064),
            .I(comm_buf_3_4));
    InMux I__3143 (
            .O(N__22061),
            .I(N__22058));
    LocalMux I__3142 (
            .O(N__22058),
            .I(N__22055));
    Span4Mux_v I__3141 (
            .O(N__22055),
            .I(N__22052));
    Odrv4 I__3140 (
            .O(N__22052),
            .I(comm_buf_2_4));
    CascadeMux I__3139 (
            .O(N__22049),
            .I(n15403_cascade_));
    CascadeMux I__3138 (
            .O(N__22046),
            .I(n16479_cascade_));
    InMux I__3137 (
            .O(N__22043),
            .I(N__22040));
    LocalMux I__3136 (
            .O(N__22040),
            .I(N__22037));
    Span4Mux_v I__3135 (
            .O(N__22037),
            .I(N__22034));
    Span4Mux_h I__3134 (
            .O(N__22034),
            .I(N__22031));
    Sp12to4 I__3133 (
            .O(N__22031),
            .I(N__22028));
    Odrv12 I__3132 (
            .O(N__22028),
            .I(buf_data4_3));
    CascadeMux I__3131 (
            .O(N__22025),
            .I(N__22022));
    InMux I__3130 (
            .O(N__22022),
            .I(N__22019));
    LocalMux I__3129 (
            .O(N__22019),
            .I(N__22016));
    Span4Mux_h I__3128 (
            .O(N__22016),
            .I(N__22013));
    Odrv4 I__3127 (
            .O(N__22013),
            .I(comm_buf_11_3));
    InMux I__3126 (
            .O(N__22010),
            .I(N__22007));
    LocalMux I__3125 (
            .O(N__22007),
            .I(N__22004));
    Span4Mux_h I__3124 (
            .O(N__22004),
            .I(N__22001));
    Span4Mux_h I__3123 (
            .O(N__22001),
            .I(N__21998));
    Odrv4 I__3122 (
            .O(N__21998),
            .I(buf_data4_4));
    InMux I__3121 (
            .O(N__21995),
            .I(N__21992));
    LocalMux I__3120 (
            .O(N__21992),
            .I(N__21989));
    Span4Mux_h I__3119 (
            .O(N__21989),
            .I(N__21986));
    Odrv4 I__3118 (
            .O(N__21986),
            .I(buf_data4_5));
    CascadeMux I__3117 (
            .O(N__21983),
            .I(N__21980));
    InMux I__3116 (
            .O(N__21980),
            .I(N__21977));
    LocalMux I__3115 (
            .O(N__21977),
            .I(comm_buf_11_5));
    InMux I__3114 (
            .O(N__21974),
            .I(N__21971));
    LocalMux I__3113 (
            .O(N__21971),
            .I(N__21968));
    Span4Mux_h I__3112 (
            .O(N__21968),
            .I(N__21965));
    Span4Mux_h I__3111 (
            .O(N__21965),
            .I(N__21962));
    Odrv4 I__3110 (
            .O(N__21962),
            .I(buf_data4_6));
    InMux I__3109 (
            .O(N__21959),
            .I(N__21956));
    LocalMux I__3108 (
            .O(N__21956),
            .I(N__21953));
    Span4Mux_v I__3107 (
            .O(N__21953),
            .I(N__21950));
    Span4Mux_h I__3106 (
            .O(N__21950),
            .I(N__21947));
    Odrv4 I__3105 (
            .O(N__21947),
            .I(buf_data4_7));
    CascadeMux I__3104 (
            .O(N__21944),
            .I(N__21941));
    InMux I__3103 (
            .O(N__21941),
            .I(N__21938));
    LocalMux I__3102 (
            .O(N__21938),
            .I(N__21935));
    Odrv4 I__3101 (
            .O(N__21935),
            .I(comm_buf_11_7));
    InMux I__3100 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__3099 (
            .O(N__21929),
            .I(N__21926));
    Span4Mux_v I__3098 (
            .O(N__21926),
            .I(N__21923));
    Span4Mux_h I__3097 (
            .O(N__21923),
            .I(N__21920));
    Sp12to4 I__3096 (
            .O(N__21920),
            .I(N__21917));
    Odrv12 I__3095 (
            .O(N__21917),
            .I(buf_data4_0));
    InMux I__3094 (
            .O(N__21914),
            .I(N__21911));
    LocalMux I__3093 (
            .O(N__21911),
            .I(comm_buf_11_0));
    InMux I__3092 (
            .O(N__21908),
            .I(N__21905));
    LocalMux I__3091 (
            .O(N__21905),
            .I(N__21902));
    Span4Mux_h I__3090 (
            .O(N__21902),
            .I(N__21899));
    Span4Mux_h I__3089 (
            .O(N__21899),
            .I(N__21896));
    Span4Mux_h I__3088 (
            .O(N__21896),
            .I(N__21893));
    Span4Mux_v I__3087 (
            .O(N__21893),
            .I(N__21890));
    Odrv4 I__3086 (
            .O(N__21890),
            .I(buf_data3_15));
    InMux I__3085 (
            .O(N__21887),
            .I(N__21884));
    LocalMux I__3084 (
            .O(N__21884),
            .I(N__21881));
    Odrv4 I__3083 (
            .O(N__21881),
            .I(comm_buf_7_7));
    InMux I__3082 (
            .O(N__21878),
            .I(N__21875));
    LocalMux I__3081 (
            .O(N__21875),
            .I(N__21872));
    Sp12to4 I__3080 (
            .O(N__21872),
            .I(N__21869));
    Span12Mux_h I__3079 (
            .O(N__21869),
            .I(N__21866));
    Span12Mux_v I__3078 (
            .O(N__21866),
            .I(N__21863));
    Odrv12 I__3077 (
            .O(N__21863),
            .I(buf_data3_8));
    CascadeMux I__3076 (
            .O(N__21860),
            .I(N__21857));
    InMux I__3075 (
            .O(N__21857),
            .I(N__21854));
    LocalMux I__3074 (
            .O(N__21854),
            .I(N__21851));
    Odrv4 I__3073 (
            .O(N__21851),
            .I(comm_buf_7_0));
    InMux I__3072 (
            .O(N__21848),
            .I(N__21845));
    LocalMux I__3071 (
            .O(N__21845),
            .I(N__21842));
    Span4Mux_h I__3070 (
            .O(N__21842),
            .I(N__21839));
    Span4Mux_v I__3069 (
            .O(N__21839),
            .I(N__21836));
    Span4Mux_h I__3068 (
            .O(N__21836),
            .I(N__21833));
    Span4Mux_h I__3067 (
            .O(N__21833),
            .I(N__21830));
    Odrv4 I__3066 (
            .O(N__21830),
            .I(buf_data3_14));
    InMux I__3065 (
            .O(N__21827),
            .I(N__21824));
    LocalMux I__3064 (
            .O(N__21824),
            .I(N__21821));
    Odrv4 I__3063 (
            .O(N__21821),
            .I(comm_buf_3_7));
    InMux I__3062 (
            .O(N__21818),
            .I(N__21815));
    LocalMux I__3061 (
            .O(N__21815),
            .I(N__21812));
    Span12Mux_h I__3060 (
            .O(N__21812),
            .I(N__21809));
    Odrv12 I__3059 (
            .O(N__21809),
            .I(comm_buf_2_7));
    CascadeMux I__3058 (
            .O(N__21806),
            .I(n15382_cascade_));
    CascadeMux I__3057 (
            .O(N__21803),
            .I(n16383_cascade_));
    CascadeMux I__3056 (
            .O(N__21800),
            .I(n16494_cascade_));
    InMux I__3055 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__3054 (
            .O(N__21794),
            .I(n16497));
    InMux I__3053 (
            .O(N__21791),
            .I(N__21788));
    LocalMux I__3052 (
            .O(N__21788),
            .I(n15450));
    CascadeMux I__3051 (
            .O(N__21785),
            .I(n15451_cascade_));
    InMux I__3050 (
            .O(N__21782),
            .I(N__21779));
    LocalMux I__3049 (
            .O(N__21779),
            .I(n16380));
    InMux I__3048 (
            .O(N__21776),
            .I(N__21773));
    LocalMux I__3047 (
            .O(N__21773),
            .I(N__21770));
    Span12Mux_h I__3046 (
            .O(N__21770),
            .I(N__21767));
    Odrv12 I__3045 (
            .O(N__21767),
            .I(buf_data4_1));
    InMux I__3044 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__3043 (
            .O(N__21761),
            .I(N__21758));
    Span4Mux_h I__3042 (
            .O(N__21758),
            .I(N__21755));
    Span4Mux_h I__3041 (
            .O(N__21755),
            .I(N__21752));
    Span4Mux_h I__3040 (
            .O(N__21752),
            .I(N__21749));
    Odrv4 I__3039 (
            .O(N__21749),
            .I(buf_data4_2));
    CascadeMux I__3038 (
            .O(N__21746),
            .I(N__21743));
    InMux I__3037 (
            .O(N__21743),
            .I(N__21740));
    LocalMux I__3036 (
            .O(N__21740),
            .I(N__21737));
    Odrv4 I__3035 (
            .O(N__21737),
            .I(comm_buf_11_2));
    CascadeMux I__3034 (
            .O(N__21734),
            .I(N__21731));
    InMux I__3033 (
            .O(N__21731),
            .I(N__21728));
    LocalMux I__3032 (
            .O(N__21728),
            .I(N__21724));
    CascadeMux I__3031 (
            .O(N__21727),
            .I(N__21720));
    Span4Mux_v I__3030 (
            .O(N__21724),
            .I(N__21717));
    InMux I__3029 (
            .O(N__21723),
            .I(N__21712));
    InMux I__3028 (
            .O(N__21720),
            .I(N__21712));
    Odrv4 I__3027 (
            .O(N__21717),
            .I(cmd_rdadctmp_14));
    LocalMux I__3026 (
            .O(N__21712),
            .I(cmd_rdadctmp_14));
    InMux I__3025 (
            .O(N__21707),
            .I(N__21704));
    LocalMux I__3024 (
            .O(N__21704),
            .I(N__21701));
    Span4Mux_h I__3023 (
            .O(N__21701),
            .I(N__21698));
    Span4Mux_v I__3022 (
            .O(N__21698),
            .I(N__21695));
    Span4Mux_v I__3021 (
            .O(N__21695),
            .I(N__21691));
    InMux I__3020 (
            .O(N__21694),
            .I(N__21688));
    Span4Mux_h I__3019 (
            .O(N__21691),
            .I(N__21685));
    LocalMux I__3018 (
            .O(N__21688),
            .I(buf_adcdata1_6));
    Odrv4 I__3017 (
            .O(N__21685),
            .I(buf_adcdata1_6));
    CascadeMux I__3016 (
            .O(N__21680),
            .I(N__21677));
    InMux I__3015 (
            .O(N__21677),
            .I(N__21673));
    InMux I__3014 (
            .O(N__21676),
            .I(N__21670));
    LocalMux I__3013 (
            .O(N__21673),
            .I(N__21667));
    LocalMux I__3012 (
            .O(N__21670),
            .I(N__21664));
    Span4Mux_h I__3011 (
            .O(N__21667),
            .I(N__21658));
    Span4Mux_v I__3010 (
            .O(N__21664),
            .I(N__21658));
    InMux I__3009 (
            .O(N__21663),
            .I(N__21655));
    Odrv4 I__3008 (
            .O(N__21658),
            .I(cmd_rdadctmp_15_adj_1097));
    LocalMux I__3007 (
            .O(N__21655),
            .I(cmd_rdadctmp_15_adj_1097));
    IoInMux I__3006 (
            .O(N__21650),
            .I(N__21647));
    LocalMux I__3005 (
            .O(N__21647),
            .I(N__21644));
    IoSpan4Mux I__3004 (
            .O(N__21644),
            .I(N__21641));
    Span4Mux_s2_v I__3003 (
            .O(N__21641),
            .I(N__21638));
    Span4Mux_h I__3002 (
            .O(N__21638),
            .I(N__21635));
    Sp12to4 I__3001 (
            .O(N__21635),
            .I(N__21631));
    CascadeMux I__3000 (
            .O(N__21634),
            .I(N__21628));
    Span12Mux_s9_v I__2999 (
            .O(N__21631),
            .I(N__21625));
    InMux I__2998 (
            .O(N__21628),
            .I(N__21622));
    Odrv12 I__2997 (
            .O(N__21625),
            .I(M_SCLK4));
    LocalMux I__2996 (
            .O(N__21622),
            .I(M_SCLK4));
    InMux I__2995 (
            .O(N__21617),
            .I(N__21614));
    LocalMux I__2994 (
            .O(N__21614),
            .I(N__21611));
    Span4Mux_h I__2993 (
            .O(N__21611),
            .I(N__21607));
    InMux I__2992 (
            .O(N__21610),
            .I(N__21604));
    Odrv4 I__2991 (
            .O(N__21607),
            .I(\comm_spi.n10434 ));
    LocalMux I__2990 (
            .O(N__21604),
            .I(\comm_spi.n10434 ));
    InMux I__2989 (
            .O(N__21599),
            .I(N__21594));
    InMux I__2988 (
            .O(N__21598),
            .I(N__21589));
    InMux I__2987 (
            .O(N__21597),
            .I(N__21589));
    LocalMux I__2986 (
            .O(N__21594),
            .I(N__21586));
    LocalMux I__2985 (
            .O(N__21589),
            .I(comm_tx_buf_0));
    Odrv12 I__2984 (
            .O(N__21586),
            .I(comm_tx_buf_0));
    SRMux I__2983 (
            .O(N__21581),
            .I(N__21578));
    LocalMux I__2982 (
            .O(N__21578),
            .I(N__21575));
    Odrv12 I__2981 (
            .O(N__21575),
            .I(\comm_spi.data_tx_7__N_834 ));
    InMux I__2980 (
            .O(N__21572),
            .I(N__21569));
    LocalMux I__2979 (
            .O(N__21569),
            .I(n16428));
    InMux I__2978 (
            .O(N__21566),
            .I(N__21563));
    LocalMux I__2977 (
            .O(N__21563),
            .I(N__21560));
    Span12Mux_v I__2976 (
            .O(N__21560),
            .I(N__21557));
    Odrv12 I__2975 (
            .O(N__21557),
            .I(buf_data2_20));
    InMux I__2974 (
            .O(N__21554),
            .I(N__21551));
    LocalMux I__2973 (
            .O(N__21551),
            .I(N__21548));
    Span4Mux_v I__2972 (
            .O(N__21548),
            .I(N__21545));
    Odrv4 I__2971 (
            .O(N__21545),
            .I(n4104));
    CascadeMux I__2970 (
            .O(N__21542),
            .I(\ADC_VAC2.n17_cascade_ ));
    InMux I__2969 (
            .O(N__21539),
            .I(N__21535));
    CascadeMux I__2968 (
            .O(N__21538),
            .I(N__21532));
    LocalMux I__2967 (
            .O(N__21535),
            .I(N__21529));
    InMux I__2966 (
            .O(N__21532),
            .I(N__21526));
    Odrv4 I__2965 (
            .O(N__21529),
            .I(cmd_rdadctmp_2_adj_1110));
    LocalMux I__2964 (
            .O(N__21526),
            .I(cmd_rdadctmp_2_adj_1110));
    InMux I__2963 (
            .O(N__21521),
            .I(N__21517));
    CascadeMux I__2962 (
            .O(N__21520),
            .I(N__21514));
    LocalMux I__2961 (
            .O(N__21517),
            .I(N__21511));
    InMux I__2960 (
            .O(N__21514),
            .I(N__21508));
    Odrv4 I__2959 (
            .O(N__21511),
            .I(cmd_rdadctmp_3_adj_1109));
    LocalMux I__2958 (
            .O(N__21508),
            .I(cmd_rdadctmp_3_adj_1109));
    CascadeMux I__2957 (
            .O(N__21503),
            .I(N__21499));
    CascadeMux I__2956 (
            .O(N__21502),
            .I(N__21496));
    InMux I__2955 (
            .O(N__21499),
            .I(N__21493));
    InMux I__2954 (
            .O(N__21496),
            .I(N__21490));
    LocalMux I__2953 (
            .O(N__21493),
            .I(N__21487));
    LocalMux I__2952 (
            .O(N__21490),
            .I(acadc_dtrig2));
    Odrv4 I__2951 (
            .O(N__21487),
            .I(acadc_dtrig2));
    InMux I__2950 (
            .O(N__21482),
            .I(N__21478));
    InMux I__2949 (
            .O(N__21481),
            .I(N__21475));
    LocalMux I__2948 (
            .O(N__21478),
            .I(acadc_dtrig1));
    LocalMux I__2947 (
            .O(N__21475),
            .I(acadc_dtrig1));
    InMux I__2946 (
            .O(N__21470),
            .I(N__21464));
    InMux I__2945 (
            .O(N__21469),
            .I(N__21464));
    LocalMux I__2944 (
            .O(N__21464),
            .I(acadc_dtrig4));
    InMux I__2943 (
            .O(N__21461),
            .I(N__21455));
    InMux I__2942 (
            .O(N__21460),
            .I(N__21455));
    LocalMux I__2941 (
            .O(N__21455),
            .I(acadc_dtrig3));
    InMux I__2940 (
            .O(N__21452),
            .I(\ADC_VAC2.n13991 ));
    InMux I__2939 (
            .O(N__21449),
            .I(\ADC_VAC2.n13992 ));
    InMux I__2938 (
            .O(N__21446),
            .I(\ADC_VAC2.n13993 ));
    InMux I__2937 (
            .O(N__21443),
            .I(\ADC_VAC2.n13994 ));
    InMux I__2936 (
            .O(N__21440),
            .I(N__21436));
    InMux I__2935 (
            .O(N__21439),
            .I(N__21433));
    LocalMux I__2934 (
            .O(N__21436),
            .I(\ADC_VAC2.bit_cnt_1 ));
    LocalMux I__2933 (
            .O(N__21433),
            .I(\ADC_VAC2.bit_cnt_1 ));
    CascadeMux I__2932 (
            .O(N__21428),
            .I(N__21424));
    InMux I__2931 (
            .O(N__21427),
            .I(N__21421));
    InMux I__2930 (
            .O(N__21424),
            .I(N__21418));
    LocalMux I__2929 (
            .O(N__21421),
            .I(\ADC_VAC2.bit_cnt_7 ));
    LocalMux I__2928 (
            .O(N__21418),
            .I(\ADC_VAC2.bit_cnt_7 ));
    CascadeMux I__2927 (
            .O(N__21413),
            .I(\ADC_VAC2.n15261_cascade_ ));
    InMux I__2926 (
            .O(N__21410),
            .I(N__21407));
    LocalMux I__2925 (
            .O(N__21407),
            .I(\ADC_VAC2.n15595 ));
    CEMux I__2924 (
            .O(N__21404),
            .I(N__21401));
    LocalMux I__2923 (
            .O(N__21401),
            .I(\ADC_VAC2.n15262 ));
    CascadeMux I__2922 (
            .O(N__21398),
            .I(N__21394));
    InMux I__2921 (
            .O(N__21397),
            .I(N__21391));
    InMux I__2920 (
            .O(N__21394),
            .I(N__21388));
    LocalMux I__2919 (
            .O(N__21391),
            .I(\ADC_VAC2.bit_cnt_6 ));
    LocalMux I__2918 (
            .O(N__21388),
            .I(\ADC_VAC2.bit_cnt_6 ));
    InMux I__2917 (
            .O(N__21383),
            .I(N__21379));
    InMux I__2916 (
            .O(N__21382),
            .I(N__21376));
    LocalMux I__2915 (
            .O(N__21379),
            .I(\ADC_VAC2.bit_cnt_0 ));
    LocalMux I__2914 (
            .O(N__21376),
            .I(\ADC_VAC2.bit_cnt_0 ));
    InMux I__2913 (
            .O(N__21371),
            .I(N__21368));
    LocalMux I__2912 (
            .O(N__21368),
            .I(\ADC_VAC2.n16 ));
    InMux I__2911 (
            .O(N__21365),
            .I(N__21362));
    LocalMux I__2910 (
            .O(N__21362),
            .I(N__21359));
    Span4Mux_v I__2909 (
            .O(N__21359),
            .I(N__21356));
    Sp12to4 I__2908 (
            .O(N__21356),
            .I(N__21352));
    CascadeMux I__2907 (
            .O(N__21355),
            .I(N__21349));
    Span12Mux_h I__2906 (
            .O(N__21352),
            .I(N__21346));
    InMux I__2905 (
            .O(N__21349),
            .I(N__21343));
    Span12Mux_v I__2904 (
            .O(N__21346),
            .I(N__21340));
    LocalMux I__2903 (
            .O(N__21343),
            .I(buf_adcdata1_22));
    Odrv12 I__2902 (
            .O(N__21340),
            .I(buf_adcdata1_22));
    CascadeMux I__2901 (
            .O(N__21335),
            .I(N__21332));
    InMux I__2900 (
            .O(N__21332),
            .I(N__21328));
    CascadeMux I__2899 (
            .O(N__21331),
            .I(N__21324));
    LocalMux I__2898 (
            .O(N__21328),
            .I(N__21321));
    InMux I__2897 (
            .O(N__21327),
            .I(N__21318));
    InMux I__2896 (
            .O(N__21324),
            .I(N__21315));
    Odrv4 I__2895 (
            .O(N__21321),
            .I(cmd_rdadctmp_24_adj_1052));
    LocalMux I__2894 (
            .O(N__21318),
            .I(cmd_rdadctmp_24_adj_1052));
    LocalMux I__2893 (
            .O(N__21315),
            .I(cmd_rdadctmp_24_adj_1052));
    InMux I__2892 (
            .O(N__21308),
            .I(N__21305));
    LocalMux I__2891 (
            .O(N__21305),
            .I(N__21301));
    InMux I__2890 (
            .O(N__21304),
            .I(N__21298));
    Span12Mux_h I__2889 (
            .O(N__21301),
            .I(N__21295));
    LocalMux I__2888 (
            .O(N__21298),
            .I(buf_adcdata2_16));
    Odrv12 I__2887 (
            .O(N__21295),
            .I(buf_adcdata2_16));
    InMux I__2886 (
            .O(N__21290),
            .I(N__21283));
    InMux I__2885 (
            .O(N__21289),
            .I(N__21283));
    InMux I__2884 (
            .O(N__21288),
            .I(N__21280));
    LocalMux I__2883 (
            .O(N__21283),
            .I(cmd_rdadctmp_29));
    LocalMux I__2882 (
            .O(N__21280),
            .I(cmd_rdadctmp_29));
    CascadeMux I__2881 (
            .O(N__21275),
            .I(N__21270));
    InMux I__2880 (
            .O(N__21274),
            .I(N__21263));
    InMux I__2879 (
            .O(N__21273),
            .I(N__21263));
    InMux I__2878 (
            .O(N__21270),
            .I(N__21263));
    LocalMux I__2877 (
            .O(N__21263),
            .I(cmd_rdadctmp_30));
    InMux I__2876 (
            .O(N__21260),
            .I(N__21257));
    LocalMux I__2875 (
            .O(N__21257),
            .I(N__21254));
    Span4Mux_h I__2874 (
            .O(N__21254),
            .I(N__21251));
    Sp12to4 I__2873 (
            .O(N__21251),
            .I(N__21247));
    InMux I__2872 (
            .O(N__21250),
            .I(N__21244));
    Span12Mux_v I__2871 (
            .O(N__21247),
            .I(N__21241));
    LocalMux I__2870 (
            .O(N__21244),
            .I(buf_adcdata1_1));
    Odrv12 I__2869 (
            .O(N__21241),
            .I(buf_adcdata1_1));
    InMux I__2868 (
            .O(N__21236),
            .I(bfn_9_13_0_));
    InMux I__2867 (
            .O(N__21233),
            .I(\ADC_VAC2.n13988 ));
    InMux I__2866 (
            .O(N__21230),
            .I(\ADC_VAC2.n13989 ));
    InMux I__2865 (
            .O(N__21227),
            .I(\ADC_VAC2.n13990 ));
    IoInMux I__2864 (
            .O(N__21224),
            .I(N__21221));
    LocalMux I__2863 (
            .O(N__21221),
            .I(N__21218));
    Span12Mux_s3_v I__2862 (
            .O(N__21218),
            .I(N__21215));
    Span12Mux_v I__2861 (
            .O(N__21215),
            .I(N__21211));
    InMux I__2860 (
            .O(N__21214),
            .I(N__21208));
    Odrv12 I__2859 (
            .O(N__21211),
            .I(DDS_MOSI1));
    LocalMux I__2858 (
            .O(N__21208),
            .I(DDS_MOSI1));
    InMux I__2857 (
            .O(N__21203),
            .I(N__21200));
    LocalMux I__2856 (
            .O(N__21200),
            .I(n15522));
    CascadeMux I__2855 (
            .O(N__21197),
            .I(N__21194));
    InMux I__2854 (
            .O(N__21194),
            .I(N__21191));
    LocalMux I__2853 (
            .O(N__21191),
            .I(n15523));
    CascadeMux I__2852 (
            .O(N__21188),
            .I(n16398_cascade_));
    CascadeMux I__2851 (
            .O(N__21185),
            .I(n16401_cascade_));
    CascadeMux I__2850 (
            .O(N__21182),
            .I(n109_adj_1155_cascade_));
    CascadeMux I__2849 (
            .O(N__21179),
            .I(n8048_cascade_));
    InMux I__2848 (
            .O(N__21176),
            .I(N__21173));
    LocalMux I__2847 (
            .O(N__21173),
            .I(N__21170));
    Odrv4 I__2846 (
            .O(N__21170),
            .I(n15578));
    InMux I__2845 (
            .O(N__21167),
            .I(N__21164));
    LocalMux I__2844 (
            .O(N__21164),
            .I(N__21161));
    Sp12to4 I__2843 (
            .O(N__21161),
            .I(N__21158));
    Span12Mux_v I__2842 (
            .O(N__21158),
            .I(N__21154));
    CascadeMux I__2841 (
            .O(N__21157),
            .I(N__21151));
    Span12Mux_v I__2840 (
            .O(N__21154),
            .I(N__21148));
    InMux I__2839 (
            .O(N__21151),
            .I(N__21145));
    Span12Mux_h I__2838 (
            .O(N__21148),
            .I(N__21142));
    LocalMux I__2837 (
            .O(N__21145),
            .I(buf_adcdata1_21));
    Odrv12 I__2836 (
            .O(N__21142),
            .I(buf_adcdata1_21));
    InMux I__2835 (
            .O(N__21137),
            .I(N__21134));
    LocalMux I__2834 (
            .O(N__21134),
            .I(N__21131));
    Span4Mux_v I__2833 (
            .O(N__21131),
            .I(N__21128));
    Odrv4 I__2832 (
            .O(N__21128),
            .I(comm_buf_3_7_N_501_2));
    InMux I__2831 (
            .O(N__21125),
            .I(N__21122));
    LocalMux I__2830 (
            .O(N__21122),
            .I(N__21119));
    Odrv4 I__2829 (
            .O(N__21119),
            .I(comm_buf_3_2));
    InMux I__2828 (
            .O(N__21116),
            .I(N__21113));
    LocalMux I__2827 (
            .O(N__21113),
            .I(N__21110));
    Span4Mux_h I__2826 (
            .O(N__21110),
            .I(N__21107));
    Odrv4 I__2825 (
            .O(N__21107),
            .I(comm_buf_3_3));
    InMux I__2824 (
            .O(N__21104),
            .I(N__21101));
    LocalMux I__2823 (
            .O(N__21101),
            .I(N__21098));
    Span12Mux_h I__2822 (
            .O(N__21098),
            .I(N__21095));
    Odrv12 I__2821 (
            .O(N__21095),
            .I(buf_data4_19));
    InMux I__2820 (
            .O(N__21092),
            .I(N__21089));
    LocalMux I__2819 (
            .O(N__21089),
            .I(N__21086));
    Span4Mux_v I__2818 (
            .O(N__21086),
            .I(N__21083));
    Sp12to4 I__2817 (
            .O(N__21083),
            .I(N__21080));
    Odrv12 I__2816 (
            .O(N__21080),
            .I(comm_buf_9_3));
    InMux I__2815 (
            .O(N__21077),
            .I(N__21074));
    LocalMux I__2814 (
            .O(N__21074),
            .I(N__21071));
    Span12Mux_v I__2813 (
            .O(N__21071),
            .I(N__21068));
    Span12Mux_h I__2812 (
            .O(N__21068),
            .I(N__21065));
    Odrv12 I__2811 (
            .O(N__21065),
            .I(buf_data4_20));
    CascadeMux I__2810 (
            .O(N__21062),
            .I(n66_adj_1153_cascade_));
    IoInMux I__2809 (
            .O(N__21059),
            .I(N__21056));
    LocalMux I__2808 (
            .O(N__21056),
            .I(N__21053));
    IoSpan4Mux I__2807 (
            .O(N__21053),
            .I(N__21050));
    IoSpan4Mux I__2806 (
            .O(N__21050),
            .I(N__21047));
    Sp12to4 I__2805 (
            .O(N__21047),
            .I(N__21043));
    CascadeMux I__2804 (
            .O(N__21046),
            .I(N__21040));
    Span12Mux_s7_v I__2803 (
            .O(N__21043),
            .I(N__21037));
    InMux I__2802 (
            .O(N__21040),
            .I(N__21034));
    Odrv12 I__2801 (
            .O(N__21037),
            .I(DDS_SCK1));
    LocalMux I__2800 (
            .O(N__21034),
            .I(DDS_SCK1));
    InMux I__2799 (
            .O(N__21029),
            .I(N__21026));
    LocalMux I__2798 (
            .O(N__21026),
            .I(N__21023));
    Span4Mux_h I__2797 (
            .O(N__21023),
            .I(N__21020));
    Odrv4 I__2796 (
            .O(N__21020),
            .I(n16431));
    InMux I__2795 (
            .O(N__21017),
            .I(N__21014));
    LocalMux I__2794 (
            .O(N__21014),
            .I(N__21011));
    Span4Mux_v I__2793 (
            .O(N__21011),
            .I(N__21008));
    Odrv4 I__2792 (
            .O(N__21008),
            .I(comm_buf_4_0));
    CascadeMux I__2791 (
            .O(N__21005),
            .I(n16506_cascade_));
    InMux I__2790 (
            .O(N__21002),
            .I(N__20999));
    LocalMux I__2789 (
            .O(N__20999),
            .I(N__20996));
    Span4Mux_v I__2788 (
            .O(N__20996),
            .I(N__20993));
    Odrv4 I__2787 (
            .O(N__20993),
            .I(comm_buf_5_0));
    CascadeMux I__2786 (
            .O(N__20990),
            .I(N__20987));
    InMux I__2785 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__2784 (
            .O(N__20984),
            .I(n16509));
    InMux I__2783 (
            .O(N__20981),
            .I(N__20978));
    LocalMux I__2782 (
            .O(N__20978),
            .I(N__20975));
    Span4Mux_v I__2781 (
            .O(N__20975),
            .I(N__20972));
    Odrv4 I__2780 (
            .O(N__20972),
            .I(n15424));
    CascadeMux I__2779 (
            .O(N__20969),
            .I(N__20966));
    InMux I__2778 (
            .O(N__20966),
            .I(N__20963));
    LocalMux I__2777 (
            .O(N__20963),
            .I(n15412));
    InMux I__2776 (
            .O(N__20960),
            .I(N__20957));
    LocalMux I__2775 (
            .O(N__20957),
            .I(N__20954));
    Odrv12 I__2774 (
            .O(N__20954),
            .I(comm_buf_5_7));
    InMux I__2773 (
            .O(N__20951),
            .I(N__20948));
    LocalMux I__2772 (
            .O(N__20948),
            .I(N__20945));
    Span4Mux_h I__2771 (
            .O(N__20945),
            .I(N__20942));
    Odrv4 I__2770 (
            .O(N__20942),
            .I(comm_buf_4_7));
    CascadeMux I__2769 (
            .O(N__20939),
            .I(n16482_cascade_));
    InMux I__2768 (
            .O(N__20936),
            .I(N__20933));
    LocalMux I__2767 (
            .O(N__20933),
            .I(N__20930));
    Span4Mux_h I__2766 (
            .O(N__20930),
            .I(N__20927));
    Odrv4 I__2765 (
            .O(N__20927),
            .I(n16485));
    InMux I__2764 (
            .O(N__20924),
            .I(N__20920));
    InMux I__2763 (
            .O(N__20923),
            .I(N__20917));
    LocalMux I__2762 (
            .O(N__20920),
            .I(\comm_spi.n16911 ));
    LocalMux I__2761 (
            .O(N__20917),
            .I(\comm_spi.n16911 ));
    InMux I__2760 (
            .O(N__20912),
            .I(N__20908));
    InMux I__2759 (
            .O(N__20911),
            .I(N__20905));
    LocalMux I__2758 (
            .O(N__20908),
            .I(\comm_spi.n10433 ));
    LocalMux I__2757 (
            .O(N__20905),
            .I(\comm_spi.n10433 ));
    CascadeMux I__2756 (
            .O(N__20900),
            .I(\comm_spi.n16911_cascade_ ));
    SRMux I__2755 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__2754 (
            .O(N__20894),
            .I(N__20891));
    Span4Mux_v I__2753 (
            .O(N__20891),
            .I(N__20888));
    Odrv4 I__2752 (
            .O(N__20888),
            .I(\comm_spi.data_tx_7__N_811 ));
    SRMux I__2751 (
            .O(N__20885),
            .I(N__20882));
    LocalMux I__2750 (
            .O(N__20882),
            .I(N__20879));
    Odrv12 I__2749 (
            .O(N__20879),
            .I(\comm_spi.data_tx_7__N_831 ));
    SRMux I__2748 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__2747 (
            .O(N__20873),
            .I(\comm_spi.data_tx_7__N_812 ));
    InMux I__2746 (
            .O(N__20870),
            .I(N__20861));
    InMux I__2745 (
            .O(N__20869),
            .I(N__20861));
    InMux I__2744 (
            .O(N__20868),
            .I(N__20861));
    LocalMux I__2743 (
            .O(N__20861),
            .I(N__20858));
    Span4Mux_v I__2742 (
            .O(N__20858),
            .I(N__20855));
    Odrv4 I__2741 (
            .O(N__20855),
            .I(comm_tx_buf_1));
    InMux I__2740 (
            .O(N__20852),
            .I(N__20849));
    LocalMux I__2739 (
            .O(N__20849),
            .I(n15411));
    CascadeMux I__2738 (
            .O(N__20846),
            .I(n16446_cascade_));
    InMux I__2737 (
            .O(N__20843),
            .I(N__20840));
    LocalMux I__2736 (
            .O(N__20840),
            .I(n15391));
    InMux I__2735 (
            .O(N__20837),
            .I(N__20834));
    LocalMux I__2734 (
            .O(N__20834),
            .I(n16449));
    InMux I__2733 (
            .O(N__20831),
            .I(N__20828));
    LocalMux I__2732 (
            .O(N__20828),
            .I(N__20825));
    Span12Mux_h I__2731 (
            .O(N__20825),
            .I(N__20822));
    Odrv12 I__2730 (
            .O(N__20822),
            .I(buf_data2_3));
    InMux I__2729 (
            .O(N__20819),
            .I(N__20815));
    CascadeMux I__2728 (
            .O(N__20818),
            .I(N__20812));
    LocalMux I__2727 (
            .O(N__20815),
            .I(N__20808));
    InMux I__2726 (
            .O(N__20812),
            .I(N__20805));
    InMux I__2725 (
            .O(N__20811),
            .I(N__20802));
    Span12Mux_h I__2724 (
            .O(N__20808),
            .I(N__20797));
    LocalMux I__2723 (
            .O(N__20805),
            .I(N__20797));
    LocalMux I__2722 (
            .O(N__20802),
            .I(buf_adcdata4_3));
    Odrv12 I__2721 (
            .O(N__20797),
            .I(buf_adcdata4_3));
    InMux I__2720 (
            .O(N__20792),
            .I(N__20789));
    LocalMux I__2719 (
            .O(N__20789),
            .I(N__20786));
    Span4Mux_h I__2718 (
            .O(N__20786),
            .I(N__20783));
    Odrv4 I__2717 (
            .O(N__20783),
            .I(n4305));
    CascadeMux I__2716 (
            .O(N__20780),
            .I(N__20777));
    InMux I__2715 (
            .O(N__20777),
            .I(N__20774));
    LocalMux I__2714 (
            .O(N__20774),
            .I(N__20771));
    Span4Mux_v I__2713 (
            .O(N__20771),
            .I(N__20768));
    Sp12to4 I__2712 (
            .O(N__20768),
            .I(N__20765));
    Span12Mux_h I__2711 (
            .O(N__20765),
            .I(N__20762));
    Odrv12 I__2710 (
            .O(N__20762),
            .I(M_MISO3));
    InMux I__2709 (
            .O(N__20759),
            .I(N__20753));
    InMux I__2708 (
            .O(N__20758),
            .I(N__20753));
    LocalMux I__2707 (
            .O(N__20753),
            .I(cmd_rdadctmp_0_adj_1112));
    CascadeMux I__2706 (
            .O(N__20750),
            .I(N__20746));
    InMux I__2705 (
            .O(N__20749),
            .I(N__20743));
    InMux I__2704 (
            .O(N__20746),
            .I(N__20740));
    LocalMux I__2703 (
            .O(N__20743),
            .I(cmd_rdadctmp_1_adj_1111));
    LocalMux I__2702 (
            .O(N__20740),
            .I(cmd_rdadctmp_1_adj_1111));
    CEMux I__2701 (
            .O(N__20735),
            .I(N__20732));
    LocalMux I__2700 (
            .O(N__20732),
            .I(N__20729));
    Span4Mux_v I__2699 (
            .O(N__20729),
            .I(N__20726));
    Odrv4 I__2698 (
            .O(N__20726),
            .I(\ADC_VAC3.n12 ));
    InMux I__2697 (
            .O(N__20723),
            .I(N__20720));
    LocalMux I__2696 (
            .O(N__20720),
            .I(N__20717));
    Odrv4 I__2695 (
            .O(N__20717),
            .I(n15162));
    CascadeMux I__2694 (
            .O(N__20714),
            .I(n15162_cascade_));
    CascadeMux I__2693 (
            .O(N__20711),
            .I(n14_adj_1031_cascade_));
    IoInMux I__2692 (
            .O(N__20708),
            .I(N__20705));
    LocalMux I__2691 (
            .O(N__20705),
            .I(N__20702));
    Span4Mux_s0_v I__2690 (
            .O(N__20702),
            .I(N__20699));
    Sp12to4 I__2689 (
            .O(N__20699),
            .I(N__20696));
    Span12Mux_s11_h I__2688 (
            .O(N__20696),
            .I(N__20692));
    CascadeMux I__2687 (
            .O(N__20695),
            .I(N__20689));
    Span12Mux_v I__2686 (
            .O(N__20692),
            .I(N__20686));
    InMux I__2685 (
            .O(N__20689),
            .I(N__20683));
    Odrv12 I__2684 (
            .O(N__20686),
            .I(M_CS3));
    LocalMux I__2683 (
            .O(N__20683),
            .I(M_CS3));
    IoInMux I__2682 (
            .O(N__20678),
            .I(N__20675));
    LocalMux I__2681 (
            .O(N__20675),
            .I(N__20671));
    CascadeMux I__2680 (
            .O(N__20674),
            .I(N__20668));
    Span12Mux_s11_v I__2679 (
            .O(N__20671),
            .I(N__20665));
    InMux I__2678 (
            .O(N__20668),
            .I(N__20662));
    Odrv12 I__2677 (
            .O(N__20665),
            .I(M_SCLK3));
    LocalMux I__2676 (
            .O(N__20662),
            .I(M_SCLK3));
    InMux I__2675 (
            .O(N__20657),
            .I(N__20651));
    InMux I__2674 (
            .O(N__20656),
            .I(N__20651));
    LocalMux I__2673 (
            .O(N__20651),
            .I(cmd_rdadctmp_4_adj_1108));
    InMux I__2672 (
            .O(N__20648),
            .I(N__20645));
    LocalMux I__2671 (
            .O(N__20645),
            .I(N__20639));
    CascadeMux I__2670 (
            .O(N__20644),
            .I(N__20633));
    CascadeMux I__2669 (
            .O(N__20643),
            .I(N__20628));
    CascadeMux I__2668 (
            .O(N__20642),
            .I(N__20624));
    Span4Mux_h I__2667 (
            .O(N__20639),
            .I(N__20619));
    InMux I__2666 (
            .O(N__20638),
            .I(N__20612));
    InMux I__2665 (
            .O(N__20637),
            .I(N__20612));
    InMux I__2664 (
            .O(N__20636),
            .I(N__20612));
    InMux I__2663 (
            .O(N__20633),
            .I(N__20605));
    InMux I__2662 (
            .O(N__20632),
            .I(N__20605));
    InMux I__2661 (
            .O(N__20631),
            .I(N__20605));
    InMux I__2660 (
            .O(N__20628),
            .I(N__20594));
    InMux I__2659 (
            .O(N__20627),
            .I(N__20594));
    InMux I__2658 (
            .O(N__20624),
            .I(N__20594));
    InMux I__2657 (
            .O(N__20623),
            .I(N__20594));
    InMux I__2656 (
            .O(N__20622),
            .I(N__20594));
    Odrv4 I__2655 (
            .O(N__20619),
            .I(DTRIG_N_957));
    LocalMux I__2654 (
            .O(N__20612),
            .I(DTRIG_N_957));
    LocalMux I__2653 (
            .O(N__20605),
            .I(DTRIG_N_957));
    LocalMux I__2652 (
            .O(N__20594),
            .I(DTRIG_N_957));
    InMux I__2651 (
            .O(N__20585),
            .I(N__20582));
    LocalMux I__2650 (
            .O(N__20582),
            .I(N__20577));
    CascadeMux I__2649 (
            .O(N__20581),
            .I(N__20570));
    InMux I__2648 (
            .O(N__20580),
            .I(N__20562));
    Span4Mux_v I__2647 (
            .O(N__20577),
            .I(N__20559));
    InMux I__2646 (
            .O(N__20576),
            .I(N__20552));
    InMux I__2645 (
            .O(N__20575),
            .I(N__20552));
    InMux I__2644 (
            .O(N__20574),
            .I(N__20552));
    InMux I__2643 (
            .O(N__20573),
            .I(N__20547));
    InMux I__2642 (
            .O(N__20570),
            .I(N__20547));
    InMux I__2641 (
            .O(N__20569),
            .I(N__20536));
    InMux I__2640 (
            .O(N__20568),
            .I(N__20536));
    InMux I__2639 (
            .O(N__20567),
            .I(N__20536));
    InMux I__2638 (
            .O(N__20566),
            .I(N__20536));
    InMux I__2637 (
            .O(N__20565),
            .I(N__20536));
    LocalMux I__2636 (
            .O(N__20562),
            .I(adc_state_1));
    Odrv4 I__2635 (
            .O(N__20559),
            .I(adc_state_1));
    LocalMux I__2634 (
            .O(N__20552),
            .I(adc_state_1));
    LocalMux I__2633 (
            .O(N__20547),
            .I(adc_state_1));
    LocalMux I__2632 (
            .O(N__20536),
            .I(adc_state_1));
    CascadeMux I__2631 (
            .O(N__20525),
            .I(N__20522));
    InMux I__2630 (
            .O(N__20522),
            .I(N__20519));
    LocalMux I__2629 (
            .O(N__20519),
            .I(N__20515));
    CascadeMux I__2628 (
            .O(N__20518),
            .I(N__20511));
    Span4Mux_v I__2627 (
            .O(N__20515),
            .I(N__20508));
    InMux I__2626 (
            .O(N__20514),
            .I(N__20505));
    InMux I__2625 (
            .O(N__20511),
            .I(N__20502));
    Odrv4 I__2624 (
            .O(N__20508),
            .I(cmd_rdadctmp_11));
    LocalMux I__2623 (
            .O(N__20505),
            .I(cmd_rdadctmp_11));
    LocalMux I__2622 (
            .O(N__20502),
            .I(cmd_rdadctmp_11));
    InMux I__2621 (
            .O(N__20495),
            .I(N__20492));
    LocalMux I__2620 (
            .O(N__20492),
            .I(N__20488));
    CascadeMux I__2619 (
            .O(N__20491),
            .I(N__20485));
    Span4Mux_v I__2618 (
            .O(N__20488),
            .I(N__20482));
    InMux I__2617 (
            .O(N__20485),
            .I(N__20478));
    Sp12to4 I__2616 (
            .O(N__20482),
            .I(N__20475));
    InMux I__2615 (
            .O(N__20481),
            .I(N__20472));
    LocalMux I__2614 (
            .O(N__20478),
            .I(N__20469));
    Span12Mux_h I__2613 (
            .O(N__20475),
            .I(N__20466));
    LocalMux I__2612 (
            .O(N__20472),
            .I(buf_adcdata4_12));
    Odrv12 I__2611 (
            .O(N__20469),
            .I(buf_adcdata4_12));
    Odrv12 I__2610 (
            .O(N__20466),
            .I(buf_adcdata4_12));
    CascadeMux I__2609 (
            .O(N__20459),
            .I(N__20455));
    InMux I__2608 (
            .O(N__20458),
            .I(N__20452));
    InMux I__2607 (
            .O(N__20455),
            .I(N__20449));
    LocalMux I__2606 (
            .O(N__20452),
            .I(N__20446));
    LocalMux I__2605 (
            .O(N__20449),
            .I(N__20442));
    Span4Mux_v I__2604 (
            .O(N__20446),
            .I(N__20439));
    CascadeMux I__2603 (
            .O(N__20445),
            .I(N__20436));
    Span4Mux_h I__2602 (
            .O(N__20442),
            .I(N__20433));
    Span4Mux_v I__2601 (
            .O(N__20439),
            .I(N__20430));
    InMux I__2600 (
            .O(N__20436),
            .I(N__20427));
    Odrv4 I__2599 (
            .O(N__20433),
            .I(cmd_rdadctmp_16_adj_1060));
    Odrv4 I__2598 (
            .O(N__20430),
            .I(cmd_rdadctmp_16_adj_1060));
    LocalMux I__2597 (
            .O(N__20427),
            .I(cmd_rdadctmp_16_adj_1060));
    InMux I__2596 (
            .O(N__20420),
            .I(N__20417));
    LocalMux I__2595 (
            .O(N__20417),
            .I(N__20414));
    Span4Mux_v I__2594 (
            .O(N__20414),
            .I(N__20411));
    Sp12to4 I__2593 (
            .O(N__20411),
            .I(N__20407));
    InMux I__2592 (
            .O(N__20410),
            .I(N__20404));
    Span12Mux_h I__2591 (
            .O(N__20407),
            .I(N__20401));
    LocalMux I__2590 (
            .O(N__20404),
            .I(buf_adcdata2_8));
    Odrv12 I__2589 (
            .O(N__20401),
            .I(buf_adcdata2_8));
    CascadeMux I__2588 (
            .O(N__20396),
            .I(N__20393));
    InMux I__2587 (
            .O(N__20393),
            .I(N__20388));
    InMux I__2586 (
            .O(N__20392),
            .I(N__20385));
    InMux I__2585 (
            .O(N__20391),
            .I(N__20382));
    LocalMux I__2584 (
            .O(N__20388),
            .I(cmd_rdadctmp_9_adj_1103));
    LocalMux I__2583 (
            .O(N__20385),
            .I(cmd_rdadctmp_9_adj_1103));
    LocalMux I__2582 (
            .O(N__20382),
            .I(cmd_rdadctmp_9_adj_1103));
    InMux I__2581 (
            .O(N__20375),
            .I(N__20371));
    CascadeMux I__2580 (
            .O(N__20374),
            .I(N__20367));
    LocalMux I__2579 (
            .O(N__20371),
            .I(N__20364));
    InMux I__2578 (
            .O(N__20370),
            .I(N__20359));
    InMux I__2577 (
            .O(N__20367),
            .I(N__20359));
    Odrv4 I__2576 (
            .O(N__20364),
            .I(cmd_rdadctmp_28));
    LocalMux I__2575 (
            .O(N__20359),
            .I(cmd_rdadctmp_28));
    InMux I__2574 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__2573 (
            .O(N__20351),
            .I(N__20348));
    Span4Mux_v I__2572 (
            .O(N__20348),
            .I(N__20345));
    Span4Mux_h I__2571 (
            .O(N__20345),
            .I(N__20341));
    InMux I__2570 (
            .O(N__20344),
            .I(N__20338));
    Sp12to4 I__2569 (
            .O(N__20341),
            .I(N__20335));
    LocalMux I__2568 (
            .O(N__20338),
            .I(buf_adcdata2_17));
    Odrv12 I__2567 (
            .O(N__20335),
            .I(buf_adcdata2_17));
    InMux I__2566 (
            .O(N__20330),
            .I(N__20327));
    LocalMux I__2565 (
            .O(N__20327),
            .I(N__20323));
    CascadeMux I__2564 (
            .O(N__20326),
            .I(N__20319));
    Span4Mux_v I__2563 (
            .O(N__20323),
            .I(N__20316));
    CascadeMux I__2562 (
            .O(N__20322),
            .I(N__20313));
    InMux I__2561 (
            .O(N__20319),
            .I(N__20310));
    Span4Mux_h I__2560 (
            .O(N__20316),
            .I(N__20307));
    InMux I__2559 (
            .O(N__20313),
            .I(N__20304));
    LocalMux I__2558 (
            .O(N__20310),
            .I(cmd_rdadctmp_13_adj_1099));
    Odrv4 I__2557 (
            .O(N__20307),
            .I(cmd_rdadctmp_13_adj_1099));
    LocalMux I__2556 (
            .O(N__20304),
            .I(cmd_rdadctmp_13_adj_1099));
    CascadeMux I__2555 (
            .O(N__20297),
            .I(N__20293));
    CascadeMux I__2554 (
            .O(N__20296),
            .I(N__20289));
    InMux I__2553 (
            .O(N__20293),
            .I(N__20286));
    InMux I__2552 (
            .O(N__20292),
            .I(N__20281));
    InMux I__2551 (
            .O(N__20289),
            .I(N__20281));
    LocalMux I__2550 (
            .O(N__20286),
            .I(cmd_rdadctmp_14_adj_1098));
    LocalMux I__2549 (
            .O(N__20281),
            .I(cmd_rdadctmp_14_adj_1098));
    InMux I__2548 (
            .O(N__20276),
            .I(N__20273));
    LocalMux I__2547 (
            .O(N__20273),
            .I(N__20270));
    Sp12to4 I__2546 (
            .O(N__20270),
            .I(N__20267));
    Span12Mux_v I__2545 (
            .O(N__20267),
            .I(N__20264));
    Span12Mux_h I__2544 (
            .O(N__20264),
            .I(N__20261));
    Odrv12 I__2543 (
            .O(N__20261),
            .I(buf_data2_14));
    InMux I__2542 (
            .O(N__20258),
            .I(N__20255));
    LocalMux I__2541 (
            .O(N__20255),
            .I(N__20252));
    Odrv12 I__2540 (
            .O(N__20252),
            .I(n4058));
    InMux I__2539 (
            .O(N__20249),
            .I(N__20240));
    InMux I__2538 (
            .O(N__20248),
            .I(N__20240));
    InMux I__2537 (
            .O(N__20247),
            .I(N__20240));
    LocalMux I__2536 (
            .O(N__20240),
            .I(cmd_rdadctmp_27));
    InMux I__2535 (
            .O(N__20237),
            .I(N__20234));
    LocalMux I__2534 (
            .O(N__20234),
            .I(N__20231));
    Span4Mux_h I__2533 (
            .O(N__20231),
            .I(N__20228));
    Span4Mux_h I__2532 (
            .O(N__20228),
            .I(N__20224));
    CascadeMux I__2531 (
            .O(N__20227),
            .I(N__20221));
    Span4Mux_h I__2530 (
            .O(N__20224),
            .I(N__20218));
    InMux I__2529 (
            .O(N__20221),
            .I(N__20215));
    Span4Mux_h I__2528 (
            .O(N__20218),
            .I(N__20212));
    LocalMux I__2527 (
            .O(N__20215),
            .I(buf_adcdata1_19));
    Odrv4 I__2526 (
            .O(N__20212),
            .I(buf_adcdata1_19));
    CascadeMux I__2525 (
            .O(N__20207),
            .I(N__20203));
    CascadeMux I__2524 (
            .O(N__20206),
            .I(N__20199));
    InMux I__2523 (
            .O(N__20203),
            .I(N__20192));
    InMux I__2522 (
            .O(N__20202),
            .I(N__20192));
    InMux I__2521 (
            .O(N__20199),
            .I(N__20192));
    LocalMux I__2520 (
            .O(N__20192),
            .I(cmd_rdadctmp_25));
    InMux I__2519 (
            .O(N__20189),
            .I(N__20186));
    LocalMux I__2518 (
            .O(N__20186),
            .I(N__20183));
    Span12Mux_v I__2517 (
            .O(N__20183),
            .I(N__20179));
    CascadeMux I__2516 (
            .O(N__20182),
            .I(N__20176));
    Span12Mux_h I__2515 (
            .O(N__20179),
            .I(N__20173));
    InMux I__2514 (
            .O(N__20176),
            .I(N__20170));
    Span12Mux_v I__2513 (
            .O(N__20173),
            .I(N__20167));
    LocalMux I__2512 (
            .O(N__20170),
            .I(buf_adcdata1_20));
    Odrv12 I__2511 (
            .O(N__20167),
            .I(buf_adcdata1_20));
    CascadeMux I__2510 (
            .O(N__20162),
            .I(n84_cascade_));
    CascadeMux I__2509 (
            .O(N__20159),
            .I(n15593_cascade_));
    CascadeMux I__2508 (
            .O(N__20156),
            .I(n8045_cascade_));
    InMux I__2507 (
            .O(N__20153),
            .I(N__20150));
    LocalMux I__2506 (
            .O(N__20150),
            .I(n15573));
    InMux I__2505 (
            .O(N__20147),
            .I(N__20144));
    LocalMux I__2504 (
            .O(N__20144),
            .I(N__20141));
    Span4Mux_v I__2503 (
            .O(N__20141),
            .I(N__20138));
    Odrv4 I__2502 (
            .O(N__20138),
            .I(comm_buf_4_5));
    InMux I__2501 (
            .O(N__20135),
            .I(N__20132));
    LocalMux I__2500 (
            .O(N__20132),
            .I(N__20129));
    Odrv12 I__2499 (
            .O(N__20129),
            .I(comm_buf_4_6));
    InMux I__2498 (
            .O(N__20126),
            .I(N__20123));
    LocalMux I__2497 (
            .O(N__20123),
            .I(N__20120));
    Span4Mux_h I__2496 (
            .O(N__20120),
            .I(N__20117));
    Span4Mux_v I__2495 (
            .O(N__20117),
            .I(N__20114));
    Span4Mux_h I__2494 (
            .O(N__20114),
            .I(N__20111));
    Span4Mux_h I__2493 (
            .O(N__20111),
            .I(N__20108));
    Odrv4 I__2492 (
            .O(N__20108),
            .I(buf_data2_15));
    CascadeMux I__2491 (
            .O(N__20105),
            .I(n4057_cascade_));
    SRMux I__2490 (
            .O(N__20102),
            .I(N__20099));
    LocalMux I__2489 (
            .O(N__20099),
            .I(N__20096));
    Span4Mux_v I__2488 (
            .O(N__20096),
            .I(N__20092));
    SRMux I__2487 (
            .O(N__20095),
            .I(N__20089));
    Span4Mux_h I__2486 (
            .O(N__20092),
            .I(N__20083));
    LocalMux I__2485 (
            .O(N__20089),
            .I(N__20083));
    SRMux I__2484 (
            .O(N__20088),
            .I(N__20080));
    Span4Mux_h I__2483 (
            .O(N__20083),
            .I(N__20077));
    LocalMux I__2482 (
            .O(N__20080),
            .I(N__20074));
    Odrv4 I__2481 (
            .O(N__20077),
            .I(n10604));
    Odrv12 I__2480 (
            .O(N__20074),
            .I(n10604));
    InMux I__2479 (
            .O(N__20069),
            .I(N__20066));
    LocalMux I__2478 (
            .O(N__20066),
            .I(N__20063));
    Span4Mux_v I__2477 (
            .O(N__20063),
            .I(N__20060));
    Span4Mux_h I__2476 (
            .O(N__20060),
            .I(N__20057));
    Span4Mux_h I__2475 (
            .O(N__20057),
            .I(N__20053));
    InMux I__2474 (
            .O(N__20056),
            .I(N__20050));
    Span4Mux_h I__2473 (
            .O(N__20053),
            .I(N__20047));
    LocalMux I__2472 (
            .O(N__20050),
            .I(buf_adcdata1_17));
    Odrv4 I__2471 (
            .O(N__20047),
            .I(buf_adcdata1_17));
    InMux I__2470 (
            .O(N__20042),
            .I(N__20038));
    CascadeMux I__2469 (
            .O(N__20041),
            .I(N__20035));
    LocalMux I__2468 (
            .O(N__20038),
            .I(N__20032));
    InMux I__2467 (
            .O(N__20035),
            .I(N__20029));
    Span12Mux_h I__2466 (
            .O(N__20032),
            .I(N__20026));
    LocalMux I__2465 (
            .O(N__20029),
            .I(buf_adcdata1_18));
    Odrv12 I__2464 (
            .O(N__20026),
            .I(buf_adcdata1_18));
    CascadeMux I__2463 (
            .O(N__20021),
            .I(N__20016));
    InMux I__2462 (
            .O(N__20020),
            .I(N__20009));
    InMux I__2461 (
            .O(N__20019),
            .I(N__20009));
    InMux I__2460 (
            .O(N__20016),
            .I(N__20009));
    LocalMux I__2459 (
            .O(N__20009),
            .I(cmd_rdadctmp_26));
    CascadeMux I__2458 (
            .O(N__20006),
            .I(n16407_cascade_));
    InMux I__2457 (
            .O(N__20003),
            .I(N__20000));
    LocalMux I__2456 (
            .O(N__20000),
            .I(N__19997));
    Span4Mux_v I__2455 (
            .O(N__19997),
            .I(N__19994));
    Odrv4 I__2454 (
            .O(N__19994),
            .I(comm_buf_5_1));
    CascadeMux I__2453 (
            .O(N__19991),
            .I(N__19988));
    InMux I__2452 (
            .O(N__19988),
            .I(N__19985));
    LocalMux I__2451 (
            .O(N__19985),
            .I(N__19982));
    Span4Mux_v I__2450 (
            .O(N__19982),
            .I(N__19979));
    Odrv4 I__2449 (
            .O(N__19979),
            .I(comm_buf_4_1));
    InMux I__2448 (
            .O(N__19976),
            .I(N__19973));
    LocalMux I__2447 (
            .O(N__19973),
            .I(n16515));
    InMux I__2446 (
            .O(N__19970),
            .I(N__19967));
    LocalMux I__2445 (
            .O(N__19967),
            .I(n16512));
    InMux I__2444 (
            .O(N__19964),
            .I(N__19961));
    LocalMux I__2443 (
            .O(N__19961),
            .I(n7_adj_1240));
    CascadeMux I__2442 (
            .O(N__19958),
            .I(n16425_cascade_));
    InMux I__2441 (
            .O(N__19955),
            .I(N__19952));
    LocalMux I__2440 (
            .O(N__19952),
            .I(N__19949));
    Span4Mux_v I__2439 (
            .O(N__19949),
            .I(N__19946));
    Span4Mux_v I__2438 (
            .O(N__19946),
            .I(N__19943));
    Span4Mux_h I__2437 (
            .O(N__19943),
            .I(N__19940));
    Sp12to4 I__2436 (
            .O(N__19940),
            .I(N__19937));
    Odrv12 I__2435 (
            .O(N__19937),
            .I(buf_data2_12));
    CascadeMux I__2434 (
            .O(N__19934),
            .I(n4060_cascade_));
    CascadeMux I__2433 (
            .O(N__19931),
            .I(n16413_cascade_));
    InMux I__2432 (
            .O(N__19928),
            .I(N__19925));
    LocalMux I__2431 (
            .O(N__19925),
            .I(N__19922));
    Odrv4 I__2430 (
            .O(N__19922),
            .I(comm_buf_5_6));
    CascadeMux I__2429 (
            .O(N__19919),
            .I(n16518_cascade_));
    InMux I__2428 (
            .O(N__19916),
            .I(N__19913));
    LocalMux I__2427 (
            .O(N__19913),
            .I(n13493));
    CascadeMux I__2426 (
            .O(N__19910),
            .I(n16521_cascade_));
    InMux I__2425 (
            .O(N__19907),
            .I(N__19904));
    LocalMux I__2424 (
            .O(N__19904),
            .I(N__19901));
    Span4Mux_v I__2423 (
            .O(N__19901),
            .I(N__19898));
    Odrv4 I__2422 (
            .O(N__19898),
            .I(comm_buf_2_6));
    CascadeMux I__2421 (
            .O(N__19895),
            .I(N__19892));
    InMux I__2420 (
            .O(N__19892),
            .I(N__19889));
    LocalMux I__2419 (
            .O(N__19889),
            .I(comm_buf_3_6));
    InMux I__2418 (
            .O(N__19886),
            .I(N__19883));
    LocalMux I__2417 (
            .O(N__19883),
            .I(n16410));
    InMux I__2416 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__2415 (
            .O(N__19877),
            .I(n16491));
    InMux I__2414 (
            .O(N__19874),
            .I(N__19871));
    LocalMux I__2413 (
            .O(N__19871),
            .I(N__19868));
    Span4Mux_h I__2412 (
            .O(N__19868),
            .I(N__19865));
    Odrv4 I__2411 (
            .O(N__19865),
            .I(comm_buf_2_1));
    CascadeMux I__2410 (
            .O(N__19862),
            .I(N__19859));
    InMux I__2409 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__2408 (
            .O(N__19856),
            .I(N__19853));
    Odrv12 I__2407 (
            .O(N__19853),
            .I(comm_buf_3_1));
    CascadeMux I__2406 (
            .O(N__19850),
            .I(n16404_cascade_));
    InMux I__2405 (
            .O(N__19847),
            .I(N__19843));
    CascadeMux I__2404 (
            .O(N__19846),
            .I(N__19840));
    LocalMux I__2403 (
            .O(N__19843),
            .I(N__19837));
    InMux I__2402 (
            .O(N__19840),
            .I(N__19834));
    Odrv4 I__2401 (
            .O(N__19837),
            .I(cmd_rdadctmp_1_adj_1148));
    LocalMux I__2400 (
            .O(N__19834),
            .I(cmd_rdadctmp_1_adj_1148));
    CascadeMux I__2399 (
            .O(N__19829),
            .I(N__19826));
    InMux I__2398 (
            .O(N__19826),
            .I(N__19823));
    LocalMux I__2397 (
            .O(N__19823),
            .I(N__19820));
    Span4Mux_v I__2396 (
            .O(N__19820),
            .I(N__19817));
    Sp12to4 I__2395 (
            .O(N__19817),
            .I(N__19814));
    Span12Mux_h I__2394 (
            .O(N__19814),
            .I(N__19811));
    Span12Mux_h I__2393 (
            .O(N__19811),
            .I(N__19808));
    Odrv12 I__2392 (
            .O(N__19808),
            .I(M_MISO4));
    InMux I__2391 (
            .O(N__19805),
            .I(N__19801));
    InMux I__2390 (
            .O(N__19804),
            .I(N__19798));
    LocalMux I__2389 (
            .O(N__19801),
            .I(cmd_rdadctmp_0_adj_1149));
    LocalMux I__2388 (
            .O(N__19798),
            .I(cmd_rdadctmp_0_adj_1149));
    CascadeMux I__2387 (
            .O(N__19793),
            .I(N__19790));
    InMux I__2386 (
            .O(N__19790),
            .I(N__19787));
    LocalMux I__2385 (
            .O(N__19787),
            .I(N__19784));
    Span4Mux_h I__2384 (
            .O(N__19784),
            .I(N__19779));
    InMux I__2383 (
            .O(N__19783),
            .I(N__19776));
    InMux I__2382 (
            .O(N__19782),
            .I(N__19773));
    Odrv4 I__2381 (
            .O(N__19779),
            .I(cmd_rdadctmp_15));
    LocalMux I__2380 (
            .O(N__19776),
            .I(cmd_rdadctmp_15));
    LocalMux I__2379 (
            .O(N__19773),
            .I(cmd_rdadctmp_15));
    IoInMux I__2378 (
            .O(N__19766),
            .I(N__19763));
    LocalMux I__2377 (
            .O(N__19763),
            .I(N__19760));
    IoSpan4Mux I__2376 (
            .O(N__19760),
            .I(N__19757));
    Span4Mux_s1_v I__2375 (
            .O(N__19757),
            .I(N__19754));
    Span4Mux_v I__2374 (
            .O(N__19754),
            .I(N__19751));
    Odrv4 I__2373 (
            .O(N__19751),
            .I(M_START));
    InMux I__2372 (
            .O(N__19748),
            .I(N__19745));
    LocalMux I__2371 (
            .O(N__19745),
            .I(N__19742));
    Odrv4 I__2370 (
            .O(N__19742),
            .I(comm_buf_3_0));
    InMux I__2369 (
            .O(N__19739),
            .I(N__19736));
    LocalMux I__2368 (
            .O(N__19736),
            .I(N__19733));
    Span4Mux_v I__2367 (
            .O(N__19733),
            .I(N__19730));
    Odrv4 I__2366 (
            .O(N__19730),
            .I(comm_buf_2_0));
    CascadeMux I__2365 (
            .O(N__19727),
            .I(N__19723));
    CascadeMux I__2364 (
            .O(N__19726),
            .I(N__19719));
    InMux I__2363 (
            .O(N__19723),
            .I(N__19712));
    InMux I__2362 (
            .O(N__19722),
            .I(N__19712));
    InMux I__2361 (
            .O(N__19719),
            .I(N__19712));
    LocalMux I__2360 (
            .O(N__19712),
            .I(cmd_rdadctmp_18_adj_1131));
    CascadeMux I__2359 (
            .O(N__19709),
            .I(N__19705));
    InMux I__2358 (
            .O(N__19708),
            .I(N__19702));
    InMux I__2357 (
            .O(N__19705),
            .I(N__19699));
    LocalMux I__2356 (
            .O(N__19702),
            .I(N__19696));
    LocalMux I__2355 (
            .O(N__19699),
            .I(N__19692));
    Span12Mux_v I__2354 (
            .O(N__19696),
            .I(N__19689));
    InMux I__2353 (
            .O(N__19695),
            .I(N__19686));
    Span4Mux_v I__2352 (
            .O(N__19692),
            .I(N__19683));
    Span12Mux_h I__2351 (
            .O(N__19689),
            .I(N__19680));
    LocalMux I__2350 (
            .O(N__19686),
            .I(buf_adcdata4_10));
    Odrv4 I__2349 (
            .O(N__19683),
            .I(buf_adcdata4_10));
    Odrv12 I__2348 (
            .O(N__19680),
            .I(buf_adcdata4_10));
    CascadeMux I__2347 (
            .O(N__19673),
            .I(\ADC_VAC1.n15263_cascade_ ));
    InMux I__2346 (
            .O(N__19670),
            .I(N__19667));
    LocalMux I__2345 (
            .O(N__19667),
            .I(\ADC_VAC1.n15553 ));
    CEMux I__2344 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__2343 (
            .O(N__19661),
            .I(\ADC_VAC1.n15264 ));
    CascadeMux I__2342 (
            .O(N__19658),
            .I(N__19654));
    InMux I__2341 (
            .O(N__19657),
            .I(N__19649));
    InMux I__2340 (
            .O(N__19654),
            .I(N__19649));
    LocalMux I__2339 (
            .O(N__19649),
            .I(N__19644));
    CascadeMux I__2338 (
            .O(N__19648),
            .I(N__19641));
    CascadeMux I__2337 (
            .O(N__19647),
            .I(N__19637));
    Span4Mux_v I__2336 (
            .O(N__19644),
            .I(N__19634));
    InMux I__2335 (
            .O(N__19641),
            .I(N__19631));
    InMux I__2334 (
            .O(N__19640),
            .I(N__19628));
    InMux I__2333 (
            .O(N__19637),
            .I(N__19625));
    Span4Mux_h I__2332 (
            .O(N__19634),
            .I(N__19622));
    LocalMux I__2331 (
            .O(N__19631),
            .I(N__19615));
    LocalMux I__2330 (
            .O(N__19628),
            .I(N__19615));
    LocalMux I__2329 (
            .O(N__19625),
            .I(N__19615));
    Sp12to4 I__2328 (
            .O(N__19622),
            .I(N__19610));
    Span12Mux_v I__2327 (
            .O(N__19615),
            .I(N__19610));
    Odrv12 I__2326 (
            .O(N__19610),
            .I(M_DRDY1));
    CascadeMux I__2325 (
            .O(N__19607),
            .I(\ADC_VAC1.n17_cascade_ ));
    CEMux I__2324 (
            .O(N__19604),
            .I(N__19601));
    LocalMux I__2323 (
            .O(N__19601),
            .I(N__19598));
    Odrv4 I__2322 (
            .O(N__19598),
            .I(\ADC_VAC1.n12 ));
    CascadeMux I__2321 (
            .O(N__19595),
            .I(N__19592));
    InMux I__2320 (
            .O(N__19592),
            .I(N__19587));
    InMux I__2319 (
            .O(N__19591),
            .I(N__19584));
    CascadeMux I__2318 (
            .O(N__19590),
            .I(N__19581));
    LocalMux I__2317 (
            .O(N__19587),
            .I(N__19578));
    LocalMux I__2316 (
            .O(N__19584),
            .I(N__19575));
    InMux I__2315 (
            .O(N__19581),
            .I(N__19572));
    Odrv4 I__2314 (
            .O(N__19578),
            .I(cmd_rdadctmp_13));
    Odrv4 I__2313 (
            .O(N__19575),
            .I(cmd_rdadctmp_13));
    LocalMux I__2312 (
            .O(N__19572),
            .I(cmd_rdadctmp_13));
    CascadeMux I__2311 (
            .O(N__19565),
            .I(N__19561));
    InMux I__2310 (
            .O(N__19564),
            .I(N__19558));
    InMux I__2309 (
            .O(N__19561),
            .I(N__19555));
    LocalMux I__2308 (
            .O(N__19558),
            .I(N__19552));
    LocalMux I__2307 (
            .O(N__19555),
            .I(N__19548));
    Span4Mux_v I__2306 (
            .O(N__19552),
            .I(N__19545));
    InMux I__2305 (
            .O(N__19551),
            .I(N__19542));
    Span4Mux_h I__2304 (
            .O(N__19548),
            .I(N__19539));
    Span4Mux_h I__2303 (
            .O(N__19545),
            .I(N__19536));
    LocalMux I__2302 (
            .O(N__19542),
            .I(buf_adcdata3_5));
    Odrv4 I__2301 (
            .O(N__19539),
            .I(buf_adcdata3_5));
    Odrv4 I__2300 (
            .O(N__19536),
            .I(buf_adcdata3_5));
    InMux I__2299 (
            .O(N__19529),
            .I(N__19525));
    CascadeMux I__2298 (
            .O(N__19528),
            .I(N__19522));
    LocalMux I__2297 (
            .O(N__19525),
            .I(N__19519));
    InMux I__2296 (
            .O(N__19522),
            .I(N__19516));
    Span4Mux_h I__2295 (
            .O(N__19519),
            .I(N__19512));
    LocalMux I__2294 (
            .O(N__19516),
            .I(N__19509));
    InMux I__2293 (
            .O(N__19515),
            .I(N__19506));
    Span4Mux_v I__2292 (
            .O(N__19512),
            .I(N__19503));
    Span4Mux_v I__2291 (
            .O(N__19509),
            .I(N__19500));
    LocalMux I__2290 (
            .O(N__19506),
            .I(buf_adcdata3_6));
    Odrv4 I__2289 (
            .O(N__19503),
            .I(buf_adcdata3_6));
    Odrv4 I__2288 (
            .O(N__19500),
            .I(buf_adcdata3_6));
    CascadeMux I__2287 (
            .O(N__19493),
            .I(N__19489));
    CascadeMux I__2286 (
            .O(N__19492),
            .I(N__19485));
    InMux I__2285 (
            .O(N__19489),
            .I(N__19480));
    InMux I__2284 (
            .O(N__19488),
            .I(N__19480));
    InMux I__2283 (
            .O(N__19485),
            .I(N__19477));
    LocalMux I__2282 (
            .O(N__19480),
            .I(cmd_rdadctmp_12));
    LocalMux I__2281 (
            .O(N__19477),
            .I(cmd_rdadctmp_12));
    CascadeMux I__2280 (
            .O(N__19472),
            .I(N__19467));
    CascadeMux I__2279 (
            .O(N__19471),
            .I(N__19464));
    CascadeMux I__2278 (
            .O(N__19470),
            .I(N__19461));
    InMux I__2277 (
            .O(N__19467),
            .I(N__19456));
    InMux I__2276 (
            .O(N__19464),
            .I(N__19456));
    InMux I__2275 (
            .O(N__19461),
            .I(N__19453));
    LocalMux I__2274 (
            .O(N__19456),
            .I(cmd_rdadctmp_10_adj_1102));
    LocalMux I__2273 (
            .O(N__19453),
            .I(cmd_rdadctmp_10_adj_1102));
    InMux I__2272 (
            .O(N__19448),
            .I(N__19442));
    InMux I__2271 (
            .O(N__19447),
            .I(N__19442));
    LocalMux I__2270 (
            .O(N__19442),
            .I(N__19438));
    CascadeMux I__2269 (
            .O(N__19441),
            .I(N__19435));
    Span4Mux_h I__2268 (
            .O(N__19438),
            .I(N__19432));
    InMux I__2267 (
            .O(N__19435),
            .I(N__19429));
    Odrv4 I__2266 (
            .O(N__19432),
            .I(cmd_rdadctmp_16_adj_1133));
    LocalMux I__2265 (
            .O(N__19429),
            .I(cmd_rdadctmp_16_adj_1133));
    CascadeMux I__2264 (
            .O(N__19424),
            .I(N__19419));
    InMux I__2263 (
            .O(N__19423),
            .I(N__19412));
    InMux I__2262 (
            .O(N__19422),
            .I(N__19412));
    InMux I__2261 (
            .O(N__19419),
            .I(N__19412));
    LocalMux I__2260 (
            .O(N__19412),
            .I(cmd_rdadctmp_17_adj_1132));
    InMux I__2259 (
            .O(N__19409),
            .I(N__19406));
    LocalMux I__2258 (
            .O(N__19406),
            .I(comm_buf_4_3));
    InMux I__2257 (
            .O(N__19403),
            .I(N__19400));
    LocalMux I__2256 (
            .O(N__19400),
            .I(N__19397));
    Span4Mux_v I__2255 (
            .O(N__19397),
            .I(N__19394));
    Odrv4 I__2254 (
            .O(N__19394),
            .I(comm_buf_5_3));
    CascadeMux I__2253 (
            .O(N__19391),
            .I(n16440_cascade_));
    CascadeMux I__2252 (
            .O(N__19388),
            .I(N__19385));
    InMux I__2251 (
            .O(N__19385),
            .I(N__19382));
    LocalMux I__2250 (
            .O(N__19382),
            .I(n15423));
    InMux I__2249 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__2248 (
            .O(N__19376),
            .I(n15397));
    CascadeMux I__2247 (
            .O(N__19373),
            .I(n16392_cascade_));
    InMux I__2246 (
            .O(N__19370),
            .I(N__19367));
    LocalMux I__2245 (
            .O(N__19367),
            .I(n16443));
    CascadeMux I__2244 (
            .O(N__19364),
            .I(n16395_cascade_));
    IoInMux I__2243 (
            .O(N__19361),
            .I(N__19358));
    LocalMux I__2242 (
            .O(N__19358),
            .I(N__19355));
    IoSpan4Mux I__2241 (
            .O(N__19355),
            .I(N__19352));
    Span4Mux_s2_h I__2240 (
            .O(N__19352),
            .I(N__19349));
    Sp12to4 I__2239 (
            .O(N__19349),
            .I(N__19345));
    CascadeMux I__2238 (
            .O(N__19348),
            .I(N__19342));
    Span12Mux_v I__2237 (
            .O(N__19345),
            .I(N__19339));
    InMux I__2236 (
            .O(N__19342),
            .I(N__19336));
    Odrv12 I__2235 (
            .O(N__19339),
            .I(M_SCLK2));
    LocalMux I__2234 (
            .O(N__19336),
            .I(M_SCLK2));
    CascadeMux I__2233 (
            .O(N__19331),
            .I(n15388_cascade_));
    CascadeMux I__2232 (
            .O(N__19328),
            .I(n16389_cascade_));
    InMux I__2231 (
            .O(N__19325),
            .I(N__19322));
    LocalMux I__2230 (
            .O(N__19322),
            .I(comm_buf_4_2));
    InMux I__2229 (
            .O(N__19319),
            .I(N__19316));
    LocalMux I__2228 (
            .O(N__19316),
            .I(N__19313));
    Odrv12 I__2227 (
            .O(N__19313),
            .I(comm_buf_5_2));
    InMux I__2226 (
            .O(N__19310),
            .I(N__19307));
    LocalMux I__2225 (
            .O(N__19307),
            .I(n15448));
    CascadeMux I__2224 (
            .O(N__19304),
            .I(n15447_cascade_));
    InMux I__2223 (
            .O(N__19301),
            .I(N__19298));
    LocalMux I__2222 (
            .O(N__19298),
            .I(n16386));
    InMux I__2221 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__2220 (
            .O(N__19292),
            .I(N__19289));
    Span4Mux_h I__2219 (
            .O(N__19289),
            .I(N__19286));
    Span4Mux_h I__2218 (
            .O(N__19286),
            .I(N__19282));
    CascadeMux I__2217 (
            .O(N__19285),
            .I(N__19279));
    Span4Mux_h I__2216 (
            .O(N__19282),
            .I(N__19275));
    InMux I__2215 (
            .O(N__19279),
            .I(N__19272));
    InMux I__2214 (
            .O(N__19278),
            .I(N__19269));
    Span4Mux_h I__2213 (
            .O(N__19275),
            .I(N__19264));
    LocalMux I__2212 (
            .O(N__19272),
            .I(N__19264));
    LocalMux I__2211 (
            .O(N__19269),
            .I(buf_adcdata4_18));
    Odrv4 I__2210 (
            .O(N__19264),
            .I(buf_adcdata4_18));
    InMux I__2209 (
            .O(N__19259),
            .I(N__19256));
    LocalMux I__2208 (
            .O(N__19256),
            .I(N__19253));
    Span4Mux_v I__2207 (
            .O(N__19253),
            .I(N__19250));
    Odrv4 I__2206 (
            .O(N__19250),
            .I(comm_buf_2_3));
    InMux I__2205 (
            .O(N__19247),
            .I(N__19244));
    LocalMux I__2204 (
            .O(N__19244),
            .I(N__19241));
    Span4Mux_h I__2203 (
            .O(N__19241),
            .I(N__19238));
    Span4Mux_v I__2202 (
            .O(N__19238),
            .I(N__19235));
    Span4Mux_h I__2201 (
            .O(N__19235),
            .I(N__19232));
    Span4Mux_h I__2200 (
            .O(N__19232),
            .I(N__19229));
    Odrv4 I__2199 (
            .O(N__19229),
            .I(buf_data2_17));
    CascadeMux I__2198 (
            .O(N__19226),
            .I(n4107_cascade_));
    InMux I__2197 (
            .O(N__19223),
            .I(N__19220));
    LocalMux I__2196 (
            .O(N__19220),
            .I(N__19217));
    Span4Mux_h I__2195 (
            .O(N__19217),
            .I(N__19214));
    Span4Mux_h I__2194 (
            .O(N__19214),
            .I(N__19211));
    Span4Mux_h I__2193 (
            .O(N__19211),
            .I(N__19208));
    Span4Mux_h I__2192 (
            .O(N__19208),
            .I(N__19205));
    Odrv4 I__2191 (
            .O(N__19205),
            .I(buf_data2_18));
    CEMux I__2190 (
            .O(N__19202),
            .I(N__19198));
    CEMux I__2189 (
            .O(N__19201),
            .I(N__19195));
    LocalMux I__2188 (
            .O(N__19198),
            .I(N__19192));
    LocalMux I__2187 (
            .O(N__19195),
            .I(N__19189));
    Span4Mux_v I__2186 (
            .O(N__19192),
            .I(N__19186));
    Span4Mux_v I__2185 (
            .O(N__19189),
            .I(N__19183));
    Odrv4 I__2184 (
            .O(N__19186),
            .I(n8787));
    Odrv4 I__2183 (
            .O(N__19183),
            .I(n8787));
    SRMux I__2182 (
            .O(N__19178),
            .I(N__19175));
    LocalMux I__2181 (
            .O(N__19175),
            .I(N__19171));
    SRMux I__2180 (
            .O(N__19174),
            .I(N__19168));
    Span4Mux_v I__2179 (
            .O(N__19171),
            .I(N__19165));
    LocalMux I__2178 (
            .O(N__19168),
            .I(N__19162));
    Span4Mux_h I__2177 (
            .O(N__19165),
            .I(N__19157));
    Span4Mux_v I__2176 (
            .O(N__19162),
            .I(N__19157));
    Odrv4 I__2175 (
            .O(N__19157),
            .I(n10599));
    CascadeMux I__2174 (
            .O(N__19154),
            .I(N__19151));
    InMux I__2173 (
            .O(N__19151),
            .I(N__19148));
    LocalMux I__2172 (
            .O(N__19148),
            .I(comm_buf_2_2));
    InMux I__2171 (
            .O(N__19145),
            .I(\ADC_VAC1.n13987 ));
    InMux I__2170 (
            .O(N__19142),
            .I(N__19138));
    InMux I__2169 (
            .O(N__19141),
            .I(N__19135));
    LocalMux I__2168 (
            .O(N__19138),
            .I(\ADC_VAC1.bit_cnt_7 ));
    LocalMux I__2167 (
            .O(N__19135),
            .I(\ADC_VAC1.bit_cnt_7 ));
    CEMux I__2166 (
            .O(N__19130),
            .I(N__19127));
    LocalMux I__2165 (
            .O(N__19127),
            .I(N__19124));
    Odrv4 I__2164 (
            .O(N__19124),
            .I(\ADC_VAC1.n9312 ));
    SRMux I__2163 (
            .O(N__19121),
            .I(N__19118));
    LocalMux I__2162 (
            .O(N__19118),
            .I(\ADC_VAC1.n10667 ));
    CascadeMux I__2161 (
            .O(N__19115),
            .I(n16470_cascade_));
    InMux I__2160 (
            .O(N__19112),
            .I(N__19109));
    LocalMux I__2159 (
            .O(N__19109),
            .I(N__19106));
    Span4Mux_h I__2158 (
            .O(N__19106),
            .I(N__19103));
    Odrv4 I__2157 (
            .O(N__19103),
            .I(comm_buf_5_5));
    InMux I__2156 (
            .O(N__19100),
            .I(N__19097));
    LocalMux I__2155 (
            .O(N__19097),
            .I(N__19094));
    Span4Mux_h I__2154 (
            .O(N__19094),
            .I(N__19091));
    Odrv4 I__2153 (
            .O(N__19091),
            .I(comm_buf_2_5));
    CascadeMux I__2152 (
            .O(N__19088),
            .I(n16416_cascade_));
    InMux I__2151 (
            .O(N__19085),
            .I(N__19082));
    LocalMux I__2150 (
            .O(N__19082),
            .I(n16473));
    CascadeMux I__2149 (
            .O(N__19079),
            .I(n16419_cascade_));
    CascadeMux I__2148 (
            .O(N__19076),
            .I(n7_adj_1238_cascade_));
    InMux I__2147 (
            .O(N__19073),
            .I(N__19070));
    LocalMux I__2146 (
            .O(N__19070),
            .I(N__19067));
    Span4Mux_v I__2145 (
            .O(N__19067),
            .I(N__19064));
    Sp12to4 I__2144 (
            .O(N__19064),
            .I(N__19061));
    Span12Mux_h I__2143 (
            .O(N__19061),
            .I(N__19058));
    Odrv12 I__2142 (
            .O(N__19058),
            .I(buf_data2_21));
    CascadeMux I__2141 (
            .O(N__19055),
            .I(n4103_cascade_));
    CascadeMux I__2140 (
            .O(N__19052),
            .I(N__19049));
    InMux I__2139 (
            .O(N__19049),
            .I(N__19046));
    LocalMux I__2138 (
            .O(N__19046),
            .I(comm_buf_3_5));
    CascadeMux I__2137 (
            .O(N__19043),
            .I(\ADC_VAC1.n15360_cascade_ ));
    InMux I__2136 (
            .O(N__19040),
            .I(N__19036));
    InMux I__2135 (
            .O(N__19039),
            .I(N__19033));
    LocalMux I__2134 (
            .O(N__19036),
            .I(\ADC_VAC1.bit_cnt_0 ));
    LocalMux I__2133 (
            .O(N__19033),
            .I(\ADC_VAC1.bit_cnt_0 ));
    InMux I__2132 (
            .O(N__19028),
            .I(bfn_6_16_0_));
    CascadeMux I__2131 (
            .O(N__19025),
            .I(N__19021));
    InMux I__2130 (
            .O(N__19024),
            .I(N__19018));
    InMux I__2129 (
            .O(N__19021),
            .I(N__19015));
    LocalMux I__2128 (
            .O(N__19018),
            .I(\ADC_VAC1.bit_cnt_1 ));
    LocalMux I__2127 (
            .O(N__19015),
            .I(\ADC_VAC1.bit_cnt_1 ));
    InMux I__2126 (
            .O(N__19010),
            .I(\ADC_VAC1.n13981 ));
    InMux I__2125 (
            .O(N__19007),
            .I(N__19003));
    InMux I__2124 (
            .O(N__19006),
            .I(N__19000));
    LocalMux I__2123 (
            .O(N__19003),
            .I(\ADC_VAC1.bit_cnt_2 ));
    LocalMux I__2122 (
            .O(N__19000),
            .I(\ADC_VAC1.bit_cnt_2 ));
    InMux I__2121 (
            .O(N__18995),
            .I(\ADC_VAC1.n13982 ));
    InMux I__2120 (
            .O(N__18992),
            .I(N__18988));
    InMux I__2119 (
            .O(N__18991),
            .I(N__18985));
    LocalMux I__2118 (
            .O(N__18988),
            .I(\ADC_VAC1.bit_cnt_3 ));
    LocalMux I__2117 (
            .O(N__18985),
            .I(\ADC_VAC1.bit_cnt_3 ));
    InMux I__2116 (
            .O(N__18980),
            .I(\ADC_VAC1.n13983 ));
    InMux I__2115 (
            .O(N__18977),
            .I(N__18973));
    InMux I__2114 (
            .O(N__18976),
            .I(N__18970));
    LocalMux I__2113 (
            .O(N__18973),
            .I(\ADC_VAC1.bit_cnt_4 ));
    LocalMux I__2112 (
            .O(N__18970),
            .I(\ADC_VAC1.bit_cnt_4 ));
    InMux I__2111 (
            .O(N__18965),
            .I(\ADC_VAC1.n13984 ));
    InMux I__2110 (
            .O(N__18962),
            .I(N__18958));
    InMux I__2109 (
            .O(N__18961),
            .I(N__18955));
    LocalMux I__2108 (
            .O(N__18958),
            .I(N__18952));
    LocalMux I__2107 (
            .O(N__18955),
            .I(\ADC_VAC1.bit_cnt_5 ));
    Odrv4 I__2106 (
            .O(N__18952),
            .I(\ADC_VAC1.bit_cnt_5 ));
    InMux I__2105 (
            .O(N__18947),
            .I(\ADC_VAC1.n13985 ));
    InMux I__2104 (
            .O(N__18944),
            .I(N__18940));
    InMux I__2103 (
            .O(N__18943),
            .I(N__18937));
    LocalMux I__2102 (
            .O(N__18940),
            .I(\ADC_VAC1.bit_cnt_6 ));
    LocalMux I__2101 (
            .O(N__18937),
            .I(\ADC_VAC1.bit_cnt_6 ));
    InMux I__2100 (
            .O(N__18932),
            .I(\ADC_VAC1.n13986 ));
    InMux I__2099 (
            .O(N__18929),
            .I(N__18926));
    LocalMux I__2098 (
            .O(N__18926),
            .I(n15168));
    CascadeMux I__2097 (
            .O(N__18923),
            .I(n15168_cascade_));
    IoInMux I__2096 (
            .O(N__18920),
            .I(N__18917));
    LocalMux I__2095 (
            .O(N__18917),
            .I(N__18914));
    IoSpan4Mux I__2094 (
            .O(N__18914),
            .I(N__18911));
    Span4Mux_s3_h I__2093 (
            .O(N__18911),
            .I(N__18908));
    Span4Mux_h I__2092 (
            .O(N__18908),
            .I(N__18904));
    InMux I__2091 (
            .O(N__18907),
            .I(N__18901));
    Odrv4 I__2090 (
            .O(N__18904),
            .I(M_CS1));
    LocalMux I__2089 (
            .O(N__18901),
            .I(M_CS1));
    InMux I__2088 (
            .O(N__18896),
            .I(N__18893));
    LocalMux I__2087 (
            .O(N__18893),
            .I(n14_adj_1039));
    IoInMux I__2086 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__2085 (
            .O(N__18887),
            .I(N__18884));
    IoSpan4Mux I__2084 (
            .O(N__18884),
            .I(N__18881));
    Span4Mux_s3_h I__2083 (
            .O(N__18881),
            .I(N__18877));
    CascadeMux I__2082 (
            .O(N__18880),
            .I(N__18874));
    Span4Mux_h I__2081 (
            .O(N__18877),
            .I(N__18871));
    InMux I__2080 (
            .O(N__18874),
            .I(N__18868));
    Odrv4 I__2079 (
            .O(N__18871),
            .I(M_SCLK1));
    LocalMux I__2078 (
            .O(N__18868),
            .I(M_SCLK1));
    CascadeMux I__2077 (
            .O(N__18863),
            .I(\ADC_VAC1.n9312_cascade_ ));
    CascadeMux I__2076 (
            .O(N__18860),
            .I(\ADC_VAC1.n15338_cascade_ ));
    InMux I__2075 (
            .O(N__18857),
            .I(N__18853));
    InMux I__2074 (
            .O(N__18856),
            .I(N__18850));
    LocalMux I__2073 (
            .O(N__18853),
            .I(cmd_rdadctmp_2));
    LocalMux I__2072 (
            .O(N__18850),
            .I(cmd_rdadctmp_2));
    InMux I__2071 (
            .O(N__18845),
            .I(N__18839));
    InMux I__2070 (
            .O(N__18844),
            .I(N__18839));
    LocalMux I__2069 (
            .O(N__18839),
            .I(cmd_rdadctmp_7));
    CascadeMux I__2068 (
            .O(N__18836),
            .I(N__18833));
    InMux I__2067 (
            .O(N__18833),
            .I(N__18827));
    InMux I__2066 (
            .O(N__18832),
            .I(N__18827));
    LocalMux I__2065 (
            .O(N__18827),
            .I(cmd_rdadctmp_6));
    CascadeMux I__2064 (
            .O(N__18824),
            .I(N__18821));
    InMux I__2063 (
            .O(N__18821),
            .I(N__18815));
    InMux I__2062 (
            .O(N__18820),
            .I(N__18815));
    LocalMux I__2061 (
            .O(N__18815),
            .I(cmd_rdadctmp_5));
    CascadeMux I__2060 (
            .O(N__18812),
            .I(N__18808));
    CascadeMux I__2059 (
            .O(N__18811),
            .I(N__18805));
    InMux I__2058 (
            .O(N__18808),
            .I(N__18800));
    InMux I__2057 (
            .O(N__18805),
            .I(N__18800));
    LocalMux I__2056 (
            .O(N__18800),
            .I(cmd_rdadctmp_3));
    CascadeMux I__2055 (
            .O(N__18797),
            .I(N__18794));
    InMux I__2054 (
            .O(N__18794),
            .I(N__18788));
    InMux I__2053 (
            .O(N__18793),
            .I(N__18788));
    LocalMux I__2052 (
            .O(N__18788),
            .I(cmd_rdadctmp_4));
    InMux I__2051 (
            .O(N__18785),
            .I(N__18782));
    LocalMux I__2050 (
            .O(N__18782),
            .I(N__18779));
    Span12Mux_s10_h I__2049 (
            .O(N__18779),
            .I(N__18775));
    InMux I__2048 (
            .O(N__18778),
            .I(N__18772));
    Span12Mux_h I__2047 (
            .O(N__18775),
            .I(N__18769));
    LocalMux I__2046 (
            .O(N__18772),
            .I(buf_adcdata1_3));
    Odrv12 I__2045 (
            .O(N__18769),
            .I(buf_adcdata1_3));
    CascadeMux I__2044 (
            .O(N__18764),
            .I(N__18761));
    InMux I__2043 (
            .O(N__18761),
            .I(N__18757));
    InMux I__2042 (
            .O(N__18760),
            .I(N__18754));
    LocalMux I__2041 (
            .O(N__18757),
            .I(N__18750));
    LocalMux I__2040 (
            .O(N__18754),
            .I(N__18747));
    InMux I__2039 (
            .O(N__18753),
            .I(N__18744));
    Span4Mux_h I__2038 (
            .O(N__18750),
            .I(N__18739));
    Span4Mux_h I__2037 (
            .O(N__18747),
            .I(N__18739));
    LocalMux I__2036 (
            .O(N__18744),
            .I(buf_adcdata3_4));
    Odrv4 I__2035 (
            .O(N__18739),
            .I(buf_adcdata3_4));
    CascadeMux I__2034 (
            .O(N__18734),
            .I(N__18730));
    CascadeMux I__2033 (
            .O(N__18733),
            .I(N__18727));
    InMux I__2032 (
            .O(N__18730),
            .I(N__18722));
    InMux I__2031 (
            .O(N__18727),
            .I(N__18722));
    LocalMux I__2030 (
            .O(N__18722),
            .I(cmd_rdadctmp_1));
    InMux I__2029 (
            .O(N__18719),
            .I(N__18716));
    LocalMux I__2028 (
            .O(N__18716),
            .I(N__18712));
    CascadeMux I__2027 (
            .O(N__18715),
            .I(N__18709));
    Span4Mux_h I__2026 (
            .O(N__18712),
            .I(N__18705));
    InMux I__2025 (
            .O(N__18709),
            .I(N__18702));
    InMux I__2024 (
            .O(N__18708),
            .I(N__18699));
    Span4Mux_v I__2023 (
            .O(N__18705),
            .I(N__18696));
    LocalMux I__2022 (
            .O(N__18702),
            .I(N__18693));
    LocalMux I__2021 (
            .O(N__18699),
            .I(buf_adcdata3_7));
    Odrv4 I__2020 (
            .O(N__18696),
            .I(buf_adcdata3_7));
    Odrv12 I__2019 (
            .O(N__18693),
            .I(buf_adcdata3_7));
    CascadeMux I__2018 (
            .O(N__18686),
            .I(N__18683));
    InMux I__2017 (
            .O(N__18683),
            .I(N__18680));
    LocalMux I__2016 (
            .O(N__18680),
            .I(N__18677));
    Span4Mux_v I__2015 (
            .O(N__18677),
            .I(N__18674));
    Span4Mux_h I__2014 (
            .O(N__18674),
            .I(N__18671));
    Span4Mux_h I__2013 (
            .O(N__18671),
            .I(N__18668));
    Odrv4 I__2012 (
            .O(N__18668),
            .I(M_MISO1));
    InMux I__2011 (
            .O(N__18665),
            .I(N__18659));
    InMux I__2010 (
            .O(N__18664),
            .I(N__18659));
    LocalMux I__2009 (
            .O(N__18659),
            .I(cmd_rdadctmp_0));
    InMux I__2008 (
            .O(N__18656),
            .I(N__18652));
    CascadeMux I__2007 (
            .O(N__18655),
            .I(N__18649));
    LocalMux I__2006 (
            .O(N__18652),
            .I(N__18645));
    InMux I__2005 (
            .O(N__18649),
            .I(N__18640));
    InMux I__2004 (
            .O(N__18648),
            .I(N__18640));
    Odrv4 I__2003 (
            .O(N__18645),
            .I(cmd_rdadctmp_12_adj_1100));
    LocalMux I__2002 (
            .O(N__18640),
            .I(cmd_rdadctmp_12_adj_1100));
    InMux I__2001 (
            .O(N__18635),
            .I(N__18632));
    LocalMux I__2000 (
            .O(N__18632),
            .I(N__18629));
    Span4Mux_h I__1999 (
            .O(N__18629),
            .I(N__18625));
    InMux I__1998 (
            .O(N__18628),
            .I(N__18622));
    Span4Mux_v I__1997 (
            .O(N__18625),
            .I(N__18619));
    LocalMux I__1996 (
            .O(N__18622),
            .I(buf_adcdata1_4));
    Odrv4 I__1995 (
            .O(N__18619),
            .I(buf_adcdata1_4));
    SRMux I__1994 (
            .O(N__18614),
            .I(N__18609));
    SRMux I__1993 (
            .O(N__18613),
            .I(N__18606));
    SRMux I__1992 (
            .O(N__18612),
            .I(N__18603));
    LocalMux I__1991 (
            .O(N__18609),
            .I(N__18600));
    LocalMux I__1990 (
            .O(N__18606),
            .I(N__18597));
    LocalMux I__1989 (
            .O(N__18603),
            .I(N__18594));
    Span4Mux_h I__1988 (
            .O(N__18600),
            .I(N__18591));
    Odrv12 I__1987 (
            .O(N__18597),
            .I(n10590));
    Odrv12 I__1986 (
            .O(N__18594),
            .I(n10590));
    Odrv4 I__1985 (
            .O(N__18591),
            .I(n10590));
    InMux I__1984 (
            .O(N__18584),
            .I(N__18580));
    InMux I__1983 (
            .O(N__18583),
            .I(N__18577));
    LocalMux I__1982 (
            .O(N__18580),
            .I(N__18574));
    LocalMux I__1981 (
            .O(N__18577),
            .I(secclk_cnt_21));
    Odrv4 I__1980 (
            .O(N__18574),
            .I(secclk_cnt_21));
    InMux I__1979 (
            .O(N__18569),
            .I(N__18565));
    InMux I__1978 (
            .O(N__18568),
            .I(N__18562));
    LocalMux I__1977 (
            .O(N__18565),
            .I(N__18559));
    LocalMux I__1976 (
            .O(N__18562),
            .I(secclk_cnt_19));
    Odrv4 I__1975 (
            .O(N__18559),
            .I(secclk_cnt_19));
    CascadeMux I__1974 (
            .O(N__18554),
            .I(N__18551));
    InMux I__1973 (
            .O(N__18551),
            .I(N__18548));
    LocalMux I__1972 (
            .O(N__18548),
            .I(N__18544));
    InMux I__1971 (
            .O(N__18547),
            .I(N__18541));
    Span4Mux_v I__1970 (
            .O(N__18544),
            .I(N__18538));
    LocalMux I__1969 (
            .O(N__18541),
            .I(secclk_cnt_12));
    Odrv4 I__1968 (
            .O(N__18538),
            .I(secclk_cnt_12));
    InMux I__1967 (
            .O(N__18533),
            .I(N__18529));
    InMux I__1966 (
            .O(N__18532),
            .I(N__18526));
    LocalMux I__1965 (
            .O(N__18529),
            .I(N__18523));
    LocalMux I__1964 (
            .O(N__18526),
            .I(secclk_cnt_22));
    Odrv12 I__1963 (
            .O(N__18523),
            .I(secclk_cnt_22));
    InMux I__1962 (
            .O(N__18518),
            .I(N__18515));
    LocalMux I__1961 (
            .O(N__18515),
            .I(N__18512));
    Span12Mux_v I__1960 (
            .O(N__18512),
            .I(N__18509));
    Odrv12 I__1959 (
            .O(N__18509),
            .I(n14_adj_1163));
    InMux I__1958 (
            .O(N__18506),
            .I(N__18503));
    LocalMux I__1957 (
            .O(N__18503),
            .I(N__18500));
    Span4Mux_h I__1956 (
            .O(N__18500),
            .I(N__18497));
    Span4Mux_v I__1955 (
            .O(N__18497),
            .I(N__18494));
    Sp12to4 I__1954 (
            .O(N__18494),
            .I(N__18491));
    Span12Mux_v I__1953 (
            .O(N__18491),
            .I(N__18488));
    Odrv12 I__1952 (
            .O(N__18488),
            .I(buf_data2_10));
    CascadeMux I__1951 (
            .O(N__18485),
            .I(n4062_cascade_));
    InMux I__1950 (
            .O(N__18482),
            .I(N__18479));
    LocalMux I__1949 (
            .O(N__18479),
            .I(N__18476));
    Span4Mux_v I__1948 (
            .O(N__18476),
            .I(N__18472));
    CascadeMux I__1947 (
            .O(N__18475),
            .I(N__18469));
    Span4Mux_h I__1946 (
            .O(N__18472),
            .I(N__18466));
    InMux I__1945 (
            .O(N__18469),
            .I(N__18463));
    Span4Mux_h I__1944 (
            .O(N__18466),
            .I(N__18460));
    LocalMux I__1943 (
            .O(N__18463),
            .I(N__18454));
    Span4Mux_h I__1942 (
            .O(N__18460),
            .I(N__18454));
    InMux I__1941 (
            .O(N__18459),
            .I(N__18451));
    Span4Mux_h I__1940 (
            .O(N__18454),
            .I(N__18448));
    LocalMux I__1939 (
            .O(N__18451),
            .I(buf_adcdata3_2));
    Odrv4 I__1938 (
            .O(N__18448),
            .I(buf_adcdata3_2));
    CascadeMux I__1937 (
            .O(N__18443),
            .I(N__18439));
    InMux I__1936 (
            .O(N__18442),
            .I(N__18431));
    InMux I__1935 (
            .O(N__18439),
            .I(N__18431));
    InMux I__1934 (
            .O(N__18438),
            .I(N__18431));
    LocalMux I__1933 (
            .O(N__18431),
            .I(cmd_rdadctmp_11_adj_1101));
    CascadeMux I__1932 (
            .O(N__18428),
            .I(n8787_cascade_));
    InMux I__1931 (
            .O(N__18425),
            .I(N__18422));
    LocalMux I__1930 (
            .O(N__18422),
            .I(N__18419));
    Span4Mux_v I__1929 (
            .O(N__18419),
            .I(N__18416));
    Sp12to4 I__1928 (
            .O(N__18416),
            .I(N__18413));
    Span12Mux_h I__1927 (
            .O(N__18413),
            .I(N__18410));
    Odrv12 I__1926 (
            .O(N__18410),
            .I(buf_data1_2));
    CascadeMux I__1925 (
            .O(N__18407),
            .I(n4150_cascade_));
    InMux I__1924 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__1923 (
            .O(N__18401),
            .I(N__18398));
    Odrv12 I__1922 (
            .O(N__18398),
            .I(buf_data1_4));
    CascadeMux I__1921 (
            .O(N__18395),
            .I(n4148_cascade_));
    InMux I__1920 (
            .O(N__18392),
            .I(N__18389));
    LocalMux I__1919 (
            .O(N__18389),
            .I(N__18386));
    Span4Mux_h I__1918 (
            .O(N__18386),
            .I(N__18383));
    Odrv4 I__1917 (
            .O(N__18383),
            .I(buf_data1_5));
    CascadeMux I__1916 (
            .O(N__18380),
            .I(n4147_cascade_));
    CEMux I__1915 (
            .O(N__18377),
            .I(N__18372));
    CEMux I__1914 (
            .O(N__18376),
            .I(N__18369));
    CEMux I__1913 (
            .O(N__18375),
            .I(N__18366));
    LocalMux I__1912 (
            .O(N__18372),
            .I(n8738));
    LocalMux I__1911 (
            .O(N__18369),
            .I(n8738));
    LocalMux I__1910 (
            .O(N__18366),
            .I(n8738));
    InMux I__1909 (
            .O(N__18359),
            .I(N__18356));
    LocalMux I__1908 (
            .O(N__18356),
            .I(N__18353));
    Odrv4 I__1907 (
            .O(N__18353),
            .I(buf_data1_7));
    InMux I__1906 (
            .O(N__18350),
            .I(N__18347));
    LocalMux I__1905 (
            .O(N__18347),
            .I(N__18344));
    Odrv4 I__1904 (
            .O(N__18344),
            .I(n4145));
    InMux I__1903 (
            .O(N__18341),
            .I(N__18338));
    LocalMux I__1902 (
            .O(N__18338),
            .I(n4152));
    CascadeMux I__1901 (
            .O(N__18335),
            .I(n15131_cascade_));
    CascadeMux I__1900 (
            .O(N__18332),
            .I(n8738_cascade_));
    CEMux I__1899 (
            .O(N__18329),
            .I(N__18326));
    LocalMux I__1898 (
            .O(N__18326),
            .I(N__18322));
    CEMux I__1897 (
            .O(N__18325),
            .I(N__18319));
    Span4Mux_v I__1896 (
            .O(N__18322),
            .I(N__18316));
    LocalMux I__1895 (
            .O(N__18319),
            .I(N__18313));
    Span4Mux_h I__1894 (
            .O(N__18316),
            .I(N__18310));
    Span4Mux_h I__1893 (
            .O(N__18313),
            .I(N__18307));
    Odrv4 I__1892 (
            .O(N__18310),
            .I(n8847));
    Odrv4 I__1891 (
            .O(N__18307),
            .I(n8847));
    CascadeMux I__1890 (
            .O(N__18302),
            .I(n8847_cascade_));
    SRMux I__1889 (
            .O(N__18299),
            .I(N__18295));
    SRMux I__1888 (
            .O(N__18298),
            .I(N__18292));
    LocalMux I__1887 (
            .O(N__18295),
            .I(n10611));
    LocalMux I__1886 (
            .O(N__18292),
            .I(n10611));
    CascadeMux I__1885 (
            .O(N__18287),
            .I(N__18284));
    InMux I__1884 (
            .O(N__18284),
            .I(N__18278));
    InMux I__1883 (
            .O(N__18283),
            .I(N__18278));
    LocalMux I__1882 (
            .O(N__18278),
            .I(cmd_rdadctmp_7_adj_1142));
    CascadeMux I__1881 (
            .O(N__18275),
            .I(N__18271));
    CascadeMux I__1880 (
            .O(N__18274),
            .I(N__18268));
    InMux I__1879 (
            .O(N__18271),
            .I(N__18262));
    InMux I__1878 (
            .O(N__18268),
            .I(N__18262));
    InMux I__1877 (
            .O(N__18267),
            .I(N__18259));
    LocalMux I__1876 (
            .O(N__18262),
            .I(cmd_rdadctmp_8_adj_1141));
    LocalMux I__1875 (
            .O(N__18259),
            .I(cmd_rdadctmp_8_adj_1141));
    InMux I__1874 (
            .O(N__18254),
            .I(N__18250));
    InMux I__1873 (
            .O(N__18253),
            .I(N__18247));
    LocalMux I__1872 (
            .O(N__18250),
            .I(cmd_rdadctmp_5_adj_1144));
    LocalMux I__1871 (
            .O(N__18247),
            .I(cmd_rdadctmp_5_adj_1144));
    InMux I__1870 (
            .O(N__18242),
            .I(N__18236));
    InMux I__1869 (
            .O(N__18241),
            .I(N__18236));
    LocalMux I__1868 (
            .O(N__18236),
            .I(cmd_rdadctmp_6_adj_1143));
    CascadeMux I__1867 (
            .O(N__18233),
            .I(N__18230));
    InMux I__1866 (
            .O(N__18230),
            .I(N__18227));
    LocalMux I__1865 (
            .O(N__18227),
            .I(N__18224));
    Span4Mux_h I__1864 (
            .O(N__18224),
            .I(N__18221));
    Span4Mux_v I__1863 (
            .O(N__18221),
            .I(N__18216));
    InMux I__1862 (
            .O(N__18220),
            .I(N__18213));
    InMux I__1861 (
            .O(N__18219),
            .I(N__18210));
    Odrv4 I__1860 (
            .O(N__18216),
            .I(cmd_rdadctmp_11_adj_1138));
    LocalMux I__1859 (
            .O(N__18213),
            .I(cmd_rdadctmp_11_adj_1138));
    LocalMux I__1858 (
            .O(N__18210),
            .I(cmd_rdadctmp_11_adj_1138));
    CascadeMux I__1857 (
            .O(N__18203),
            .I(N__18199));
    InMux I__1856 (
            .O(N__18202),
            .I(N__18196));
    InMux I__1855 (
            .O(N__18199),
            .I(N__18193));
    LocalMux I__1854 (
            .O(N__18196),
            .I(cmd_rdadctmp_4_adj_1145));
    LocalMux I__1853 (
            .O(N__18193),
            .I(cmd_rdadctmp_4_adj_1145));
    CascadeMux I__1852 (
            .O(N__18188),
            .I(N__18184));
    InMux I__1851 (
            .O(N__18187),
            .I(N__18179));
    InMux I__1850 (
            .O(N__18184),
            .I(N__18179));
    LocalMux I__1849 (
            .O(N__18179),
            .I(cmd_rdadctmp_3_adj_1146));
    CascadeMux I__1848 (
            .O(N__18176),
            .I(N__18172));
    InMux I__1847 (
            .O(N__18175),
            .I(N__18169));
    InMux I__1846 (
            .O(N__18172),
            .I(N__18166));
    LocalMux I__1845 (
            .O(N__18169),
            .I(cmd_rdadctmp_2_adj_1147));
    LocalMux I__1844 (
            .O(N__18166),
            .I(cmd_rdadctmp_2_adj_1147));
    CascadeMux I__1843 (
            .O(N__18161),
            .I(N__18158));
    InMux I__1842 (
            .O(N__18158),
            .I(N__18155));
    LocalMux I__1841 (
            .O(N__18155),
            .I(N__18152));
    Span4Mux_v I__1840 (
            .O(N__18152),
            .I(N__18147));
    InMux I__1839 (
            .O(N__18151),
            .I(N__18144));
    CascadeMux I__1838 (
            .O(N__18150),
            .I(N__18141));
    Span4Mux_v I__1837 (
            .O(N__18147),
            .I(N__18138));
    LocalMux I__1836 (
            .O(N__18144),
            .I(N__18135));
    InMux I__1835 (
            .O(N__18141),
            .I(N__18132));
    Odrv4 I__1834 (
            .O(N__18138),
            .I(cmd_rdadctmp_12_adj_1137));
    Odrv4 I__1833 (
            .O(N__18135),
            .I(cmd_rdadctmp_12_adj_1137));
    LocalMux I__1832 (
            .O(N__18132),
            .I(cmd_rdadctmp_12_adj_1137));
    InMux I__1831 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__1830 (
            .O(N__18122),
            .I(N__18117));
    InMux I__1829 (
            .O(N__18121),
            .I(N__18114));
    InMux I__1828 (
            .O(N__18120),
            .I(N__18111));
    Span4Mux_v I__1827 (
            .O(N__18117),
            .I(N__18108));
    LocalMux I__1826 (
            .O(N__18114),
            .I(buf_adcdata4_4));
    LocalMux I__1825 (
            .O(N__18111),
            .I(buf_adcdata4_4));
    Odrv4 I__1824 (
            .O(N__18108),
            .I(buf_adcdata4_4));
    InMux I__1823 (
            .O(N__18101),
            .I(N__18098));
    LocalMux I__1822 (
            .O(N__18098),
            .I(N__18095));
    Span4Mux_v I__1821 (
            .O(N__18095),
            .I(N__18092));
    Odrv4 I__1820 (
            .O(N__18092),
            .I(buf_data1_6));
    InMux I__1819 (
            .O(N__18089),
            .I(N__18086));
    LocalMux I__1818 (
            .O(N__18086),
            .I(N__18083));
    Span4Mux_h I__1817 (
            .O(N__18083),
            .I(N__18080));
    Odrv4 I__1816 (
            .O(N__18080),
            .I(n4146));
    InMux I__1815 (
            .O(N__18077),
            .I(N__18074));
    LocalMux I__1814 (
            .O(N__18074),
            .I(N__18071));
    Span4Mux_h I__1813 (
            .O(N__18071),
            .I(N__18068));
    Sp12to4 I__1812 (
            .O(N__18068),
            .I(N__18065));
    Span12Mux_h I__1811 (
            .O(N__18065),
            .I(N__18062));
    Odrv12 I__1810 (
            .O(N__18062),
            .I(buf_data1_0));
    InMux I__1809 (
            .O(N__18059),
            .I(N__18056));
    LocalMux I__1808 (
            .O(N__18056),
            .I(N__18051));
    InMux I__1807 (
            .O(N__18055),
            .I(N__18048));
    CascadeMux I__1806 (
            .O(N__18054),
            .I(N__18045));
    Span4Mux_v I__1805 (
            .O(N__18051),
            .I(N__18042));
    LocalMux I__1804 (
            .O(N__18048),
            .I(N__18039));
    InMux I__1803 (
            .O(N__18045),
            .I(N__18036));
    Odrv4 I__1802 (
            .O(N__18042),
            .I(cmd_rdadctmp_15_adj_1134));
    Odrv4 I__1801 (
            .O(N__18039),
            .I(cmd_rdadctmp_15_adj_1134));
    LocalMux I__1800 (
            .O(N__18036),
            .I(cmd_rdadctmp_15_adj_1134));
    InMux I__1799 (
            .O(N__18029),
            .I(N__18026));
    LocalMux I__1798 (
            .O(N__18026),
            .I(N__18023));
    Span4Mux_v I__1797 (
            .O(N__18023),
            .I(N__18020));
    Span4Mux_v I__1796 (
            .O(N__18020),
            .I(N__18017));
    Sp12to4 I__1795 (
            .O(N__18017),
            .I(N__18012));
    InMux I__1794 (
            .O(N__18016),
            .I(N__18009));
    InMux I__1793 (
            .O(N__18015),
            .I(N__18006));
    Span12Mux_h I__1792 (
            .O(N__18012),
            .I(N__18003));
    LocalMux I__1791 (
            .O(N__18009),
            .I(N__18000));
    LocalMux I__1790 (
            .O(N__18006),
            .I(buf_adcdata4_0));
    Odrv12 I__1789 (
            .O(N__18003),
            .I(buf_adcdata4_0));
    Odrv12 I__1788 (
            .O(N__18000),
            .I(buf_adcdata4_0));
    InMux I__1787 (
            .O(N__17993),
            .I(N__17990));
    LocalMux I__1786 (
            .O(N__17990),
            .I(N__17987));
    Span4Mux_v I__1785 (
            .O(N__17987),
            .I(N__17983));
    CascadeMux I__1784 (
            .O(N__17986),
            .I(N__17980));
    Span4Mux_v I__1783 (
            .O(N__17983),
            .I(N__17977));
    InMux I__1782 (
            .O(N__17980),
            .I(N__17973));
    Sp12to4 I__1781 (
            .O(N__17977),
            .I(N__17970));
    InMux I__1780 (
            .O(N__17976),
            .I(N__17967));
    LocalMux I__1779 (
            .O(N__17973),
            .I(N__17964));
    Span12Mux_h I__1778 (
            .O(N__17970),
            .I(N__17961));
    LocalMux I__1777 (
            .O(N__17967),
            .I(buf_adcdata4_1));
    Odrv12 I__1776 (
            .O(N__17964),
            .I(buf_adcdata4_1));
    Odrv12 I__1775 (
            .O(N__17961),
            .I(buf_adcdata4_1));
    CascadeMux I__1774 (
            .O(N__17954),
            .I(N__17950));
    CascadeMux I__1773 (
            .O(N__17953),
            .I(N__17947));
    InMux I__1772 (
            .O(N__17950),
            .I(N__17939));
    InMux I__1771 (
            .O(N__17947),
            .I(N__17939));
    InMux I__1770 (
            .O(N__17946),
            .I(N__17939));
    LocalMux I__1769 (
            .O(N__17939),
            .I(cmd_rdadctmp_9_adj_1140));
    CascadeMux I__1768 (
            .O(N__17936),
            .I(N__17932));
    InMux I__1767 (
            .O(N__17935),
            .I(N__17924));
    InMux I__1766 (
            .O(N__17932),
            .I(N__17924));
    InMux I__1765 (
            .O(N__17931),
            .I(N__17924));
    LocalMux I__1764 (
            .O(N__17924),
            .I(cmd_rdadctmp_10_adj_1139));
    InMux I__1763 (
            .O(N__17921),
            .I(N__17918));
    LocalMux I__1762 (
            .O(N__17918),
            .I(N__17915));
    Span4Mux_v I__1761 (
            .O(N__17915),
            .I(N__17911));
    InMux I__1760 (
            .O(N__17914),
            .I(N__17907));
    Sp12to4 I__1759 (
            .O(N__17911),
            .I(N__17904));
    CascadeMux I__1758 (
            .O(N__17910),
            .I(N__17901));
    LocalMux I__1757 (
            .O(N__17907),
            .I(N__17896));
    Span12Mux_s11_h I__1756 (
            .O(N__17904),
            .I(N__17896));
    InMux I__1755 (
            .O(N__17901),
            .I(N__17893));
    Span12Mux_h I__1754 (
            .O(N__17896),
            .I(N__17890));
    LocalMux I__1753 (
            .O(N__17893),
            .I(buf_adcdata4_2));
    Odrv12 I__1752 (
            .O(N__17890),
            .I(buf_adcdata4_2));
    InMux I__1751 (
            .O(N__17885),
            .I(N__17881));
    InMux I__1750 (
            .O(N__17884),
            .I(N__17878));
    LocalMux I__1749 (
            .O(N__17881),
            .I(N__17875));
    LocalMux I__1748 (
            .O(N__17878),
            .I(buf_adcdata2_4));
    Odrv4 I__1747 (
            .O(N__17875),
            .I(buf_adcdata2_4));
    CascadeMux I__1746 (
            .O(N__17870),
            .I(N__17865));
    CascadeMux I__1745 (
            .O(N__17869),
            .I(N__17862));
    CascadeMux I__1744 (
            .O(N__17868),
            .I(N__17859));
    InMux I__1743 (
            .O(N__17865),
            .I(N__17856));
    InMux I__1742 (
            .O(N__17862),
            .I(N__17851));
    InMux I__1741 (
            .O(N__17859),
            .I(N__17851));
    LocalMux I__1740 (
            .O(N__17856),
            .I(cmd_rdadctmp_13_adj_1063));
    LocalMux I__1739 (
            .O(N__17851),
            .I(cmd_rdadctmp_13_adj_1063));
    InMux I__1738 (
            .O(N__17846),
            .I(N__17839));
    InMux I__1737 (
            .O(N__17845),
            .I(N__17839));
    InMux I__1736 (
            .O(N__17844),
            .I(N__17836));
    LocalMux I__1735 (
            .O(N__17839),
            .I(cmd_rdadctmp_14_adj_1062));
    LocalMux I__1734 (
            .O(N__17836),
            .I(cmd_rdadctmp_14_adj_1062));
    CascadeMux I__1733 (
            .O(N__17831),
            .I(N__17826));
    InMux I__1732 (
            .O(N__17830),
            .I(N__17823));
    InMux I__1731 (
            .O(N__17829),
            .I(N__17818));
    InMux I__1730 (
            .O(N__17826),
            .I(N__17818));
    LocalMux I__1729 (
            .O(N__17823),
            .I(cmd_rdadctmp_11_adj_1065));
    LocalMux I__1728 (
            .O(N__17818),
            .I(cmd_rdadctmp_11_adj_1065));
    CascadeMux I__1727 (
            .O(N__17813),
            .I(N__17809));
    CascadeMux I__1726 (
            .O(N__17812),
            .I(N__17805));
    InMux I__1725 (
            .O(N__17809),
            .I(N__17800));
    InMux I__1724 (
            .O(N__17808),
            .I(N__17800));
    InMux I__1723 (
            .O(N__17805),
            .I(N__17797));
    LocalMux I__1722 (
            .O(N__17800),
            .I(cmd_rdadctmp_12_adj_1064));
    LocalMux I__1721 (
            .O(N__17797),
            .I(cmd_rdadctmp_12_adj_1064));
    InMux I__1720 (
            .O(N__17792),
            .I(N__17789));
    LocalMux I__1719 (
            .O(N__17789),
            .I(N__17785));
    InMux I__1718 (
            .O(N__17788),
            .I(N__17782));
    Span4Mux_v I__1717 (
            .O(N__17785),
            .I(N__17779));
    LocalMux I__1716 (
            .O(N__17782),
            .I(buf_adcdata1_5));
    Odrv4 I__1715 (
            .O(N__17779),
            .I(buf_adcdata1_5));
    InMux I__1714 (
            .O(N__17774),
            .I(N__17771));
    LocalMux I__1713 (
            .O(N__17771),
            .I(N__17767));
    InMux I__1712 (
            .O(N__17770),
            .I(N__17764));
    Span4Mux_v I__1711 (
            .O(N__17767),
            .I(N__17761));
    LocalMux I__1710 (
            .O(N__17764),
            .I(buf_adcdata1_7));
    Odrv4 I__1709 (
            .O(N__17761),
            .I(buf_adcdata1_7));
    CascadeMux I__1708 (
            .O(N__17756),
            .I(N__17753));
    InMux I__1707 (
            .O(N__17753),
            .I(N__17749));
    InMux I__1706 (
            .O(N__17752),
            .I(N__17746));
    LocalMux I__1705 (
            .O(N__17749),
            .I(N__17740));
    LocalMux I__1704 (
            .O(N__17746),
            .I(N__17740));
    InMux I__1703 (
            .O(N__17745),
            .I(N__17737));
    Span4Mux_v I__1702 (
            .O(N__17740),
            .I(N__17734));
    LocalMux I__1701 (
            .O(N__17737),
            .I(buf_adcdata4_5));
    Odrv4 I__1700 (
            .O(N__17734),
            .I(buf_adcdata4_5));
    CascadeMux I__1699 (
            .O(N__17729),
            .I(N__17724));
    InMux I__1698 (
            .O(N__17728),
            .I(N__17717));
    InMux I__1697 (
            .O(N__17727),
            .I(N__17717));
    InMux I__1696 (
            .O(N__17724),
            .I(N__17717));
    LocalMux I__1695 (
            .O(N__17717),
            .I(cmd_rdadctmp_13_adj_1136));
    InMux I__1694 (
            .O(N__17714),
            .I(N__17711));
    LocalMux I__1693 (
            .O(N__17711),
            .I(N__17706));
    CascadeMux I__1692 (
            .O(N__17710),
            .I(N__17703));
    CascadeMux I__1691 (
            .O(N__17709),
            .I(N__17700));
    Span4Mux_h I__1690 (
            .O(N__17706),
            .I(N__17697));
    InMux I__1689 (
            .O(N__17703),
            .I(N__17692));
    InMux I__1688 (
            .O(N__17700),
            .I(N__17692));
    Odrv4 I__1687 (
            .O(N__17697),
            .I(cmd_rdadctmp_14_adj_1135));
    LocalMux I__1686 (
            .O(N__17692),
            .I(cmd_rdadctmp_14_adj_1135));
    CascadeMux I__1685 (
            .O(N__17687),
            .I(N__17684));
    InMux I__1684 (
            .O(N__17684),
            .I(N__17681));
    LocalMux I__1683 (
            .O(N__17681),
            .I(N__17677));
    InMux I__1682 (
            .O(N__17680),
            .I(N__17674));
    Span4Mux_h I__1681 (
            .O(N__17677),
            .I(N__17668));
    LocalMux I__1680 (
            .O(N__17674),
            .I(N__17668));
    InMux I__1679 (
            .O(N__17673),
            .I(N__17665));
    Span4Mux_v I__1678 (
            .O(N__17668),
            .I(N__17662));
    LocalMux I__1677 (
            .O(N__17665),
            .I(buf_adcdata4_6));
    Odrv4 I__1676 (
            .O(N__17662),
            .I(buf_adcdata4_6));
    InMux I__1675 (
            .O(N__17657),
            .I(N__17654));
    LocalMux I__1674 (
            .O(N__17654),
            .I(N__17650));
    InMux I__1673 (
            .O(N__17653),
            .I(N__17647));
    Span4Mux_h I__1672 (
            .O(N__17650),
            .I(N__17644));
    LocalMux I__1671 (
            .O(N__17647),
            .I(buf_adcdata2_5));
    Odrv4 I__1670 (
            .O(N__17644),
            .I(buf_adcdata2_5));
    InMux I__1669 (
            .O(N__17639),
            .I(N__17635));
    CascadeMux I__1668 (
            .O(N__17638),
            .I(N__17632));
    LocalMux I__1667 (
            .O(N__17635),
            .I(N__17629));
    InMux I__1666 (
            .O(N__17632),
            .I(N__17626));
    Span4Mux_h I__1665 (
            .O(N__17629),
            .I(N__17623));
    LocalMux I__1664 (
            .O(N__17626),
            .I(buf_adcdata2_6));
    Odrv4 I__1663 (
            .O(N__17623),
            .I(buf_adcdata2_6));
    InMux I__1662 (
            .O(N__17618),
            .I(N__17614));
    CascadeMux I__1661 (
            .O(N__17617),
            .I(N__17611));
    LocalMux I__1660 (
            .O(N__17614),
            .I(N__17608));
    InMux I__1659 (
            .O(N__17611),
            .I(N__17605));
    Span4Mux_h I__1658 (
            .O(N__17608),
            .I(N__17602));
    LocalMux I__1657 (
            .O(N__17605),
            .I(buf_adcdata2_7));
    Odrv4 I__1656 (
            .O(N__17602),
            .I(buf_adcdata2_7));
    CascadeMux I__1655 (
            .O(N__17597),
            .I(N__17592));
    InMux I__1654 (
            .O(N__17596),
            .I(N__17585));
    InMux I__1653 (
            .O(N__17595),
            .I(N__17585));
    InMux I__1652 (
            .O(N__17592),
            .I(N__17585));
    LocalMux I__1651 (
            .O(N__17585),
            .I(cmd_rdadctmp_15_adj_1061));
    InMux I__1650 (
            .O(N__17582),
            .I(N__17579));
    LocalMux I__1649 (
            .O(N__17579),
            .I(N__17576));
    Span4Mux_v I__1648 (
            .O(N__17576),
            .I(N__17573));
    Span4Mux_v I__1647 (
            .O(N__17573),
            .I(N__17569));
    CascadeMux I__1646 (
            .O(N__17572),
            .I(N__17566));
    Sp12to4 I__1645 (
            .O(N__17569),
            .I(N__17563));
    InMux I__1644 (
            .O(N__17566),
            .I(N__17560));
    Span12Mux_h I__1643 (
            .O(N__17563),
            .I(N__17557));
    LocalMux I__1642 (
            .O(N__17560),
            .I(buf_adcdata2_3));
    Odrv12 I__1641 (
            .O(N__17557),
            .I(buf_adcdata2_3));
    InMux I__1640 (
            .O(N__17552),
            .I(N__17549));
    LocalMux I__1639 (
            .O(N__17549),
            .I(n4301));
    InMux I__1638 (
            .O(N__17546),
            .I(N__17543));
    LocalMux I__1637 (
            .O(N__17543),
            .I(N__17540));
    Sp12to4 I__1636 (
            .O(N__17540),
            .I(N__17537));
    Span12Mux_v I__1635 (
            .O(N__17537),
            .I(N__17534));
    Span12Mux_h I__1634 (
            .O(N__17534),
            .I(N__17531));
    Odrv12 I__1633 (
            .O(N__17531),
            .I(buf_data2_0));
    InMux I__1632 (
            .O(N__17528),
            .I(N__17525));
    LocalMux I__1631 (
            .O(N__17525),
            .I(N__17522));
    Span12Mux_h I__1630 (
            .O(N__17522),
            .I(N__17519));
    Odrv12 I__1629 (
            .O(N__17519),
            .I(buf_data2_1));
    InMux I__1628 (
            .O(N__17516),
            .I(N__17513));
    LocalMux I__1627 (
            .O(N__17513),
            .I(N__17510));
    Span4Mux_v I__1626 (
            .O(N__17510),
            .I(N__17507));
    Sp12to4 I__1625 (
            .O(N__17507),
            .I(N__17504));
    Span12Mux_h I__1624 (
            .O(N__17504),
            .I(N__17501));
    Odrv12 I__1623 (
            .O(N__17501),
            .I(buf_data2_2));
    InMux I__1622 (
            .O(N__17498),
            .I(N__17495));
    LocalMux I__1621 (
            .O(N__17495),
            .I(n4307));
    InMux I__1620 (
            .O(N__17492),
            .I(N__17489));
    LocalMux I__1619 (
            .O(N__17489),
            .I(n4306));
    InMux I__1618 (
            .O(N__17486),
            .I(N__17483));
    LocalMux I__1617 (
            .O(N__17483),
            .I(n4308));
    InMux I__1616 (
            .O(N__17480),
            .I(N__17477));
    LocalMux I__1615 (
            .O(N__17477),
            .I(buf_data2_6));
    InMux I__1614 (
            .O(N__17474),
            .I(N__17469));
    InMux I__1613 (
            .O(N__17473),
            .I(N__17464));
    InMux I__1612 (
            .O(N__17472),
            .I(N__17464));
    LocalMux I__1611 (
            .O(N__17469),
            .I(buf_adcdata4_7));
    LocalMux I__1610 (
            .O(N__17464),
            .I(buf_adcdata4_7));
    InMux I__1609 (
            .O(N__17459),
            .I(N__17456));
    LocalMux I__1608 (
            .O(N__17456),
            .I(buf_data2_7));
    CascadeMux I__1607 (
            .O(N__17453),
            .I(N__17450));
    InMux I__1606 (
            .O(N__17450),
            .I(N__17447));
    LocalMux I__1605 (
            .O(N__17447),
            .I(N__17444));
    Odrv4 I__1604 (
            .O(N__17444),
            .I(buf_data2_4));
    CascadeMux I__1603 (
            .O(N__17441),
            .I(n4304_cascade_));
    InMux I__1602 (
            .O(N__17438),
            .I(N__17435));
    LocalMux I__1601 (
            .O(N__17435),
            .I(buf_data2_5));
    CascadeMux I__1600 (
            .O(N__17432),
            .I(n4303_cascade_));
    InMux I__1599 (
            .O(N__17429),
            .I(N__17426));
    LocalMux I__1598 (
            .O(N__17426),
            .I(n4302));
    CascadeMux I__1597 (
            .O(N__17423),
            .I(N__17419));
    InMux I__1596 (
            .O(N__17422),
            .I(N__17414));
    InMux I__1595 (
            .O(N__17419),
            .I(N__17414));
    LocalMux I__1594 (
            .O(N__17414),
            .I(cmd_rdadctmp_5_adj_1071));
    CascadeMux I__1593 (
            .O(N__17411),
            .I(N__17407));
    InMux I__1592 (
            .O(N__17410),
            .I(N__17402));
    InMux I__1591 (
            .O(N__17407),
            .I(N__17402));
    LocalMux I__1590 (
            .O(N__17402),
            .I(cmd_rdadctmp_3_adj_1073));
    InMux I__1589 (
            .O(N__17399),
            .I(N__17393));
    InMux I__1588 (
            .O(N__17398),
            .I(N__17393));
    LocalMux I__1587 (
            .O(N__17393),
            .I(cmd_rdadctmp_4_adj_1072));
    CascadeMux I__1586 (
            .O(N__17390),
            .I(n14_adj_1035_cascade_));
    IoInMux I__1585 (
            .O(N__17387),
            .I(N__17384));
    LocalMux I__1584 (
            .O(N__17384),
            .I(N__17381));
    IoSpan4Mux I__1583 (
            .O(N__17381),
            .I(N__17378));
    Span4Mux_s2_h I__1582 (
            .O(N__17378),
            .I(N__17374));
    CascadeMux I__1581 (
            .O(N__17377),
            .I(N__17371));
    Span4Mux_h I__1580 (
            .O(N__17374),
            .I(N__17368));
    InMux I__1579 (
            .O(N__17371),
            .I(N__17365));
    Odrv4 I__1578 (
            .O(N__17368),
            .I(M_CS2));
    LocalMux I__1577 (
            .O(N__17365),
            .I(M_CS2));
    InMux I__1576 (
            .O(N__17360),
            .I(N__17356));
    InMux I__1575 (
            .O(N__17359),
            .I(N__17353));
    LocalMux I__1574 (
            .O(N__17356),
            .I(n15165));
    LocalMux I__1573 (
            .O(N__17353),
            .I(n15165));
    InMux I__1572 (
            .O(N__17348),
            .I(N__17345));
    LocalMux I__1571 (
            .O(N__17345),
            .I(N__17342));
    Span4Mux_v I__1570 (
            .O(N__17342),
            .I(N__17339));
    Span4Mux_v I__1569 (
            .O(N__17339),
            .I(N__17336));
    Span4Mux_h I__1568 (
            .O(N__17336),
            .I(N__17333));
    Odrv4 I__1567 (
            .O(N__17333),
            .I(M_MISO2));
    CascadeMux I__1566 (
            .O(N__17330),
            .I(n8302_cascade_));
    InMux I__1565 (
            .O(N__17327),
            .I(N__17323));
    CascadeMux I__1564 (
            .O(N__17326),
            .I(N__17320));
    LocalMux I__1563 (
            .O(N__17323),
            .I(N__17317));
    InMux I__1562 (
            .O(N__17320),
            .I(N__17314));
    Odrv4 I__1561 (
            .O(N__17317),
            .I(cmd_rdadctmp_2_adj_1074));
    LocalMux I__1560 (
            .O(N__17314),
            .I(cmd_rdadctmp_2_adj_1074));
    InMux I__1559 (
            .O(N__17309),
            .I(N__17303));
    InMux I__1558 (
            .O(N__17308),
            .I(N__17303));
    LocalMux I__1557 (
            .O(N__17303),
            .I(cmd_rdadctmp_0_adj_1076));
    CascadeMux I__1556 (
            .O(N__17300),
            .I(N__17296));
    InMux I__1555 (
            .O(N__17299),
            .I(N__17291));
    InMux I__1554 (
            .O(N__17296),
            .I(N__17291));
    LocalMux I__1553 (
            .O(N__17291),
            .I(cmd_rdadctmp_1_adj_1075));
    InMux I__1552 (
            .O(N__17288),
            .I(n14029));
    InMux I__1551 (
            .O(N__17285),
            .I(n14030));
    InMux I__1550 (
            .O(N__17282),
            .I(N__17279));
    LocalMux I__1549 (
            .O(N__17279),
            .I(N__17272));
    ClkMux I__1548 (
            .O(N__17278),
            .I(N__17261));
    ClkMux I__1547 (
            .O(N__17277),
            .I(N__17261));
    ClkMux I__1546 (
            .O(N__17276),
            .I(N__17261));
    ClkMux I__1545 (
            .O(N__17275),
            .I(N__17261));
    Glb2LocalMux I__1544 (
            .O(N__17272),
            .I(N__17261));
    GlobalMux I__1543 (
            .O(N__17261),
            .I(clk_16MHz));
    SRMux I__1542 (
            .O(N__17258),
            .I(N__17254));
    SRMux I__1541 (
            .O(N__17257),
            .I(N__17251));
    LocalMux I__1540 (
            .O(N__17254),
            .I(N__17247));
    LocalMux I__1539 (
            .O(N__17251),
            .I(N__17244));
    SRMux I__1538 (
            .O(N__17250),
            .I(N__17241));
    Span4Mux_h I__1537 (
            .O(N__17247),
            .I(N__17238));
    Span4Mux_h I__1536 (
            .O(N__17244),
            .I(N__17235));
    LocalMux I__1535 (
            .O(N__17241),
            .I(N__17232));
    Odrv4 I__1534 (
            .O(N__17238),
            .I(n10522));
    Odrv4 I__1533 (
            .O(N__17235),
            .I(n10522));
    Odrv4 I__1532 (
            .O(N__17232),
            .I(n10522));
    InMux I__1531 (
            .O(N__17225),
            .I(N__17222));
    LocalMux I__1530 (
            .O(N__17222),
            .I(N__17219));
    Span4Mux_v I__1529 (
            .O(N__17219),
            .I(N__17216));
    Sp12to4 I__1528 (
            .O(N__17216),
            .I(N__17212));
    CascadeMux I__1527 (
            .O(N__17215),
            .I(N__17209));
    Span12Mux_h I__1526 (
            .O(N__17212),
            .I(N__17206));
    InMux I__1525 (
            .O(N__17209),
            .I(N__17203));
    Span12Mux_h I__1524 (
            .O(N__17206),
            .I(N__17200));
    LocalMux I__1523 (
            .O(N__17203),
            .I(buf_adcdata2_0));
    Odrv12 I__1522 (
            .O(N__17200),
            .I(buf_adcdata2_0));
    InMux I__1521 (
            .O(N__17195),
            .I(N__17186));
    InMux I__1520 (
            .O(N__17194),
            .I(N__17186));
    InMux I__1519 (
            .O(N__17193),
            .I(N__17186));
    LocalMux I__1518 (
            .O(N__17186),
            .I(cmd_rdadctmp_8_adj_1068));
    CascadeMux I__1517 (
            .O(N__17183),
            .I(N__17180));
    InMux I__1516 (
            .O(N__17180),
            .I(N__17174));
    InMux I__1515 (
            .O(N__17179),
            .I(N__17174));
    LocalMux I__1514 (
            .O(N__17174),
            .I(cmd_rdadctmp_7_adj_1069));
    CascadeMux I__1513 (
            .O(N__17171),
            .I(N__17168));
    InMux I__1512 (
            .O(N__17168),
            .I(N__17165));
    LocalMux I__1511 (
            .O(N__17165),
            .I(N__17161));
    InMux I__1510 (
            .O(N__17164),
            .I(N__17158));
    Odrv4 I__1509 (
            .O(N__17161),
            .I(cmd_rdadctmp_6_adj_1070));
    LocalMux I__1508 (
            .O(N__17158),
            .I(cmd_rdadctmp_6_adj_1070));
    CascadeMux I__1507 (
            .O(N__17153),
            .I(N__17150));
    InMux I__1506 (
            .O(N__17150),
            .I(N__17146));
    InMux I__1505 (
            .O(N__17149),
            .I(N__17143));
    LocalMux I__1504 (
            .O(N__17146),
            .I(N__17140));
    LocalMux I__1503 (
            .O(N__17143),
            .I(secclk_cnt_13));
    Odrv4 I__1502 (
            .O(N__17140),
            .I(secclk_cnt_13));
    InMux I__1501 (
            .O(N__17135),
            .I(n14021));
    InMux I__1500 (
            .O(N__17132),
            .I(N__17128));
    InMux I__1499 (
            .O(N__17131),
            .I(N__17125));
    LocalMux I__1498 (
            .O(N__17128),
            .I(secclk_cnt_14));
    LocalMux I__1497 (
            .O(N__17125),
            .I(secclk_cnt_14));
    InMux I__1496 (
            .O(N__17120),
            .I(n14022));
    InMux I__1495 (
            .O(N__17117),
            .I(N__17113));
    InMux I__1494 (
            .O(N__17116),
            .I(N__17110));
    LocalMux I__1493 (
            .O(N__17113),
            .I(secclk_cnt_15));
    LocalMux I__1492 (
            .O(N__17110),
            .I(secclk_cnt_15));
    InMux I__1491 (
            .O(N__17105),
            .I(n14023));
    InMux I__1490 (
            .O(N__17102),
            .I(N__17098));
    InMux I__1489 (
            .O(N__17101),
            .I(N__17095));
    LocalMux I__1488 (
            .O(N__17098),
            .I(N__17092));
    LocalMux I__1487 (
            .O(N__17095),
            .I(secclk_cnt_16));
    Odrv4 I__1486 (
            .O(N__17092),
            .I(secclk_cnt_16));
    InMux I__1485 (
            .O(N__17087),
            .I(bfn_3_9_0_));
    InMux I__1484 (
            .O(N__17084),
            .I(N__17080));
    InMux I__1483 (
            .O(N__17083),
            .I(N__17077));
    LocalMux I__1482 (
            .O(N__17080),
            .I(secclk_cnt_17));
    LocalMux I__1481 (
            .O(N__17077),
            .I(secclk_cnt_17));
    InMux I__1480 (
            .O(N__17072),
            .I(n14025));
    InMux I__1479 (
            .O(N__17069),
            .I(N__17065));
    InMux I__1478 (
            .O(N__17068),
            .I(N__17062));
    LocalMux I__1477 (
            .O(N__17065),
            .I(secclk_cnt_18));
    LocalMux I__1476 (
            .O(N__17062),
            .I(secclk_cnt_18));
    InMux I__1475 (
            .O(N__17057),
            .I(n14026));
    InMux I__1474 (
            .O(N__17054),
            .I(n14027));
    InMux I__1473 (
            .O(N__17051),
            .I(N__17047));
    InMux I__1472 (
            .O(N__17050),
            .I(N__17044));
    LocalMux I__1471 (
            .O(N__17047),
            .I(secclk_cnt_20));
    LocalMux I__1470 (
            .O(N__17044),
            .I(secclk_cnt_20));
    InMux I__1469 (
            .O(N__17039),
            .I(n14028));
    InMux I__1468 (
            .O(N__17036),
            .I(N__17032));
    InMux I__1467 (
            .O(N__17035),
            .I(N__17029));
    LocalMux I__1466 (
            .O(N__17032),
            .I(secclk_cnt_4));
    LocalMux I__1465 (
            .O(N__17029),
            .I(secclk_cnt_4));
    InMux I__1464 (
            .O(N__17024),
            .I(n14012));
    InMux I__1463 (
            .O(N__17021),
            .I(N__17017));
    InMux I__1462 (
            .O(N__17020),
            .I(N__17014));
    LocalMux I__1461 (
            .O(N__17017),
            .I(secclk_cnt_5));
    LocalMux I__1460 (
            .O(N__17014),
            .I(secclk_cnt_5));
    InMux I__1459 (
            .O(N__17009),
            .I(n14013));
    InMux I__1458 (
            .O(N__17006),
            .I(N__17002));
    InMux I__1457 (
            .O(N__17005),
            .I(N__16999));
    LocalMux I__1456 (
            .O(N__17002),
            .I(secclk_cnt_6));
    LocalMux I__1455 (
            .O(N__16999),
            .I(secclk_cnt_6));
    InMux I__1454 (
            .O(N__16994),
            .I(n14014));
    InMux I__1453 (
            .O(N__16991),
            .I(N__16987));
    InMux I__1452 (
            .O(N__16990),
            .I(N__16984));
    LocalMux I__1451 (
            .O(N__16987),
            .I(secclk_cnt_7));
    LocalMux I__1450 (
            .O(N__16984),
            .I(secclk_cnt_7));
    InMux I__1449 (
            .O(N__16979),
            .I(n14015));
    InMux I__1448 (
            .O(N__16976),
            .I(N__16972));
    InMux I__1447 (
            .O(N__16975),
            .I(N__16969));
    LocalMux I__1446 (
            .O(N__16972),
            .I(secclk_cnt_8));
    LocalMux I__1445 (
            .O(N__16969),
            .I(secclk_cnt_8));
    InMux I__1444 (
            .O(N__16964),
            .I(bfn_3_8_0_));
    InMux I__1443 (
            .O(N__16961),
            .I(N__16957));
    InMux I__1442 (
            .O(N__16960),
            .I(N__16954));
    LocalMux I__1441 (
            .O(N__16957),
            .I(secclk_cnt_9));
    LocalMux I__1440 (
            .O(N__16954),
            .I(secclk_cnt_9));
    InMux I__1439 (
            .O(N__16949),
            .I(n14017));
    CascadeMux I__1438 (
            .O(N__16946),
            .I(N__16942));
    InMux I__1437 (
            .O(N__16945),
            .I(N__16939));
    InMux I__1436 (
            .O(N__16942),
            .I(N__16936));
    LocalMux I__1435 (
            .O(N__16939),
            .I(secclk_cnt_10));
    LocalMux I__1434 (
            .O(N__16936),
            .I(secclk_cnt_10));
    InMux I__1433 (
            .O(N__16931),
            .I(n14018));
    CascadeMux I__1432 (
            .O(N__16928),
            .I(N__16924));
    InMux I__1431 (
            .O(N__16927),
            .I(N__16921));
    InMux I__1430 (
            .O(N__16924),
            .I(N__16918));
    LocalMux I__1429 (
            .O(N__16921),
            .I(secclk_cnt_11));
    LocalMux I__1428 (
            .O(N__16918),
            .I(secclk_cnt_11));
    InMux I__1427 (
            .O(N__16913),
            .I(n14019));
    InMux I__1426 (
            .O(N__16910),
            .I(n14020));
    InMux I__1425 (
            .O(N__16907),
            .I(N__16904));
    LocalMux I__1424 (
            .O(N__16904),
            .I(n28));
    InMux I__1423 (
            .O(N__16901),
            .I(N__16898));
    LocalMux I__1422 (
            .O(N__16898),
            .I(n26_adj_1180));
    InMux I__1421 (
            .O(N__16895),
            .I(N__16892));
    LocalMux I__1420 (
            .O(N__16892),
            .I(n10));
    IoInMux I__1419 (
            .O(N__16889),
            .I(N__16886));
    LocalMux I__1418 (
            .O(N__16886),
            .I(N__16883));
    Span4Mux_s2_v I__1417 (
            .O(N__16883),
            .I(N__16880));
    Span4Mux_v I__1416 (
            .O(N__16880),
            .I(N__16877));
    Odrv4 I__1415 (
            .O(N__16877),
            .I(DDS_MCLK1));
    InMux I__1414 (
            .O(N__16874),
            .I(N__16870));
    InMux I__1413 (
            .O(N__16873),
            .I(N__16867));
    LocalMux I__1412 (
            .O(N__16870),
            .I(secclk_cnt_0));
    LocalMux I__1411 (
            .O(N__16867),
            .I(secclk_cnt_0));
    InMux I__1410 (
            .O(N__16862),
            .I(bfn_3_7_0_));
    CascadeMux I__1409 (
            .O(N__16859),
            .I(N__16855));
    InMux I__1408 (
            .O(N__16858),
            .I(N__16852));
    InMux I__1407 (
            .O(N__16855),
            .I(N__16849));
    LocalMux I__1406 (
            .O(N__16852),
            .I(secclk_cnt_1));
    LocalMux I__1405 (
            .O(N__16849),
            .I(secclk_cnt_1));
    InMux I__1404 (
            .O(N__16844),
            .I(n14009));
    InMux I__1403 (
            .O(N__16841),
            .I(N__16837));
    InMux I__1402 (
            .O(N__16840),
            .I(N__16834));
    LocalMux I__1401 (
            .O(N__16837),
            .I(secclk_cnt_2));
    LocalMux I__1400 (
            .O(N__16834),
            .I(secclk_cnt_2));
    InMux I__1399 (
            .O(N__16829),
            .I(n14010));
    InMux I__1398 (
            .O(N__16826),
            .I(N__16822));
    InMux I__1397 (
            .O(N__16825),
            .I(N__16819));
    LocalMux I__1396 (
            .O(N__16822),
            .I(secclk_cnt_3));
    LocalMux I__1395 (
            .O(N__16819),
            .I(secclk_cnt_3));
    InMux I__1394 (
            .O(N__16814),
            .I(n14011));
    CascadeMux I__1393 (
            .O(N__16811),
            .I(n25_cascade_));
    InMux I__1392 (
            .O(N__16808),
            .I(N__16805));
    LocalMux I__1391 (
            .O(N__16805),
            .I(n27_adj_1173));
    CascadeMux I__1390 (
            .O(N__16802),
            .I(n14114_cascade_));
    CascadeMux I__1389 (
            .O(N__16799),
            .I(n10522_cascade_));
    IoInMux I__1388 (
            .O(N__16796),
            .I(N__16793));
    LocalMux I__1387 (
            .O(N__16793),
            .I(N__16790));
    IoSpan4Mux I__1386 (
            .O(N__16790),
            .I(N__16787));
    Span4Mux_s1_v I__1385 (
            .O(N__16787),
            .I(N__16784));
    Sp12to4 I__1384 (
            .O(N__16784),
            .I(N__16781));
    Span12Mux_v I__1383 (
            .O(N__16781),
            .I(N__16777));
    InMux I__1382 (
            .O(N__16780),
            .I(N__16774));
    Odrv12 I__1381 (
            .O(N__16777),
            .I(TEST_LED));
    LocalMux I__1380 (
            .O(N__16774),
            .I(TEST_LED));
    IoInMux I__1379 (
            .O(N__16769),
            .I(N__16766));
    LocalMux I__1378 (
            .O(N__16766),
            .I(N__16763));
    IoSpan4Mux I__1377 (
            .O(N__16763),
            .I(N__16760));
    IoSpan4Mux I__1376 (
            .O(N__16760),
            .I(N__16757));
    Odrv4 I__1375 (
            .O(N__16757),
            .I(ICE_SYSCLK));
    IoInMux I__1374 (
            .O(N__16754),
            .I(N__16750));
    IoInMux I__1373 (
            .O(N__16753),
            .I(N__16746));
    LocalMux I__1372 (
            .O(N__16750),
            .I(N__16742));
    IoInMux I__1371 (
            .O(N__16749),
            .I(N__16739));
    LocalMux I__1370 (
            .O(N__16746),
            .I(N__16736));
    IoInMux I__1369 (
            .O(N__16745),
            .I(N__16733));
    IoSpan4Mux I__1368 (
            .O(N__16742),
            .I(N__16730));
    LocalMux I__1367 (
            .O(N__16739),
            .I(N__16727));
    IoSpan4Mux I__1366 (
            .O(N__16736),
            .I(N__16722));
    LocalMux I__1365 (
            .O(N__16733),
            .I(N__16722));
    Span4Mux_s1_v I__1364 (
            .O(N__16730),
            .I(N__16719));
    Span4Mux_s1_v I__1363 (
            .O(N__16727),
            .I(N__16716));
    IoSpan4Mux I__1362 (
            .O(N__16722),
            .I(N__16713));
    Sp12to4 I__1361 (
            .O(N__16719),
            .I(N__16710));
    Sp12to4 I__1360 (
            .O(N__16716),
            .I(N__16707));
    Span4Mux_s2_h I__1359 (
            .O(N__16713),
            .I(N__16704));
    Span12Mux_s9_v I__1358 (
            .O(N__16710),
            .I(N__16701));
    Span12Mux_h I__1357 (
            .O(N__16707),
            .I(N__16698));
    Sp12to4 I__1356 (
            .O(N__16704),
            .I(N__16695));
    Span12Mux_v I__1355 (
            .O(N__16701),
            .I(N__16692));
    Span12Mux_v I__1354 (
            .O(N__16698),
            .I(N__16689));
    Span12Mux_v I__1353 (
            .O(N__16695),
            .I(N__16686));
    Span12Mux_h I__1352 (
            .O(N__16692),
            .I(N__16683));
    Span12Mux_v I__1351 (
            .O(N__16689),
            .I(N__16678));
    Span12Mux_h I__1350 (
            .O(N__16686),
            .I(N__16678));
    Odrv12 I__1349 (
            .O(N__16683),
            .I(M_CLK4));
    Odrv12 I__1348 (
            .O(N__16678),
            .I(M_CLK4));
    IoInMux I__1347 (
            .O(N__16673),
            .I(N__16670));
    LocalMux I__1346 (
            .O(N__16670),
            .I(N__16667));
    IoSpan4Mux I__1345 (
            .O(N__16667),
            .I(N__16664));
    Sp12to4 I__1344 (
            .O(N__16664),
            .I(N__16661));
    Span12Mux_s3_v I__1343 (
            .O(N__16661),
            .I(N__16658));
    Span12Mux_h I__1342 (
            .O(N__16658),
            .I(N__16655));
    Odrv12 I__1341 (
            .O(N__16655),
            .I(ICE_GPMO_2));
    INV \INVcomm_spi.bit_cnt_1603__i3C  (
            .O(\INVcomm_spi.bit_cnt_1603__i3C_net ),
            .I(N__42424));
    INV INVdata_count_i0_i8C (
            .O(INVdata_count_i0_i8C_net),
            .I(N__51309));
    INV INVdata_count_i0_i0C (
            .O(INVdata_count_i0_i0C_net),
            .I(N__51303));
    INV INVdata_cntvec_i0_i8C (
            .O(INVdata_cntvec_i0_i8C_net),
            .I(N__51294));
    INV INVdata_cntvec_i0_i0C (
            .O(INVdata_cntvec_i0_i0C_net),
            .I(N__51283));
    INV \INVcomm_spi.MISO_48_7334_7335_setC  (
            .O(\INVcomm_spi.MISO_48_7334_7335_setC_net ),
            .I(N__51131));
    INV \INVcomm_spi.MISO_48_7334_7335_resetC  (
            .O(\INVcomm_spi.MISO_48_7334_7335_resetC_net ),
            .I(N__51116));
    INV INVacadc_trig_329C (
            .O(INVacadc_trig_329C_net),
            .I(N__51281));
    INV \INVcomm_spi.imiso_83_7340_7341_setC  (
            .O(\INVcomm_spi.imiso_83_7340_7341_setC_net ),
            .I(N__42420));
    INV \INVcomm_spi.data_valid_85C  (
            .O(\INVcomm_spi.data_valid_85C_net ),
            .I(N__51123));
    INV INVacadc_skipcnt_i0_i9C (
            .O(INVacadc_skipcnt_i0_i9C_net),
            .I(N__51268));
    INV INVacadc_skipcnt_i0_i1C (
            .O(INVacadc_skipcnt_i0_i1C_net),
            .I(N__51252));
    INV INVacadc_skipcnt_i0_i0C (
            .O(INVacadc_skipcnt_i0_i0C_net),
            .I(N__51236));
    INV INVeis_state_i0C (
            .O(INVeis_state_i0C_net),
            .I(N__51184));
    INV INVeis_end_328C (
            .O(INVeis_end_328C_net),
            .I(N__51166));
    INV \INVcomm_spi.imiso_83_7340_7341_resetC  (
            .O(\INVcomm_spi.imiso_83_7340_7341_resetC_net ),
            .I(N__42440));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN_net),
            .I(N__51260));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN_net),
            .I(N__51288));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN_net),
            .I(N__51175));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN_net),
            .I(N__51306));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN_net),
            .I(N__51210));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN_net),
            .I(N__51227));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN_net),
            .I(N__51314));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN_net),
            .I(N__51135));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN_net),
            .I(N__51193));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN_net),
            .I(N__51318));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN_net),
            .I(N__51157));
    INV INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN (
            .O(INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN_net),
            .I(N__51320));
    defparam IN_MUX_bfv_3_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_7_0_));
    defparam IN_MUX_bfv_3_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_8_0_ (
            .carryinitin(n14016),
            .carryinitout(bfn_3_8_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(n14024),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(n13966_THRU_CRY_6_THRU_CO),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(n13974),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(n13958),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(n13949),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(n14038),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(n14047),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_6_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_16_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam i11_4_lut_adj_191_LC_2_7_3.C_ON=1'b0;
    defparam i11_4_lut_adj_191_LC_2_7_3.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_191_LC_2_7_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_191_LC_2_7_3 (
            .in0(N__17005),
            .in1(N__17131),
            .in2(N__16946),
            .in3(N__16825),
            .lcout(n27_adj_1173),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_2_8_0.C_ON=1'b0;
    defparam i9_4_lut_LC_2_8_0.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_2_8_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_2_8_0 (
            .in0(N__17116),
            .in1(N__16975),
            .in2(N__16859),
            .in3(N__17020),
            .lcout(),
            .ltout(n25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_193_LC_2_8_1.C_ON=1'b0;
    defparam i15_4_lut_adj_193_LC_2_8_1.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_193_LC_2_8_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_193_LC_2_8_1 (
            .in0(N__16907),
            .in1(N__16901),
            .in2(N__16811),
            .in3(N__16808),
            .lcout(),
            .ltout(n14114_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_194_LC_2_8_2.C_ON=1'b0;
    defparam i7_4_lut_adj_194_LC_2_8_2.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_194_LC_2_8_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 i7_4_lut_adj_194_LC_2_8_2 (
            .in0(N__17050),
            .in1(N__16895),
            .in2(N__16802),
            .in3(N__18518),
            .lcout(n10522),
            .ltout(n10522_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SecClk_321_LC_2_8_3.C_ON=1'b0;
    defparam SecClk_321_LC_2_8_3.SEQ_MODE=4'b1000;
    defparam SecClk_321_LC_2_8_3.LUT_INIT=16'b0101101001011010;
    LogicCell40 SecClk_321_LC_2_8_3 (
            .in0(N__16780),
            .in1(_gnd_net_),
            .in2(N__16799),
            .in3(_gnd_net_),
            .lcout(TEST_LED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17277),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_189_LC_2_8_4.C_ON=1'b0;
    defparam i12_4_lut_adj_189_LC_2_8_4.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_189_LC_2_8_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_189_LC_2_8_4 (
            .in0(N__17068),
            .in1(N__16873),
            .in2(N__16928),
            .in3(N__17035),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_190_LC_2_8_5.C_ON=1'b0;
    defparam i10_4_lut_adj_190_LC_2_8_5.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_190_LC_2_8_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_190_LC_2_8_5 (
            .in0(N__17102),
            .in1(N__16990),
            .in2(N__17153),
            .in3(N__16840),
            .lcout(n26_adj_1180),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_2_9_1.C_ON=1'b0;
    defparam i2_2_lut_LC_2_9_1.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_2_9_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2_2_lut_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(N__16960),
            .in2(_gnd_net_),
            .in3(N__17083),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_58_LC_2_14_2.C_ON=1'b0;
    defparam i1_2_lut_adj_58_LC_2_14_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_58_LC_2_14_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_58_LC_2_14_2 (
            .in0(_gnd_net_),
            .in1(N__36410),
            .in2(_gnd_net_),
            .in3(N__35617),
            .lcout(n15165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_16MHz_I_0_1_lut_LC_3_1_2.C_ON=1'b0;
    defparam clk_16MHz_I_0_1_lut_LC_3_1_2.SEQ_MODE=4'b0000;
    defparam clk_16MHz_I_0_1_lut_LC_3_1_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 clk_16MHz_I_0_1_lut_LC_3_1_2 (
            .in0(N__17282),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DDS_MCLK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secclk_cnt_1601_1602__i1_LC_3_7_0.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i1_LC_3_7_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i1_LC_3_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i1_LC_3_7_0 (
            .in0(_gnd_net_),
            .in1(N__16874),
            .in2(_gnd_net_),
            .in3(N__16862),
            .lcout(secclk_cnt_0),
            .ltout(),
            .carryin(bfn_3_7_0_),
            .carryout(n14009),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i2_LC_3_7_1.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i2_LC_3_7_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i2_LC_3_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i2_LC_3_7_1 (
            .in0(_gnd_net_),
            .in1(N__16858),
            .in2(_gnd_net_),
            .in3(N__16844),
            .lcout(secclk_cnt_1),
            .ltout(),
            .carryin(n14009),
            .carryout(n14010),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i3_LC_3_7_2.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i3_LC_3_7_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i3_LC_3_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i3_LC_3_7_2 (
            .in0(_gnd_net_),
            .in1(N__16841),
            .in2(_gnd_net_),
            .in3(N__16829),
            .lcout(secclk_cnt_2),
            .ltout(),
            .carryin(n14010),
            .carryout(n14011),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i4_LC_3_7_3.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i4_LC_3_7_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i4_LC_3_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i4_LC_3_7_3 (
            .in0(_gnd_net_),
            .in1(N__16826),
            .in2(_gnd_net_),
            .in3(N__16814),
            .lcout(secclk_cnt_3),
            .ltout(),
            .carryin(n14011),
            .carryout(n14012),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i5_LC_3_7_4.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i5_LC_3_7_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i5_LC_3_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i5_LC_3_7_4 (
            .in0(_gnd_net_),
            .in1(N__17036),
            .in2(_gnd_net_),
            .in3(N__17024),
            .lcout(secclk_cnt_4),
            .ltout(),
            .carryin(n14012),
            .carryout(n14013),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i6_LC_3_7_5.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i6_LC_3_7_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i6_LC_3_7_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i6_LC_3_7_5 (
            .in0(_gnd_net_),
            .in1(N__17021),
            .in2(_gnd_net_),
            .in3(N__17009),
            .lcout(secclk_cnt_5),
            .ltout(),
            .carryin(n14013),
            .carryout(n14014),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i7_LC_3_7_6.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i7_LC_3_7_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i7_LC_3_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i7_LC_3_7_6 (
            .in0(_gnd_net_),
            .in1(N__17006),
            .in2(_gnd_net_),
            .in3(N__16994),
            .lcout(secclk_cnt_6),
            .ltout(),
            .carryin(n14014),
            .carryout(n14015),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i8_LC_3_7_7.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i8_LC_3_7_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i8_LC_3_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i8_LC_3_7_7 (
            .in0(_gnd_net_),
            .in1(N__16991),
            .in2(_gnd_net_),
            .in3(N__16979),
            .lcout(secclk_cnt_7),
            .ltout(),
            .carryin(n14015),
            .carryout(n14016),
            .clk(N__17275),
            .ce(),
            .sr(N__17257));
    defparam secclk_cnt_1601_1602__i9_LC_3_8_0.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i9_LC_3_8_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i9_LC_3_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i9_LC_3_8_0 (
            .in0(_gnd_net_),
            .in1(N__16976),
            .in2(_gnd_net_),
            .in3(N__16964),
            .lcout(secclk_cnt_8),
            .ltout(),
            .carryin(bfn_3_8_0_),
            .carryout(n14017),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i10_LC_3_8_1.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i10_LC_3_8_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i10_LC_3_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i10_LC_3_8_1 (
            .in0(_gnd_net_),
            .in1(N__16961),
            .in2(_gnd_net_),
            .in3(N__16949),
            .lcout(secclk_cnt_9),
            .ltout(),
            .carryin(n14017),
            .carryout(n14018),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i11_LC_3_8_2.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i11_LC_3_8_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i11_LC_3_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i11_LC_3_8_2 (
            .in0(_gnd_net_),
            .in1(N__16945),
            .in2(_gnd_net_),
            .in3(N__16931),
            .lcout(secclk_cnt_10),
            .ltout(),
            .carryin(n14018),
            .carryout(n14019),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i12_LC_3_8_3.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i12_LC_3_8_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i12_LC_3_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i12_LC_3_8_3 (
            .in0(_gnd_net_),
            .in1(N__16927),
            .in2(_gnd_net_),
            .in3(N__16913),
            .lcout(secclk_cnt_11),
            .ltout(),
            .carryin(n14019),
            .carryout(n14020),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i13_LC_3_8_4.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i13_LC_3_8_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i13_LC_3_8_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i13_LC_3_8_4 (
            .in0(_gnd_net_),
            .in1(N__18547),
            .in2(_gnd_net_),
            .in3(N__16910),
            .lcout(secclk_cnt_12),
            .ltout(),
            .carryin(n14020),
            .carryout(n14021),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i14_LC_3_8_5.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i14_LC_3_8_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i14_LC_3_8_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i14_LC_3_8_5 (
            .in0(_gnd_net_),
            .in1(N__17149),
            .in2(_gnd_net_),
            .in3(N__17135),
            .lcout(secclk_cnt_13),
            .ltout(),
            .carryin(n14021),
            .carryout(n14022),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i15_LC_3_8_6.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i15_LC_3_8_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i15_LC_3_8_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i15_LC_3_8_6 (
            .in0(_gnd_net_),
            .in1(N__17132),
            .in2(_gnd_net_),
            .in3(N__17120),
            .lcout(secclk_cnt_14),
            .ltout(),
            .carryin(n14022),
            .carryout(n14023),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i16_LC_3_8_7.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i16_LC_3_8_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i16_LC_3_8_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i16_LC_3_8_7 (
            .in0(_gnd_net_),
            .in1(N__17117),
            .in2(_gnd_net_),
            .in3(N__17105),
            .lcout(secclk_cnt_15),
            .ltout(),
            .carryin(n14023),
            .carryout(n14024),
            .clk(N__17276),
            .ce(),
            .sr(N__17250));
    defparam secclk_cnt_1601_1602__i17_LC_3_9_0.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i17_LC_3_9_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i17_LC_3_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i17_LC_3_9_0 (
            .in0(_gnd_net_),
            .in1(N__17101),
            .in2(_gnd_net_),
            .in3(N__17087),
            .lcout(secclk_cnt_16),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(n14025),
            .clk(N__17278),
            .ce(),
            .sr(N__17258));
    defparam secclk_cnt_1601_1602__i18_LC_3_9_1.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i18_LC_3_9_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i18_LC_3_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i18_LC_3_9_1 (
            .in0(_gnd_net_),
            .in1(N__17084),
            .in2(_gnd_net_),
            .in3(N__17072),
            .lcout(secclk_cnt_17),
            .ltout(),
            .carryin(n14025),
            .carryout(n14026),
            .clk(N__17278),
            .ce(),
            .sr(N__17258));
    defparam secclk_cnt_1601_1602__i19_LC_3_9_2.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i19_LC_3_9_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i19_LC_3_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i19_LC_3_9_2 (
            .in0(_gnd_net_),
            .in1(N__17069),
            .in2(_gnd_net_),
            .in3(N__17057),
            .lcout(secclk_cnt_18),
            .ltout(),
            .carryin(n14026),
            .carryout(n14027),
            .clk(N__17278),
            .ce(),
            .sr(N__17258));
    defparam secclk_cnt_1601_1602__i20_LC_3_9_3.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i20_LC_3_9_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i20_LC_3_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i20_LC_3_9_3 (
            .in0(_gnd_net_),
            .in1(N__18568),
            .in2(_gnd_net_),
            .in3(N__17054),
            .lcout(secclk_cnt_19),
            .ltout(),
            .carryin(n14027),
            .carryout(n14028),
            .clk(N__17278),
            .ce(),
            .sr(N__17258));
    defparam secclk_cnt_1601_1602__i21_LC_3_9_4.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i21_LC_3_9_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i21_LC_3_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i21_LC_3_9_4 (
            .in0(_gnd_net_),
            .in1(N__17051),
            .in2(_gnd_net_),
            .in3(N__17039),
            .lcout(secclk_cnt_20),
            .ltout(),
            .carryin(n14028),
            .carryout(n14029),
            .clk(N__17278),
            .ce(),
            .sr(N__17258));
    defparam secclk_cnt_1601_1602__i22_LC_3_9_5.C_ON=1'b1;
    defparam secclk_cnt_1601_1602__i22_LC_3_9_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i22_LC_3_9_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i22_LC_3_9_5 (
            .in0(_gnd_net_),
            .in1(N__18583),
            .in2(_gnd_net_),
            .in3(N__17288),
            .lcout(secclk_cnt_21),
            .ltout(),
            .carryin(n14029),
            .carryout(n14030),
            .clk(N__17278),
            .ce(),
            .sr(N__17258));
    defparam secclk_cnt_1601_1602__i23_LC_3_9_6.C_ON=1'b0;
    defparam secclk_cnt_1601_1602__i23_LC_3_9_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_1601_1602__i23_LC_3_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_1601_1602__i23_LC_3_9_6 (
            .in0(_gnd_net_),
            .in1(N__18532),
            .in2(_gnd_net_),
            .in3(N__17285),
            .lcout(secclk_cnt_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17278),
            .ce(),
            .sr(N__17258));
    defparam \ADC_VAC2.ADC_DATA_i0_LC_3_10_0 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i0_LC_3_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i0_LC_3_10_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i0_LC_3_10_0  (
            .in0(N__53685),
            .in1(N__53436),
            .in2(N__17215),
            .in3(N__17195),
            .lcout(buf_adcdata2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i9_LC_3_10_2 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i9_LC_3_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i9_LC_3_10_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i9_LC_3_10_2  (
            .in0(N__46004),
            .in1(N__53437),
            .in2(N__42931),
            .in3(N__17194),
            .lcout(cmd_rdadctmp_9_adj_1067),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i8_LC_3_10_4 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i8_LC_3_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i8_LC_3_10_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i8_LC_3_10_4  (
            .in0(N__46003),
            .in1(N__17193),
            .in2(N__17183),
            .in3(N__53438),
            .lcout(cmd_rdadctmp_8_adj_1068),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i7_LC_3_10_5 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i7_LC_3_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i7_LC_3_10_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i7_LC_3_10_5  (
            .in0(N__53435),
            .in1(N__17179),
            .in2(N__17171),
            .in3(N__46002),
            .lcout(cmd_rdadctmp_7_adj_1069),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51275),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i10_LC_3_10_7 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i10_LC_3_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i10_LC_3_10_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i10_LC_3_10_7  (
            .in0(N__53434),
            .in1(N__42927),
            .in2(N__46696),
            .in3(N__46001),
            .lcout(cmd_rdadctmp_10_adj_1066),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51275),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_17_LC_3_12_2.C_ON=1'b0;
    defparam i1_2_lut_adj_17_LC_3_12_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_17_LC_3_12_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_17_LC_3_12_2 (
            .in0(_gnd_net_),
            .in1(N__36449),
            .in2(_gnd_net_),
            .in3(N__35616),
            .lcout(n15150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i6_LC_3_13_0 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i6_LC_3_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i6_LC_3_13_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i6_LC_3_13_0  (
            .in0(N__53391),
            .in1(N__17164),
            .in2(N__46038),
            .in3(N__17422),
            .lcout(cmd_rdadctmp_6_adj_1070),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51307),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i3_LC_3_13_1 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i3_LC_3_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i3_LC_3_13_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i3_LC_3_13_1  (
            .in0(N__17327),
            .in1(N__45993),
            .in2(N__17411),
            .in3(N__53392),
            .lcout(cmd_rdadctmp_3_adj_1073),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51307),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i5_LC_3_13_3 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i5_LC_3_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i5_LC_3_13_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i5_LC_3_13_3  (
            .in0(N__17399),
            .in1(N__45997),
            .in2(N__17423),
            .in3(N__53393),
            .lcout(cmd_rdadctmp_5_adj_1071),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51307),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i4_LC_3_13_4 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i4_LC_3_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i4_LC_3_13_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i4_LC_3_13_4  (
            .in0(N__53390),
            .in1(N__17410),
            .in2(N__46037),
            .in3(N__17398),
            .lcout(cmd_rdadctmp_4_adj_1072),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51307),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.adc_state_i2_LC_3_14_0 .C_ON=1'b0;
    defparam \ADC_VAC2.adc_state_i2_LC_3_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.adc_state_i2_LC_3_14_0 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \ADC_VAC2.adc_state_i2_LC_3_14_0  (
            .in0(N__36429),
            .in1(N__53335),
            .in2(_gnd_net_),
            .in3(N__35618),
            .lcout(DTRIG_N_957_adj_1077),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51311),
            .ce(N__35503),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_207_LC_3_15_1.C_ON=1'b0;
    defparam i1_4_lut_adj_207_LC_3_15_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_207_LC_3_15_1.LUT_INIT=16'b0000111100000110;
    LogicCell40 i1_4_lut_adj_207_LC_3_15_1 (
            .in0(N__36428),
            .in1(N__53404),
            .in2(N__17377),
            .in3(N__35608),
            .lcout(),
            .ltout(n14_adj_1035_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.CS_37_LC_3_15_2 .C_ON=1'b0;
    defparam \ADC_VAC2.CS_37_LC_3_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.CS_37_LC_3_15_2 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \ADC_VAC2.CS_37_LC_3_15_2  (
            .in0(N__53405),
            .in1(N__30185),
            .in2(N__17390),
            .in3(N__17360),
            .lcout(M_CS2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51315),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i1_3_lut_adj_4_LC_3_15_3 .C_ON=1'b0;
    defparam \ADC_VAC2.i1_3_lut_adj_4_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i1_3_lut_adj_4_LC_3_15_3 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \ADC_VAC2.i1_3_lut_adj_4_LC_3_15_3  (
            .in0(N__30186),
            .in1(N__17359),
            .in2(_gnd_net_),
            .in3(N__53403),
            .lcout(n8302),
            .ltout(n8302_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i0_LC_3_15_4 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i0_LC_3_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i0_LC_3_15_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i0_LC_3_15_4  (
            .in0(N__53406),
            .in1(N__17348),
            .in2(N__17330),
            .in3(N__17308),
            .lcout(cmd_rdadctmp_0_adj_1076),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51315),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i2_LC_3_15_5 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i2_LC_3_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i2_LC_3_15_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i2_LC_3_15_5  (
            .in0(N__45949),
            .in1(N__17299),
            .in2(N__17326),
            .in3(N__53408),
            .lcout(cmd_rdadctmp_2_adj_1074),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51315),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i1_LC_3_15_6 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i1_LC_3_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i1_LC_3_15_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i1_LC_3_15_6  (
            .in0(N__53407),
            .in1(N__17309),
            .in2(N__17300),
            .in3(N__45948),
            .lcout(cmd_rdadctmp_1_adj_1075),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51315),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i7_LC_5_5_3 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i7_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i7_LC_5_5_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i7_LC_5_5_3  (
            .in0(N__27527),
            .in1(N__18059),
            .in2(N__25967),
            .in3(N__17473),
            .lcout(buf_adcdata4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51159),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1525_i7_4_lut_LC_5_5_4.C_ON=1'b0;
    defparam mux_1525_i7_4_lut_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam mux_1525_i7_4_lut_LC_5_5_4.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1525_i7_4_lut_LC_5_5_4 (
            .in0(N__17480),
            .in1(N__48060),
            .in2(N__17687),
            .in3(N__47339),
            .lcout(n4302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i3_LC_5_5_6 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i3_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i3_LC_5_5_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_VAC4.ADC_DATA_i3_LC_5_5_6  (
            .in0(N__20811),
            .in1(N__25962),
            .in2(N__18233),
            .in3(N__27528),
            .lcout(buf_adcdata4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51159),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1525_i8_4_lut_LC_5_5_7.C_ON=1'b0;
    defparam mux_1525_i8_4_lut_LC_5_5_7.SEQ_MODE=4'b0000;
    defparam mux_1525_i8_4_lut_LC_5_5_7.LUT_INIT=16'b1010111000000100;
    LogicCell40 mux_1525_i8_4_lut_LC_5_5_7 (
            .in0(N__47338),
            .in1(N__17472),
            .in2(N__48085),
            .in3(N__17459),
            .lcout(n4301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1525_i5_4_lut_LC_5_6_0.C_ON=1'b0;
    defparam mux_1525_i5_4_lut_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam mux_1525_i5_4_lut_LC_5_6_0.LUT_INIT=16'b1111000001000100;
    LogicCell40 mux_1525_i5_4_lut_LC_5_6_0 (
            .in0(N__48072),
            .in1(N__18120),
            .in2(N__17453),
            .in3(N__47322),
            .lcout(),
            .ltout(n4304_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_5__i4_LC_5_6_1.C_ON=1'b0;
    defparam comm_buf_5__i4_LC_5_6_1.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i4_LC_5_6_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_5__i4_LC_5_6_1 (
            .in0(_gnd_net_),
            .in1(N__39903),
            .in2(N__17441),
            .in3(N__50274),
            .lcout(comm_buf_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51176),
            .ce(N__18325),
            .sr(N__18298));
    defparam mux_1525_i6_4_lut_LC_5_6_2.C_ON=1'b0;
    defparam mux_1525_i6_4_lut_LC_5_6_2.SEQ_MODE=4'b0000;
    defparam mux_1525_i6_4_lut_LC_5_6_2.LUT_INIT=16'b1100110001010000;
    LogicCell40 mux_1525_i6_4_lut_LC_5_6_2 (
            .in0(N__48073),
            .in1(N__17438),
            .in2(N__17756),
            .in3(N__47323),
            .lcout(),
            .ltout(n4303_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_5__i5_LC_5_6_3.C_ON=1'b0;
    defparam comm_buf_5__i5_LC_5_6_3.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i5_LC_5_6_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_5__i5_LC_5_6_3 (
            .in0(_gnd_net_),
            .in1(N__39797),
            .in2(N__17432),
            .in3(N__50275),
            .lcout(comm_buf_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51176),
            .ce(N__18325),
            .sr(N__18298));
    defparam comm_buf_5__i6_LC_5_6_5.C_ON=1'b0;
    defparam comm_buf_5__i6_LC_5_6_5.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i6_LC_5_6_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i6_LC_5_6_5 (
            .in0(N__40693),
            .in1(N__17429),
            .in2(_gnd_net_),
            .in3(N__50276),
            .lcout(comm_buf_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51176),
            .ce(N__18325),
            .sr(N__18298));
    defparam comm_buf_5__i7_LC_5_6_7.C_ON=1'b0;
    defparam comm_buf_5__i7_LC_5_6_7.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i7_LC_5_6_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i7_LC_5_6_7 (
            .in0(N__39338),
            .in1(N__17552),
            .in2(_gnd_net_),
            .in3(N__50277),
            .lcout(comm_buf_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51176),
            .ce(N__18325),
            .sr(N__18298));
    defparam comm_buf_2__i6_LC_5_7_1.C_ON=1'b0;
    defparam comm_buf_2__i6_LC_5_7_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i6_LC_5_7_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i6_LC_5_7_1 (
            .in0(N__40739),
            .in1(N__18089),
            .in2(_gnd_net_),
            .in3(N__50340),
            .lcout(comm_buf_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51194),
            .ce(N__18377),
            .sr(N__18613));
    defparam comm_buf_2__i7_LC_5_7_3.C_ON=1'b0;
    defparam comm_buf_2__i7_LC_5_7_3.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i7_LC_5_7_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_2__i7_LC_5_7_3 (
            .in0(N__18350),
            .in1(N__39397),
            .in2(_gnd_net_),
            .in3(N__50341),
            .lcout(comm_buf_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51194),
            .ce(N__18377),
            .sr(N__18613));
    defparam mux_1525_i1_4_lut_LC_5_7_4.C_ON=1'b0;
    defparam mux_1525_i1_4_lut_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam mux_1525_i1_4_lut_LC_5_7_4.LUT_INIT=16'b1000101110001000;
    LogicCell40 mux_1525_i1_4_lut_LC_5_7_4 (
            .in0(N__17546),
            .in1(N__47230),
            .in2(N__48086),
            .in3(N__18016),
            .lcout(n4308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1525_i2_4_lut_LC_5_7_5.C_ON=1'b0;
    defparam mux_1525_i2_4_lut_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam mux_1525_i2_4_lut_LC_5_7_5.LUT_INIT=16'b1011101000010000;
    LogicCell40 mux_1525_i2_4_lut_LC_5_7_5 (
            .in0(N__47231),
            .in1(N__48067),
            .in2(N__17986),
            .in3(N__17528),
            .lcout(n4307),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1525_i3_4_lut_LC_5_7_6.C_ON=1'b0;
    defparam mux_1525_i3_4_lut_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam mux_1525_i3_4_lut_LC_5_7_6.LUT_INIT=16'b1010000010101100;
    LogicCell40 mux_1525_i3_4_lut_LC_5_7_6 (
            .in0(N__17516),
            .in1(N__17914),
            .in2(N__47336),
            .in3(N__48068),
            .lcout(n4306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_5__i1_LC_5_8_0.C_ON=1'b0;
    defparam comm_buf_5__i1_LC_5_8_0.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i1_LC_5_8_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i1_LC_5_8_0 (
            .in0(N__44180),
            .in1(N__17498),
            .in2(_gnd_net_),
            .in3(N__50273),
            .lcout(comm_buf_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51211),
            .ce(N__18329),
            .sr(N__18299));
    defparam comm_buf_5__i2_LC_5_8_1.C_ON=1'b0;
    defparam comm_buf_5__i2_LC_5_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i2_LC_5_8_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i2_LC_5_8_1 (
            .in0(N__50270),
            .in1(N__40124),
            .in2(_gnd_net_),
            .in3(N__17492),
            .lcout(comm_buf_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51211),
            .ce(N__18329),
            .sr(N__18299));
    defparam comm_buf_5__i0_LC_5_8_2.C_ON=1'b0;
    defparam comm_buf_5__i0_LC_5_8_2.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i0_LC_5_8_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_5__i0_LC_5_8_2 (
            .in0(N__17486),
            .in1(N__50272),
            .in2(_gnd_net_),
            .in3(N__39215),
            .lcout(comm_buf_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51211),
            .ce(N__18329),
            .sr(N__18299));
    defparam comm_buf_5__i3_LC_5_8_3.C_ON=1'b0;
    defparam comm_buf_5__i3_LC_5_8_3.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i3_LC_5_8_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i3_LC_5_8_3 (
            .in0(N__50271),
            .in1(N__44921),
            .in2(_gnd_net_),
            .in3(N__20792),
            .lcout(comm_buf_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51211),
            .ce(N__18329),
            .sr(N__18299));
    defparam \ADC_VAC2.ADC_DATA_i5_LC_5_9_0 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i5_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i5_LC_5_9_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i5_LC_5_9_0  (
            .in0(N__53702),
            .in1(N__17653),
            .in2(N__17870),
            .in3(N__53518),
            .lcout(buf_adcdata2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51228),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i6_LC_5_9_1 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i6_LC_5_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i6_LC_5_9_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i6_LC_5_9_1  (
            .in0(N__53515),
            .in1(N__53704),
            .in2(N__17638),
            .in3(N__17846),
            .lcout(buf_adcdata2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51228),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i7_LC_5_9_2 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i7_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i7_LC_5_9_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i7_LC_5_9_2  (
            .in0(N__53703),
            .in1(N__53517),
            .in2(N__17617),
            .in3(N__17596),
            .lcout(buf_adcdata2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51228),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i15_LC_5_9_3 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i15_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i15_LC_5_9_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i15_LC_5_9_3  (
            .in0(N__53516),
            .in1(N__17845),
            .in2(N__17597),
            .in3(N__46079),
            .lcout(cmd_rdadctmp_15_adj_1061),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51228),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i16_LC_5_9_4 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i16_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i16_LC_5_9_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i16_LC_5_9_4  (
            .in0(N__46080),
            .in1(N__17595),
            .in2(N__20445),
            .in3(N__53519),
            .lcout(cmd_rdadctmp_16_adj_1060),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51228),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i3_LC_5_10_2 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i3_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i3_LC_5_10_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i3_LC_5_10_2  (
            .in0(N__53695),
            .in1(N__53523),
            .in2(N__17572),
            .in3(N__17829),
            .lcout(buf_adcdata2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51244),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i11_LC_5_10_3 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i11_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i11_LC_5_10_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i11_LC_5_10_3  (
            .in0(N__53520),
            .in1(N__46695),
            .in2(N__17831),
            .in3(N__46076),
            .lcout(cmd_rdadctmp_11_adj_1065),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51244),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i15_LC_5_10_4 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i15_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i15_LC_5_10_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i15_LC_5_10_4  (
            .in0(N__17714),
            .in1(N__27415),
            .in2(N__18054),
            .in3(N__26846),
            .lcout(cmd_rdadctmp_15_adj_1134),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51244),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i13_LC_5_10_5 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i13_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i13_LC_5_10_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i13_LC_5_10_5  (
            .in0(N__53521),
            .in1(N__17808),
            .in2(N__17868),
            .in3(N__46077),
            .lcout(cmd_rdadctmp_13_adj_1063),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51244),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i4_LC_5_10_6 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i4_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i4_LC_5_10_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i4_LC_5_10_6  (
            .in0(N__53696),
            .in1(N__17884),
            .in2(N__17813),
            .in3(N__53524),
            .lcout(buf_adcdata2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51244),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i14_LC_5_10_7 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i14_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i14_LC_5_10_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i14_LC_5_10_7  (
            .in0(N__53522),
            .in1(N__17844),
            .in2(N__17869),
            .in3(N__46078),
            .lcout(cmd_rdadctmp_14_adj_1062),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51244),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i12_LC_5_11_6 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i12_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i12_LC_5_11_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i12_LC_5_11_6  (
            .in0(N__17830),
            .in1(N__46058),
            .in2(N__17812),
            .in3(N__53356),
            .lcout(cmd_rdadctmp_12_adj_1064),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51262),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i5_LC_5_11_7 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i5_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i5_LC_5_11_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i5_LC_5_11_7  (
            .in0(N__53049),
            .in1(N__17788),
            .in2(N__19595),
            .in3(N__52845),
            .lcout(buf_adcdata1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51262),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i7_LC_5_12_0 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i7_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i7_LC_5_12_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i7_LC_5_12_0  (
            .in0(N__53051),
            .in1(N__17770),
            .in2(N__19793),
            .in3(N__52847),
            .lcout(buf_adcdata1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i5_LC_5_12_2 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i5_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i5_LC_5_12_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i5_LC_5_12_2  (
            .in0(N__25940),
            .in1(N__17745),
            .in2(N__27515),
            .in3(N__17728),
            .lcout(buf_adcdata4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i13_LC_5_12_3 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i13_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i13_LC_5_12_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i13_LC_5_12_3  (
            .in0(N__27482),
            .in1(N__18151),
            .in2(N__17729),
            .in3(N__26839),
            .lcout(cmd_rdadctmp_13_adj_1136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i14_LC_5_12_4 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i14_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i14_LC_5_12_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i14_LC_5_12_4  (
            .in0(N__26838),
            .in1(N__17727),
            .in2(N__17709),
            .in3(N__27485),
            .lcout(cmd_rdadctmp_14_adj_1135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i6_LC_5_12_6 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i6_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i6_LC_5_12_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i6_LC_5_12_6  (
            .in0(N__25941),
            .in1(N__17673),
            .in2(N__17710),
            .in3(N__27484),
            .lcout(buf_adcdata4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i16_LC_5_12_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i16_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i16_LC_5_12_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i16_LC_5_12_7  (
            .in0(N__27483),
            .in1(N__18055),
            .in2(N__19441),
            .in3(N__26840),
            .lcout(cmd_rdadctmp_16_adj_1133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51276),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i0_LC_5_13_1 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i0_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i0_LC_5_13_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i0_LC_5_13_1  (
            .in0(N__25937),
            .in1(N__18015),
            .in2(N__18275),
            .in3(N__27451),
            .lcout(buf_adcdata4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51289),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i1_LC_5_13_2 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i1_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i1_LC_5_13_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i1_LC_5_13_2  (
            .in0(N__27447),
            .in1(N__25938),
            .in2(N__17954),
            .in3(N__17976),
            .lcout(buf_adcdata4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51289),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i9_LC_5_13_3 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i9_LC_5_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i9_LC_5_13_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i9_LC_5_13_3  (
            .in0(N__26843),
            .in1(N__17946),
            .in2(N__18274),
            .in3(N__27453),
            .lcout(cmd_rdadctmp_9_adj_1140),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51289),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i10_LC_5_13_4 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i10_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i10_LC_5_13_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i10_LC_5_13_4  (
            .in0(N__27449),
            .in1(N__17931),
            .in2(N__17953),
            .in3(N__26844),
            .lcout(cmd_rdadctmp_10_adj_1139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51289),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i11_LC_5_13_5 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i11_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i11_LC_5_13_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i11_LC_5_13_5  (
            .in0(N__26841),
            .in1(N__18219),
            .in2(N__17936),
            .in3(N__27452),
            .lcout(cmd_rdadctmp_11_adj_1138),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51289),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i2_LC_5_13_6 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i2_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i2_LC_5_13_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i2_LC_5_13_6  (
            .in0(N__27448),
            .in1(N__25939),
            .in2(N__17910),
            .in3(N__17935),
            .lcout(buf_adcdata4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51289),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i5_LC_5_13_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i5_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i5_LC_5_13_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i5_LC_5_13_7  (
            .in0(N__26842),
            .in1(N__27450),
            .in2(N__18203),
            .in3(N__18253),
            .lcout(cmd_rdadctmp_5_adj_1144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51289),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i7_LC_5_14_2 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i7_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i7_LC_5_14_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i7_LC_5_14_2  (
            .in0(N__26834),
            .in1(N__18242),
            .in2(N__27514),
            .in3(N__18283),
            .lcout(cmd_rdadctmp_7_adj_1142),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i8_LC_5_14_3 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i8_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i8_LC_5_14_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i8_LC_5_14_3  (
            .in0(N__18267),
            .in1(N__27472),
            .in2(N__18287),
            .in3(N__26837),
            .lcout(cmd_rdadctmp_8_adj_1141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i6_LC_5_14_4 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i6_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i6_LC_5_14_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i6_LC_5_14_4  (
            .in0(N__26833),
            .in1(N__18241),
            .in2(N__27513),
            .in3(N__18254),
            .lcout(cmd_rdadctmp_6_adj_1143),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i12_LC_5_14_5 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i12_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i12_LC_5_14_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i12_LC_5_14_5  (
            .in0(N__18220),
            .in1(N__27470),
            .in2(N__18150),
            .in3(N__26835),
            .lcout(cmd_rdadctmp_12_adj_1137),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i4_LC_5_14_6 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i4_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i4_LC_5_14_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i4_LC_5_14_6  (
            .in0(N__26832),
            .in1(N__18187),
            .in2(N__27512),
            .in3(N__18202),
            .lcout(cmd_rdadctmp_4_adj_1145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i3_LC_5_14_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i3_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i3_LC_5_14_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i3_LC_5_14_7  (
            .in0(N__18175),
            .in1(N__27471),
            .in2(N__18188),
            .in3(N__26836),
            .lcout(cmd_rdadctmp_3_adj_1146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51299),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i2_LC_5_15_2 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i2_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i2_LC_5_15_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i2_LC_5_15_2  (
            .in0(N__19847),
            .in1(N__27459),
            .in2(N__18176),
            .in3(N__26845),
            .lcout(cmd_rdadctmp_2_adj_1147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51308),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i4_LC_6_5_0 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i4_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i4_LC_6_5_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i4_LC_6_5_0  (
            .in0(N__25966),
            .in1(N__18121),
            .in2(N__18161),
            .in3(N__27526),
            .lcout(buf_adcdata4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51137),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1481_i7_4_lut_LC_6_5_1.C_ON=1'b0;
    defparam mux_1481_i7_4_lut_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam mux_1481_i7_4_lut_LC_6_5_1.LUT_INIT=16'b1000100011011000;
    LogicCell40 mux_1481_i7_4_lut_LC_6_5_1 (
            .in0(N__47324),
            .in1(N__18101),
            .in2(N__19528),
            .in3(N__48087),
            .lcout(n4146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1481_i1_4_lut_LC_6_5_4.C_ON=1'b0;
    defparam mux_1481_i1_4_lut_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam mux_1481_i1_4_lut_LC_6_5_4.LUT_INIT=16'b1000101110001000;
    LogicCell40 mux_1481_i1_4_lut_LC_6_5_4 (
            .in0(N__18077),
            .in1(N__47326),
            .in2(N__48092),
            .in3(N__43814),
            .lcout(n4152),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1481_i8_4_lut_LC_6_5_6.C_ON=1'b0;
    defparam mux_1481_i8_4_lut_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam mux_1481_i8_4_lut_LC_6_5_6.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1481_i8_4_lut_LC_6_5_6 (
            .in0(N__18359),
            .in1(N__48091),
            .in2(N__18715),
            .in3(N__47325),
            .lcout(n4145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i1_LC_6_6_0.C_ON=1'b0;
    defparam comm_buf_2__i1_LC_6_6_0.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i1_LC_6_6_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i1_LC_6_6_0 (
            .in0(N__50268),
            .in1(N__44155),
            .in2(_gnd_net_),
            .in3(N__27545),
            .lcout(comm_buf_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51148),
            .ce(N__18375),
            .sr(N__18614));
    defparam comm_buf_2__i0_LC_6_6_1.C_ON=1'b0;
    defparam comm_buf_2__i0_LC_6_6_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i0_LC_6_6_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_buf_2__i0_LC_6_6_1 (
            .in0(N__50269),
            .in1(N__18341),
            .in2(_gnd_net_),
            .in3(N__39214),
            .lcout(comm_buf_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51148),
            .ce(N__18375),
            .sr(N__18614));
    defparam i1_2_lut_adj_270_LC_6_7_0.C_ON=1'b0;
    defparam i1_2_lut_adj_270_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_270_LC_6_7_0.LUT_INIT=16'b1111111101010101;
    LogicCell40 i1_2_lut_adj_270_LC_6_7_0 (
            .in0(N__49536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52310),
            .lcout(n15221),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_3_lut_3_lut_LC_6_7_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_3_lut_3_lut_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_3_lut_3_lut_LC_6_7_1.LUT_INIT=16'b1111111110001000;
    LogicCell40 i1_2_lut_3_lut_3_lut_3_lut_LC_6_7_1 (
            .in0(N__52309),
            .in1(N__50267),
            .in2(_gnd_net_),
            .in3(N__49535),
            .lcout(n15131),
            .ltout(n15131_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_195_LC_6_7_2.C_ON=1'b0;
    defparam i1_4_lut_adj_195_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_195_LC_6_7_2.LUT_INIT=16'b1011000010100000;
    LogicCell40 i1_4_lut_adj_195_LC_6_7_2 (
            .in0(N__25558),
            .in1(N__50604),
            .in2(N__18335),
            .in3(N__27809),
            .lcout(n8738),
            .ltout(n8738_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7484_2_lut_LC_6_7_3.C_ON=1'b0;
    defparam i7484_2_lut_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam i7484_2_lut_LC_6_7_3.LUT_INIT=16'b1010000010100000;
    LogicCell40 i7484_2_lut_LC_6_7_3 (
            .in0(N__52312),
            .in1(_gnd_net_),
            .in2(N__18332),
            .in3(_gnd_net_),
            .lcout(n10590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_233_LC_6_7_4.C_ON=1'b0;
    defparam i1_4_lut_adj_233_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_233_LC_6_7_4.LUT_INIT=16'b1010001010100000;
    LogicCell40 i1_4_lut_adj_233_LC_6_7_4 (
            .in0(N__42839),
            .in1(N__50605),
            .in2(N__25572),
            .in3(N__27734),
            .lcout(n8847),
            .ltout(n8847_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7505_2_lut_LC_6_7_5.C_ON=1'b0;
    defparam i7505_2_lut_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam i7505_2_lut_LC_6_7_5.LUT_INIT=16'b1010000010100000;
    LogicCell40 i7505_2_lut_LC_6_7_5 (
            .in0(N__52313),
            .in1(_gnd_net_),
            .in2(N__18302),
            .in3(_gnd_net_),
            .lcout(n10611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_201_LC_6_7_6.C_ON=1'b0;
    defparam i1_4_lut_adj_201_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_201_LC_6_7_6.LUT_INIT=16'b1010001010100000;
    LogicCell40 i1_4_lut_adj_201_LC_6_7_6 (
            .in0(N__42838),
            .in1(N__50603),
            .in2(N__25571),
            .in3(N__27827),
            .lcout(n8787),
            .ltout(n8787_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7491_2_lut_LC_6_7_7.C_ON=1'b0;
    defparam i7491_2_lut_LC_6_7_7.SEQ_MODE=4'b0000;
    defparam i7491_2_lut_LC_6_7_7.LUT_INIT=16'b1010000010100000;
    LogicCell40 i7491_2_lut_LC_6_7_7 (
            .in0(N__52311),
            .in1(_gnd_net_),
            .in2(N__18428),
            .in3(_gnd_net_),
            .lcout(n10599),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1481_i3_4_lut_LC_6_8_0.C_ON=1'b0;
    defparam mux_1481_i3_4_lut_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam mux_1481_i3_4_lut_LC_6_8_0.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1481_i3_4_lut_LC_6_8_0 (
            .in0(N__18425),
            .in1(N__48069),
            .in2(N__18475),
            .in3(N__47319),
            .lcout(),
            .ltout(n4150_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i2_LC_6_8_1.C_ON=1'b0;
    defparam comm_buf_2__i2_LC_6_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i2_LC_6_8_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_2__i2_LC_6_8_1 (
            .in0(N__40122),
            .in1(_gnd_net_),
            .in2(N__18407),
            .in3(N__50088),
            .lcout(comm_buf_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51178),
            .ce(N__18376),
            .sr(N__18612));
    defparam comm_buf_2__i3_LC_6_8_3.C_ON=1'b0;
    defparam comm_buf_2__i3_LC_6_8_3.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i3_LC_6_8_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i3_LC_6_8_3 (
            .in0(N__44907),
            .in1(N__32582),
            .in2(_gnd_net_),
            .in3(N__50089),
            .lcout(comm_buf_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51178),
            .ce(N__18376),
            .sr(N__18612));
    defparam mux_1481_i5_4_lut_LC_6_8_4.C_ON=1'b0;
    defparam mux_1481_i5_4_lut_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam mux_1481_i5_4_lut_LC_6_8_4.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1481_i5_4_lut_LC_6_8_4 (
            .in0(N__18404),
            .in1(N__48070),
            .in2(N__18764),
            .in3(N__47320),
            .lcout(),
            .ltout(n4148_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i4_LC_6_8_5.C_ON=1'b0;
    defparam comm_buf_2__i4_LC_6_8_5.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i4_LC_6_8_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_2__i4_LC_6_8_5 (
            .in0(N__39947),
            .in1(_gnd_net_),
            .in2(N__18395),
            .in3(N__50090),
            .lcout(comm_buf_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51178),
            .ce(N__18376),
            .sr(N__18612));
    defparam mux_1481_i6_4_lut_LC_6_8_6.C_ON=1'b0;
    defparam mux_1481_i6_4_lut_LC_6_8_6.SEQ_MODE=4'b0000;
    defparam mux_1481_i6_4_lut_LC_6_8_6.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1481_i6_4_lut_LC_6_8_6 (
            .in0(N__18392),
            .in1(N__48071),
            .in2(N__19565),
            .in3(N__47321),
            .lcout(),
            .ltout(n4147_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i5_LC_6_8_7.C_ON=1'b0;
    defparam comm_buf_2__i5_LC_6_8_7.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i5_LC_6_8_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_2__i5_LC_6_8_7 (
            .in0(_gnd_net_),
            .in1(N__39809),
            .in2(N__18380),
            .in3(N__50091),
            .lcout(comm_buf_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51178),
            .ce(N__18376),
            .sr(N__18612));
    defparam i6_4_lut_adj_192_LC_6_9_0.C_ON=1'b0;
    defparam i6_4_lut_adj_192_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_192_LC_6_9_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_adj_192_LC_6_9_0 (
            .in0(N__18584),
            .in1(N__18569),
            .in2(N__18554),
            .in3(N__18533),
            .lcout(n14_adj_1163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i0_LC_6_9_2.C_ON=1'b0;
    defparam comm_buf_4__i0_LC_6_9_2.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i0_LC_6_9_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_4__i0_LC_6_9_2 (
            .in0(N__24305),
            .in1(N__50278),
            .in2(_gnd_net_),
            .in3(N__39213),
            .lcout(comm_buf_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51196),
            .ce(N__25450),
            .sr(N__20088));
    defparam comm_buf_4__i1_LC_6_9_4.C_ON=1'b0;
    defparam comm_buf_4__i1_LC_6_9_4.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i1_LC_6_9_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i1_LC_6_9_4 (
            .in0(N__44179),
            .in1(N__42632),
            .in2(_gnd_net_),
            .in3(N__50279),
            .lcout(comm_buf_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51196),
            .ce(N__25450),
            .sr(N__20088));
    defparam mux_1457_i3_4_lut_LC_6_9_5.C_ON=1'b0;
    defparam mux_1457_i3_4_lut_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam mux_1457_i3_4_lut_LC_6_9_5.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1457_i3_4_lut_LC_6_9_5 (
            .in0(N__18506),
            .in1(N__48037),
            .in2(N__19709),
            .in3(N__47290),
            .lcout(),
            .ltout(n4062_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i2_LC_6_9_6.C_ON=1'b0;
    defparam comm_buf_4__i2_LC_6_9_6.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i2_LC_6_9_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_4__i2_LC_6_9_6 (
            .in0(_gnd_net_),
            .in1(N__40123),
            .in2(N__18485),
            .in3(N__50280),
            .lcout(comm_buf_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51196),
            .ce(N__25450),
            .sr(N__20088));
    defparam comm_buf_4__i3_LC_6_10_0.C_ON=1'b0;
    defparam comm_buf_4__i3_LC_6_10_0.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i3_LC_6_10_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i3_LC_6_10_0 (
            .in0(N__44908),
            .in1(N__26516),
            .in2(_gnd_net_),
            .in3(N__50281),
            .lcout(comm_buf_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51213),
            .ce(N__25457),
            .sr(N__20102));
    defparam \ADC_VAC3.ADC_DATA_i2_LC_6_11_1 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i2_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i2_LC_6_11_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i2_LC_6_11_1  (
            .in0(N__49190),
            .in1(N__44356),
            .in2(N__19472),
            .in3(N__18459),
            .lcout(buf_adcdata3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51230),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i11_LC_6_11_3 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i11_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i11_LC_6_11_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i11_LC_6_11_3  (
            .in0(N__49193),
            .in1(N__18438),
            .in2(N__19471),
            .in3(N__48840),
            .lcout(cmd_rdadctmp_11_adj_1101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51230),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i12_LC_6_11_4 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i12_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i12_LC_6_11_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i12_LC_6_11_4  (
            .in0(N__48839),
            .in1(N__18648),
            .in2(N__18443),
            .in3(N__49194),
            .lcout(cmd_rdadctmp_12_adj_1100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51230),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i3_LC_6_11_5 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i3_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i3_LC_6_11_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i3_LC_6_11_5  (
            .in0(N__49191),
            .in1(N__44357),
            .in2(N__32619),
            .in3(N__18442),
            .lcout(buf_adcdata3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51230),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i3_LC_6_11_6 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i3_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i3_LC_6_11_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i3_LC_6_11_6  (
            .in0(N__52848),
            .in1(N__53015),
            .in2(N__20525),
            .in3(N__18778),
            .lcout(buf_adcdata1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51230),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i4_LC_6_11_7 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i4_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i4_LC_6_11_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i4_LC_6_11_7  (
            .in0(N__49192),
            .in1(N__44358),
            .in2(N__18655),
            .in3(N__18753),
            .lcout(buf_adcdata3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51230),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i1_LC_6_12_0 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i1_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i1_LC_6_12_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i1_LC_6_12_0  (
            .in0(N__52851),
            .in1(N__18665),
            .in2(N__18733),
            .in3(N__26115),
            .lcout(cmd_rdadctmp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51246),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i2_LC_6_12_2 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i2_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i2_LC_6_12_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i2_LC_6_12_2  (
            .in0(N__52852),
            .in1(N__18856),
            .in2(N__18734),
            .in3(N__26116),
            .lcout(cmd_rdadctmp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51246),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i7_LC_6_12_3 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i7_LC_6_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i7_LC_6_12_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC3.ADC_DATA_i7_LC_6_12_3  (
            .in0(N__44355),
            .in1(N__18708),
            .in2(N__21680),
            .in3(N__49201),
            .lcout(buf_adcdata3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51246),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i0_LC_6_12_4 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i0_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i0_LC_6_12_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i0_LC_6_12_4  (
            .in0(N__52849),
            .in1(N__18664),
            .in2(N__18686),
            .in3(N__26113),
            .lcout(cmd_rdadctmp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51246),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i13_LC_6_12_5 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i13_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i13_LC_6_12_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i13_LC_6_12_5  (
            .in0(N__18656),
            .in1(N__49200),
            .in2(N__20322),
            .in3(N__48814),
            .lcout(cmd_rdadctmp_13_adj_1099),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51246),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i13_LC_6_12_6 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i13_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i13_LC_6_12_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i13_LC_6_12_6  (
            .in0(N__52850),
            .in1(N__19488),
            .in2(N__19590),
            .in3(N__26114),
            .lcout(cmd_rdadctmp_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51246),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i4_LC_6_12_7 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i4_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i4_LC_6_12_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i4_LC_6_12_7  (
            .in0(N__53050),
            .in1(N__18628),
            .in2(N__19493),
            .in3(N__52853),
            .lcout(buf_adcdata1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51246),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.CS_37_LC_6_13_0 .C_ON=1'b0;
    defparam \ADC_VAC1.CS_37_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.CS_37_LC_6_13_0 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \ADC_VAC1.CS_37_LC_6_13_0  (
            .in0(N__18929),
            .in1(N__18896),
            .in2(N__19648),
            .in3(N__52674),
            .lcout(M_CS1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i24_LC_6_13_1 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i24_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i24_LC_6_13_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i24_LC_6_13_1  (
            .in0(N__52670),
            .in1(N__22715),
            .in2(N__48252),
            .in3(N__26069),
            .lcout(cmd_rdadctmp_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i8_LC_6_13_2 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i8_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i8_LC_6_13_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i8_LC_6_13_2  (
            .in0(N__26075),
            .in1(N__52677),
            .in2(N__22477),
            .in3(N__18845),
            .lcout(cmd_rdadctmp_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i3_LC_6_13_3 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i3_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i3_LC_6_13_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i3_LC_6_13_3  (
            .in0(N__52671),
            .in1(N__18857),
            .in2(N__18811),
            .in3(N__26070),
            .lcout(cmd_rdadctmp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i7_LC_6_13_4 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i7_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i7_LC_6_13_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i7_LC_6_13_4  (
            .in0(N__26074),
            .in1(N__18844),
            .in2(N__18836),
            .in3(N__52676),
            .lcout(cmd_rdadctmp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i6_LC_6_13_5 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i6_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i6_LC_6_13_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i6_LC_6_13_5  (
            .in0(N__52673),
            .in1(N__18832),
            .in2(N__18824),
            .in3(N__26073),
            .lcout(cmd_rdadctmp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i5_LC_6_13_6 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i5_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i5_LC_6_13_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i5_LC_6_13_6  (
            .in0(N__26072),
            .in1(N__18820),
            .in2(N__18797),
            .in3(N__52675),
            .lcout(cmd_rdadctmp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i4_LC_6_13_7 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i4_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i4_LC_6_13_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i4_LC_6_13_7  (
            .in0(N__52672),
            .in1(N__18793),
            .in2(N__18812),
            .in3(N__26071),
            .lcout(cmd_rdadctmp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51263),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.adc_state_i2_LC_6_14_1 .C_ON=1'b0;
    defparam \ADC_VAC1.adc_state_i2_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.adc_state_i2_LC_6_14_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_VAC1.adc_state_i2_LC_6_14_1  (
            .in0(N__52605),
            .in1(N__20627),
            .in2(_gnd_net_),
            .in3(N__20569),
            .lcout(DTRIG_N_957),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51277),
            .ce(N__19604),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.adc_state_i1_LC_6_14_2 .C_ON=1'b0;
    defparam \ADC_VAC1.adc_state_i1_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.adc_state_i1_LC_6_14_2 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \ADC_VAC1.adc_state_i1_LC_6_14_2  (
            .in0(N__20568),
            .in1(_gnd_net_),
            .in2(N__20643),
            .in3(N__52606),
            .lcout(adc_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51277),
            .ce(N__19604),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_224_LC_6_14_3.C_ON=1'b0;
    defparam i1_2_lut_adj_224_LC_6_14_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_224_LC_6_14_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_224_LC_6_14_3 (
            .in0(_gnd_net_),
            .in1(N__20623),
            .in2(_gnd_net_),
            .in3(N__20566),
            .lcout(n15168),
            .ltout(n15168_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i1_3_lut_LC_6_14_4 .C_ON=1'b0;
    defparam \ADC_VAC1.i1_3_lut_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i1_3_lut_LC_6_14_4 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \ADC_VAC1.i1_3_lut_LC_6_14_4  (
            .in0(N__19640),
            .in1(_gnd_net_),
            .in2(N__18923),
            .in3(N__52603),
            .lcout(n8272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_222_LC_6_14_6.C_ON=1'b0;
    defparam i1_4_lut_adj_222_LC_6_14_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_222_LC_6_14_6.LUT_INIT=16'b0010001100110010;
    LogicCell40 i1_4_lut_adj_222_LC_6_14_6 (
            .in0(N__20567),
            .in1(N__18907),
            .in2(N__20642),
            .in3(N__52604),
            .lcout(n14_adj_1039),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_298_LC_6_14_7.C_ON=1'b0;
    defparam i1_2_lut_adj_298_LC_6_14_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_298_LC_6_14_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_298_LC_6_14_7 (
            .in0(_gnd_net_),
            .in1(N__20622),
            .in2(_gnd_net_),
            .in3(N__20565),
            .lcout(n15153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.SCLK_35_LC_6_15_0 .C_ON=1'b0;
    defparam \ADC_VAC1.SCLK_35_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.SCLK_35_LC_6_15_0 .LUT_INIT=16'b1011000011100010;
    LogicCell40 \ADC_VAC1.SCLK_35_LC_6_15_0  (
            .in0(N__20638),
            .in1(N__52678),
            .in2(N__18880),
            .in3(N__20576),
            .lcout(M_SCLK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51290),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i1_4_lut_adj_6_LC_6_15_3 .C_ON=1'b0;
    defparam \ADC_VAC1.i1_4_lut_adj_6_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i1_4_lut_adj_6_LC_6_15_3 .LUT_INIT=16'b0001000100000010;
    LogicCell40 \ADC_VAC1.i1_4_lut_adj_6_LC_6_15_3  (
            .in0(N__20574),
            .in1(N__52616),
            .in2(N__19647),
            .in3(N__20636),
            .lcout(\ADC_VAC1.n9312 ),
            .ltout(\ADC_VAC1.n9312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i7561_2_lut_LC_6_15_4 .C_ON=1'b0;
    defparam \ADC_VAC1.i7561_2_lut_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i7561_2_lut_LC_6_15_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ADC_VAC1.i7561_2_lut_LC_6_15_4  (
            .in0(N__20637),
            .in1(_gnd_net_),
            .in2(N__18863),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC1.n10667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i12131_4_lut_LC_6_15_5 .C_ON=1'b0;
    defparam \ADC_VAC1.i12131_4_lut_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i12131_4_lut_LC_6_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC1.i12131_4_lut_LC_6_15_5  (
            .in0(N__18976),
            .in1(N__18991),
            .in2(N__19025),
            .in3(N__19006),
            .lcout(),
            .ltout(\ADC_VAC1.n15338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i12151_4_lut_LC_6_15_6 .C_ON=1'b0;
    defparam \ADC_VAC1.i12151_4_lut_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i12151_4_lut_LC_6_15_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC1.i12151_4_lut_LC_6_15_6  (
            .in0(N__18943),
            .in1(N__19039),
            .in2(N__18860),
            .in3(N__19141),
            .lcout(),
            .ltout(\ADC_VAC1.n15360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i12914_4_lut_LC_6_15_7 .C_ON=1'b0;
    defparam \ADC_VAC1.i12914_4_lut_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i12914_4_lut_LC_6_15_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_VAC1.i12914_4_lut_LC_6_15_7  (
            .in0(N__20575),
            .in1(N__18962),
            .in2(N__19043),
            .in3(N__52617),
            .lcout(\ADC_VAC1.n15553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.bit_cnt_i0_LC_6_16_0 .C_ON=1'b1;
    defparam \ADC_VAC1.bit_cnt_i0_LC_6_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i0_LC_6_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i0_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__19040),
            .in2(_gnd_net_),
            .in3(N__19028),
            .lcout(\ADC_VAC1.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_6_16_0_),
            .carryout(\ADC_VAC1.n13981 ),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam \ADC_VAC1.bit_cnt_i1_LC_6_16_1 .C_ON=1'b1;
    defparam \ADC_VAC1.bit_cnt_i1_LC_6_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i1_LC_6_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i1_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(N__19024),
            .in2(_gnd_net_),
            .in3(N__19010),
            .lcout(\ADC_VAC1.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC1.n13981 ),
            .carryout(\ADC_VAC1.n13982 ),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam \ADC_VAC1.bit_cnt_i2_LC_6_16_2 .C_ON=1'b1;
    defparam \ADC_VAC1.bit_cnt_i2_LC_6_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i2_LC_6_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i2_LC_6_16_2  (
            .in0(_gnd_net_),
            .in1(N__19007),
            .in2(_gnd_net_),
            .in3(N__18995),
            .lcout(\ADC_VAC1.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC1.n13982 ),
            .carryout(\ADC_VAC1.n13983 ),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam \ADC_VAC1.bit_cnt_i3_LC_6_16_3 .C_ON=1'b1;
    defparam \ADC_VAC1.bit_cnt_i3_LC_6_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i3_LC_6_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i3_LC_6_16_3  (
            .in0(_gnd_net_),
            .in1(N__18992),
            .in2(_gnd_net_),
            .in3(N__18980),
            .lcout(\ADC_VAC1.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC1.n13983 ),
            .carryout(\ADC_VAC1.n13984 ),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam \ADC_VAC1.bit_cnt_i4_LC_6_16_4 .C_ON=1'b1;
    defparam \ADC_VAC1.bit_cnt_i4_LC_6_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i4_LC_6_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i4_LC_6_16_4  (
            .in0(_gnd_net_),
            .in1(N__18977),
            .in2(_gnd_net_),
            .in3(N__18965),
            .lcout(\ADC_VAC1.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC1.n13984 ),
            .carryout(\ADC_VAC1.n13985 ),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam \ADC_VAC1.bit_cnt_i5_LC_6_16_5 .C_ON=1'b1;
    defparam \ADC_VAC1.bit_cnt_i5_LC_6_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i5_LC_6_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i5_LC_6_16_5  (
            .in0(_gnd_net_),
            .in1(N__18961),
            .in2(_gnd_net_),
            .in3(N__18947),
            .lcout(\ADC_VAC1.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC1.n13985 ),
            .carryout(\ADC_VAC1.n13986 ),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam \ADC_VAC1.bit_cnt_i6_LC_6_16_6 .C_ON=1'b1;
    defparam \ADC_VAC1.bit_cnt_i6_LC_6_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i6_LC_6_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i6_LC_6_16_6  (
            .in0(_gnd_net_),
            .in1(N__18944),
            .in2(_gnd_net_),
            .in3(N__18932),
            .lcout(\ADC_VAC1.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC1.n13986 ),
            .carryout(\ADC_VAC1.n13987 ),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam \ADC_VAC1.bit_cnt_i7_LC_6_16_7 .C_ON=1'b0;
    defparam \ADC_VAC1.bit_cnt_i7_LC_6_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.bit_cnt_i7_LC_6_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC1.bit_cnt_i7_LC_6_16_7  (
            .in0(_gnd_net_),
            .in1(N__19142),
            .in2(_gnd_net_),
            .in3(N__19145),
            .lcout(\ADC_VAC1.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51300),
            .ce(N__19130),
            .sr(N__19121));
    defparam comm_index_0__bdd_4_lut_13254_LC_7_5_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13254_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13254_LC_7_5_0.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_0__bdd_4_lut_13254_LC_7_5_0 (
            .in0(N__38848),
            .in1(N__23537),
            .in2(N__22205),
            .in3(N__33206),
            .lcout(),
            .ltout(n16470_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16470_bdd_4_lut_LC_7_5_1.C_ON=1'b0;
    defparam n16470_bdd_4_lut_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam n16470_bdd_4_lut_LC_7_5_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16470_bdd_4_lut_LC_7_5_1 (
            .in0(N__33207),
            .in1(N__20147),
            .in2(N__19115),
            .in3(N__19112),
            .lcout(n16473),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13205_LC_7_5_4.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13205_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13205_LC_7_5_4.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_0__bdd_4_lut_13205_LC_7_5_4 (
            .in0(N__38849),
            .in1(N__19100),
            .in2(N__19052),
            .in3(N__33208),
            .lcout(),
            .ltout(n16416_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16416_bdd_4_lut_LC_7_5_5.C_ON=1'b0;
    defparam n16416_bdd_4_lut_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam n16416_bdd_4_lut_LC_7_5_5.LUT_INIT=16'b1110001111100000;
    LogicCell40 n16416_bdd_4_lut_LC_7_5_5 (
            .in0(N__37878),
            .in1(N__33205),
            .in2(N__19088),
            .in3(N__33785),
            .lcout(),
            .ltout(n16419_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i981538_i1_3_lut_LC_7_5_6.C_ON=1'b0;
    defparam i981538_i1_3_lut_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam i981538_i1_3_lut_LC_7_5_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 i981538_i1_3_lut_LC_7_5_6 (
            .in0(_gnd_net_),
            .in1(N__19085),
            .in2(N__19079),
            .in3(N__33535),
            .lcout(),
            .ltout(n7_adj_1238_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i5_LC_7_5_7.C_ON=1'b0;
    defparam comm_tx_buf_i5_LC_7_5_7.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i5_LC_7_5_7.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_tx_buf_i5_LC_7_5_7 (
            .in0(N__33536),
            .in1(N__20936),
            .in2(N__19076),
            .in3(N__33352),
            .lcout(comm_tx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51126),
            .ce(N__43110),
            .sr(N__22393));
    defparam mux_1469_i6_4_lut_LC_7_6_0.C_ON=1'b0;
    defparam mux_1469_i6_4_lut_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam mux_1469_i6_4_lut_LC_7_6_0.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1469_i6_4_lut_LC_7_6_0 (
            .in0(N__19073),
            .in1(N__48013),
            .in2(N__23177),
            .in3(N__47335),
            .lcout(),
            .ltout(n4103_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i5_LC_7_6_1.C_ON=1'b0;
    defparam comm_buf_3__i5_LC_7_6_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i5_LC_7_6_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_3__i5_LC_7_6_1 (
            .in0(N__39796),
            .in1(_gnd_net_),
            .in2(N__19055),
            .in3(N__50112),
            .lcout(comm_buf_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51138),
            .ce(N__19202),
            .sr(N__19178));
    defparam comm_buf_3__i6_LC_7_6_3.C_ON=1'b0;
    defparam comm_buf_3__i6_LC_7_6_3.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i6_LC_7_6_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i6_LC_7_6_3 (
            .in0(N__40692),
            .in1(N__29045),
            .in2(_gnd_net_),
            .in3(N__50113),
            .lcout(comm_buf_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51138),
            .ce(N__19202),
            .sr(N__19178));
    defparam comm_buf_3__i7_LC_7_6_5.C_ON=1'b0;
    defparam comm_buf_3__i7_LC_7_6_5.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i7_LC_7_6_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i7_LC_7_6_5 (
            .in0(N__39360),
            .in1(N__45836),
            .in2(_gnd_net_),
            .in3(N__50114),
            .lcout(comm_buf_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51138),
            .ce(N__19202),
            .sr(N__19178));
    defparam comm_buf_3__i0_LC_7_7_1.C_ON=1'b0;
    defparam comm_buf_3__i0_LC_7_7_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i0_LC_7_7_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_3__i0_LC_7_7_1 (
            .in0(N__46718),
            .in1(N__50337),
            .in2(_gnd_net_),
            .in3(N__39209),
            .lcout(comm_buf_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51149),
            .ce(N__19201),
            .sr(N__19174));
    defparam mux_1469_i2_4_lut_LC_7_7_2.C_ON=1'b0;
    defparam mux_1469_i2_4_lut_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam mux_1469_i2_4_lut_LC_7_7_2.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1469_i2_4_lut_LC_7_7_2 (
            .in0(N__19247),
            .in1(N__48006),
            .in2(N__25799),
            .in3(N__47088),
            .lcout(),
            .ltout(n4107_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i1_LC_7_7_3.C_ON=1'b0;
    defparam comm_buf_3__i1_LC_7_7_3.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i1_LC_7_7_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_3__i1_LC_7_7_3 (
            .in0(N__44171),
            .in1(_gnd_net_),
            .in2(N__19226),
            .in3(N__50338),
            .lcout(comm_buf_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51149),
            .ce(N__19201),
            .sr(N__19174));
    defparam mux_1469_i3_4_lut_LC_7_7_4.C_ON=1'b0;
    defparam mux_1469_i3_4_lut_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam mux_1469_i3_4_lut_LC_7_7_4.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1469_i3_4_lut_LC_7_7_4 (
            .in0(N__19223),
            .in1(N__48005),
            .in2(N__19285),
            .in3(N__47087),
            .lcout(comm_buf_3_7_N_501_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i4_LC_7_7_7.C_ON=1'b0;
    defparam comm_buf_3__i4_LC_7_7_7.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i4_LC_7_7_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i4_LC_7_7_7 (
            .in0(N__39939),
            .in1(N__21554),
            .in2(_gnd_net_),
            .in3(N__50339),
            .lcout(comm_buf_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51149),
            .ce(N__19201),
            .sr(N__19174));
    defparam i12238_3_lut_LC_7_8_1.C_ON=1'b0;
    defparam i12238_3_lut_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam i12238_3_lut_LC_7_8_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12238_3_lut_LC_7_8_1 (
            .in0(N__22121),
            .in1(N__38840),
            .in2(_gnd_net_),
            .in3(N__23453),
            .lcout(n15448),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12178_3_lut_LC_7_8_2.C_ON=1'b0;
    defparam i12178_3_lut_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam i12178_3_lut_LC_7_8_2.LUT_INIT=16'b1111101001010000;
    LogicCell40 i12178_3_lut_LC_7_8_2 (
            .in0(N__38842),
            .in1(_gnd_net_),
            .in2(N__19154),
            .in3(N__21125),
            .lcout(),
            .ltout(n15388_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16386_bdd_4_lut_LC_7_8_3.C_ON=1'b0;
    defparam n16386_bdd_4_lut_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam n16386_bdd_4_lut_LC_7_8_3.LUT_INIT=16'b1011100110101000;
    LogicCell40 n16386_bdd_4_lut_LC_7_8_3 (
            .in0(N__19301),
            .in1(N__33522),
            .in2(N__19331),
            .in3(N__29117),
            .lcout(),
            .ltout(n16389_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i2_LC_7_8_4.C_ON=1'b0;
    defparam comm_tx_buf_i2_LC_7_8_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i2_LC_7_8_4.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_tx_buf_i2_LC_7_8_4 (
            .in0(N__33523),
            .in1(N__21029),
            .in2(N__19328),
            .in3(N__33347),
            .lcout(comm_tx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51161),
            .ce(N__43127),
            .sr(N__22348));
    defparam i12237_3_lut_LC_7_8_5.C_ON=1'b0;
    defparam i12237_3_lut_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam i12237_3_lut_LC_7_8_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 i12237_3_lut_LC_7_8_5 (
            .in0(N__19325),
            .in1(N__38841),
            .in2(_gnd_net_),
            .in3(N__19319),
            .lcout(),
            .ltout(n15447_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_13182_LC_7_8_6.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_13182_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_13182_LC_7_8_6.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_index_1__bdd_4_lut_13182_LC_7_8_6 (
            .in0(N__33521),
            .in1(N__19310),
            .in2(N__19304),
            .in3(N__33212),
            .lcout(n16386),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7554_3_lut_LC_7_9_1.C_ON=1'b0;
    defparam i7554_3_lut_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam i7554_3_lut_LC_7_9_1.LUT_INIT=16'b1000100010101010;
    LogicCell40 i7554_3_lut_LC_7_9_1 (
            .in0(N__43078),
            .in1(N__52444),
            .in2(_gnd_net_),
            .in3(N__39263),
            .lcout(n10660),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i18_LC_7_9_2 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i18_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i18_LC_7_9_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i18_LC_7_9_2  (
            .in0(N__25945),
            .in1(N__19278),
            .in2(N__25751),
            .in3(N__27511),
            .lcout(buf_adcdata4_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51179),
            .ce(),
            .sr(_gnd_net_));
    defparam i7498_2_lut_LC_7_9_3.C_ON=1'b0;
    defparam i7498_2_lut_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam i7498_2_lut_LC_7_9_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i7498_2_lut_LC_7_9_3 (
            .in0(_gnd_net_),
            .in1(N__52445),
            .in2(_gnd_net_),
            .in3(N__25448),
            .lcout(n10604),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9698_2_lut_3_lut_LC_7_9_5.C_ON=1'b0;
    defparam i9698_2_lut_3_lut_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam i9698_2_lut_3_lut_LC_7_9_5.LUT_INIT=16'b0000000000100010;
    LogicCell40 i9698_2_lut_3_lut_LC_7_9_5 (
            .in0(N__33971),
            .in1(N__50110),
            .in2(_gnd_net_),
            .in3(N__49537),
            .lcout(n14_adj_1169),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i1_3_lut_LC_7_9_7.C_ON=1'b0;
    defparam mux_1498_i1_3_lut_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam mux_1498_i1_3_lut_LC_7_9_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_1498_i1_3_lut_LC_7_9_7 (
            .in0(N__33871),
            .in1(N__24512),
            .in2(_gnd_net_),
            .in3(N__48014),
            .lcout(n4209),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12187_3_lut_LC_7_10_0.C_ON=1'b0;
    defparam i12187_3_lut_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam i12187_3_lut_LC_7_10_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12187_3_lut_LC_7_10_0 (
            .in0(N__21116),
            .in1(N__19259),
            .in2(_gnd_net_),
            .in3(N__38845),
            .lcout(n15397),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12213_3_lut_LC_7_10_1.C_ON=1'b0;
    defparam i12213_3_lut_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam i12213_3_lut_LC_7_10_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 i12213_3_lut_LC_7_10_1 (
            .in0(N__38843),
            .in1(N__19409),
            .in2(_gnd_net_),
            .in3(N__19403),
            .lcout(n15423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13230_LC_7_10_2.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13230_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13230_LC_7_10_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13230_LC_7_10_2 (
            .in0(N__23672),
            .in1(N__33209),
            .in2(N__22025),
            .in3(N__38844),
            .lcout(),
            .ltout(n16440_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16440_bdd_4_lut_LC_7_10_3.C_ON=1'b0;
    defparam n16440_bdd_4_lut_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam n16440_bdd_4_lut_LC_7_10_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16440_bdd_4_lut_LC_7_10_3 (
            .in0(N__33210),
            .in1(N__23288),
            .in2(N__19391),
            .in3(N__21092),
            .lcout(n16443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_13225_LC_7_10_4.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_13225_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_13225_LC_7_10_4.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_index_1__bdd_4_lut_13225_LC_7_10_4 (
            .in0(N__33532),
            .in1(N__33211),
            .in2(N__19388),
            .in3(N__20981),
            .lcout(),
            .ltout(n16392_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16392_bdd_4_lut_LC_7_10_5.C_ON=1'b0;
    defparam n16392_bdd_4_lut_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam n16392_bdd_4_lut_LC_7_10_5.LUT_INIT=16'b1111000011001010;
    LogicCell40 n16392_bdd_4_lut_LC_7_10_5 (
            .in0(N__31109),
            .in1(N__19379),
            .in2(N__19373),
            .in3(N__33533),
            .lcout(),
            .ltout(n16395_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i3_LC_7_10_6.C_ON=1'b0;
    defparam comm_tx_buf_i3_LC_7_10_6.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i3_LC_7_10_6.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_tx_buf_i3_LC_7_10_6 (
            .in0(N__33534),
            .in1(N__19370),
            .in2(N__19364),
            .in3(N__33348),
            .lcout(comm_tx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51197),
            .ce(N__43126),
            .sr(N__22370));
    defparam \ADC_VAC2.cmd_rdadctmp_i31_LC_7_11_3 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i31_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i31_LC_7_11_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i31_LC_7_11_3  (
            .in0(N__53354),
            .in1(N__48212),
            .in2(N__48139),
            .in3(N__46081),
            .lcout(cmd_rdadctmp_31_adj_1045),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51214),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.SCLK_35_LC_7_11_4 .C_ON=1'b0;
    defparam \ADC_VAC2.SCLK_35_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.SCLK_35_LC_7_11_4 .LUT_INIT=16'b1011000011100010;
    LogicCell40 \ADC_VAC2.SCLK_35_LC_7_11_4  (
            .in0(N__36466),
            .in1(N__53355),
            .in2(N__19348),
            .in3(N__35609),
            .lcout(M_SCLK2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51214),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i8_LC_7_11_6 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i8_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i8_LC_7_11_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i8_LC_7_11_6  (
            .in0(N__49195),
            .in1(N__43827),
            .in2(N__23999),
            .in3(N__48815),
            .lcout(cmd_rdadctmp_8_adj_1104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51214),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i1_LC_7_11_7 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i1_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i1_LC_7_11_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC3.ADC_DATA_i1_LC_7_11_7  (
            .in0(N__44354),
            .in1(N__27571),
            .in2(N__20396),
            .in3(N__49196),
            .lcout(buf_adcdata3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51214),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i5_LC_7_12_0 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i5_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i5_LC_7_12_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC3.ADC_DATA_i5_LC_7_12_0  (
            .in0(N__44352),
            .in1(N__19551),
            .in2(N__20326),
            .in3(N__49199),
            .lcout(buf_adcdata3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51231),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i6_LC_7_12_1 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i6_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i6_LC_7_12_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i6_LC_7_12_1  (
            .in0(N__49197),
            .in1(N__44353),
            .in2(N__20297),
            .in3(N__19515),
            .lcout(buf_adcdata3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51231),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i12_LC_7_12_2 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i12_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i12_LC_7_12_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i12_LC_7_12_2  (
            .in0(N__20514),
            .in1(N__52836),
            .in2(N__19492),
            .in3(N__26126),
            .lcout(cmd_rdadctmp_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51231),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i10_LC_7_12_3 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i10_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i10_LC_7_12_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i10_LC_7_12_3  (
            .in0(N__49198),
            .in1(N__20392),
            .in2(N__19470),
            .in3(N__48763),
            .lcout(cmd_rdadctmp_10_adj_1102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51231),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i8_LC_7_13_1 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i8_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i8_LC_7_13_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i8_LC_7_13_1  (
            .in0(N__27372),
            .in1(N__25926),
            .in2(N__24336),
            .in3(N__19448),
            .lcout(buf_adcdata4_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51247),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i9_LC_7_13_2 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i9_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i9_LC_7_13_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i9_LC_7_13_2  (
            .in0(N__25925),
            .in1(N__27376),
            .in2(N__42652),
            .in3(N__19423),
            .lcout(buf_adcdata4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51247),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i17_LC_7_13_3 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i17_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i17_LC_7_13_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i17_LC_7_13_3  (
            .in0(N__27373),
            .in1(N__19447),
            .in2(N__19424),
            .in3(N__26855),
            .lcout(cmd_rdadctmp_17_adj_1132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51247),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i18_LC_7_13_4 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i18_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i18_LC_7_13_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i18_LC_7_13_4  (
            .in0(N__26854),
            .in1(N__19422),
            .in2(N__19726),
            .in3(N__27378),
            .lcout(cmd_rdadctmp_18_adj_1131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51247),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i19_LC_7_13_5 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i19_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i19_LC_7_13_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i19_LC_7_13_5  (
            .in0(N__27374),
            .in1(N__19722),
            .in2(N__22500),
            .in3(N__26856),
            .lcout(cmd_rdadctmp_19_adj_1130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51247),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i10_LC_7_13_6 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i10_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i10_LC_7_13_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i10_LC_7_13_6  (
            .in0(N__25924),
            .in1(N__19695),
            .in2(N__19727),
            .in3(N__27377),
            .lcout(buf_adcdata4_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51247),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i20_LC_7_13_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i20_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i20_LC_7_13_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i20_LC_7_13_7  (
            .in0(N__27375),
            .in1(N__22656),
            .in2(N__22501),
            .in3(N__26857),
            .lcout(cmd_rdadctmp_20_adj_1129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51247),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i1_4_lut_LC_7_14_1 .C_ON=1'b0;
    defparam \ADC_VAC1.i1_4_lut_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i1_4_lut_LC_7_14_1 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_VAC1.i1_4_lut_LC_7_14_1  (
            .in0(N__20632),
            .in1(N__52619),
            .in2(N__19658),
            .in3(N__30658),
            .lcout(),
            .ltout(\ADC_VAC1.n15263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i1_2_lut_LC_7_14_2 .C_ON=1'b0;
    defparam \ADC_VAC1.i1_2_lut_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i1_2_lut_LC_7_14_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \ADC_VAC1.i1_2_lut_LC_7_14_2  (
            .in0(N__20573),
            .in1(_gnd_net_),
            .in2(N__19673),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC1.n15264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.adc_state_i0_LC_7_14_5 .C_ON=1'b0;
    defparam \ADC_VAC1.adc_state_i0_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.adc_state_i0_LC_7_14_5 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \ADC_VAC1.adc_state_i0_LC_7_14_5  (
            .in0(N__20580),
            .in1(N__52620),
            .in2(N__20644),
            .in3(N__19670),
            .lcout(adc_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51264),
            .ce(N__19664),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i30_4_lut_LC_7_14_6 .C_ON=1'b0;
    defparam \ADC_VAC1.i30_4_lut_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i30_4_lut_LC_7_14_6 .LUT_INIT=16'b1011000110000001;
    LogicCell40 \ADC_VAC1.i30_4_lut_LC_7_14_6  (
            .in0(N__30659),
            .in1(N__20631),
            .in2(N__20581),
            .in3(N__19657),
            .lcout(),
            .ltout(\ADC_VAC1.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.i13056_2_lut_LC_7_14_7 .C_ON=1'b0;
    defparam \ADC_VAC1.i13056_2_lut_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC1.i13056_2_lut_LC_7_14_7 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \ADC_VAC1.i13056_2_lut_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19607),
            .in3(N__52618),
            .lcout(\ADC_VAC1.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i15_LC_7_15_3 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i15_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i15_LC_7_15_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i15_LC_7_15_3  (
            .in0(N__26089),
            .in1(N__19782),
            .in2(N__52778),
            .in3(N__21723),
            .lcout(cmd_rdadctmp_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51278),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i14_LC_7_15_4 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i14_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i14_LC_7_15_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i14_LC_7_15_4  (
            .in0(N__19591),
            .in1(N__52679),
            .in2(N__21727),
            .in3(N__26088),
            .lcout(cmd_rdadctmp_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51278),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i1_LC_7_15_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i1_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i1_LC_7_15_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i1_LC_7_15_7  (
            .in0(N__19805),
            .in1(N__27460),
            .in2(N__19846),
            .in3(N__26858),
            .lcout(cmd_rdadctmp_1_adj_1148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51278),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i0_LC_7_16_1 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i0_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i0_LC_7_16_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i0_LC_7_16_1  (
            .in0(N__19804),
            .in1(N__27468),
            .in2(N__19829),
            .in3(N__26797),
            .lcout(cmd_rdadctmp_0_adj_1149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51291),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i16_LC_7_16_6 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i16_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i16_LC_7_16_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i16_LC_7_16_6  (
            .in0(N__19783),
            .in1(N__26127),
            .in2(N__32166),
            .in3(N__52774),
            .lcout(cmd_rdadctmp_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51291),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i17_LC_7_17_2 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i17_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i17_LC_7_17_2 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i17_LC_7_17_2  (
            .in0(N__20458),
            .in1(N__46062),
            .in2(N__46227),
            .in3(N__53402),
            .lcout(cmd_rdadctmp_17_adj_1059),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51301),
            .ce(),
            .sr(_gnd_net_));
    defparam ICE_GPMO_0_I_0_1_lut_LC_7_18_2.C_ON=1'b0;
    defparam ICE_GPMO_0_I_0_1_lut_LC_7_18_2.SEQ_MODE=4'b0000;
    defparam ICE_GPMO_0_I_0_1_lut_LC_7_18_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 ICE_GPMO_0_I_0_1_lut_LC_7_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32771),
            .lcout(M_START),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i1_7348_7349_reset_LC_8_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_7348_7349_reset_LC_8_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i1_7348_7349_reset_LC_8_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_7348_7349_reset_LC_8_4_0  (
            .in0(N__20924),
            .in1(N__20912),
            .in2(_gnd_net_),
            .in3(N__21617),
            .lcout(\comm_spi.n10460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42466),
            .ce(),
            .sr(N__20885));
    defparam comm_tx_buf_i0_LC_8_5_2.C_ON=1'b0;
    defparam comm_tx_buf_i0_LC_8_5_2.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i0_LC_8_5_2.LUT_INIT=16'b0010001011100010;
    LogicCell40 comm_tx_buf_i0_LC_8_5_2 (
            .in0(N__20837),
            .in1(N__33520),
            .in2(N__20990),
            .in3(N__33353),
            .lcout(comm_tx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51119),
            .ce(N__43134),
            .sr(N__22394));
    defparam i12201_3_lut_LC_8_5_5.C_ON=1'b0;
    defparam i12201_3_lut_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam i12201_3_lut_LC_8_5_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12201_3_lut_LC_8_5_5 (
            .in0(N__25043),
            .in1(N__23615),
            .in2(_gnd_net_),
            .in3(N__38846),
            .lcout(n15411),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12181_3_lut_LC_8_5_7.C_ON=1'b0;
    defparam i12181_3_lut_LC_8_5_7.SEQ_MODE=4'b0000;
    defparam i12181_3_lut_LC_8_5_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12181_3_lut_LC_8_5_7 (
            .in0(N__19748),
            .in1(N__19739),
            .in2(_gnd_net_),
            .in3(N__38847),
            .lcout(n15391),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16410_bdd_4_lut_LC_8_6_0.C_ON=1'b0;
    defparam n16410_bdd_4_lut_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam n16410_bdd_4_lut_LC_8_6_0.LUT_INIT=16'b1110111001010000;
    LogicCell40 n16410_bdd_4_lut_LC_8_6_0 (
            .in0(N__33106),
            .in1(N__33970),
            .in2(N__41897),
            .in3(N__19886),
            .lcout(),
            .ltout(n16413_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10400_3_lut_LC_8_6_1.C_ON=1'b0;
    defparam i10400_3_lut_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam i10400_3_lut_LC_8_6_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 i10400_3_lut_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(N__19880),
            .in2(N__19931),
            .in3(N__33349),
            .lcout(n13493),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_LC_8_6_2.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_LC_8_6_2.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_index_0__bdd_4_lut_LC_8_6_2 (
            .in0(N__38810),
            .in1(N__22229),
            .in2(N__33168),
            .in3(N__23567),
            .lcout(),
            .ltout(n16518_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16518_bdd_4_lut_LC_8_6_3.C_ON=1'b0;
    defparam n16518_bdd_4_lut_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam n16518_bdd_4_lut_LC_8_6_3.LUT_INIT=16'b1110001111100000;
    LogicCell40 n16518_bdd_4_lut_LC_8_6_3 (
            .in0(N__19928),
            .in1(N__33110),
            .in2(N__19919),
            .in3(N__20135),
            .lcout(),
            .ltout(n16521_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i6_LC_8_6_4.C_ON=1'b0;
    defparam comm_tx_buf_i6_LC_8_6_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i6_LC_8_6_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_tx_buf_i6_LC_8_6_4 (
            .in0(N__33350),
            .in1(N__19916),
            .in2(N__19910),
            .in3(N__33531),
            .lcout(comm_tx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51127),
            .ce(N__43122),
            .sr(N__22383));
    defparam comm_index_0__bdd_4_lut_13200_LC_8_6_5.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13200_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13200_LC_8_6_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13200_LC_8_6_5 (
            .in0(N__19907),
            .in1(N__33104),
            .in2(N__19895),
            .in3(N__38809),
            .lcout(n16410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16488_bdd_4_lut_LC_8_6_6.C_ON=1'b0;
    defparam n16488_bdd_4_lut_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam n16488_bdd_4_lut_LC_8_6_6.LUT_INIT=16'b1111101001000100;
    LogicCell40 n16488_bdd_4_lut_LC_8_6_6 (
            .in0(N__33105),
            .in1(N__23369),
            .in2(N__24794),
            .in3(N__25127),
            .lcout(n16491),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13195_LC_8_7_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13195_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13195_LC_8_7_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13195_LC_8_7_0 (
            .in0(N__19874),
            .in1(N__33182),
            .in2(N__19862),
            .in3(N__38839),
            .lcout(),
            .ltout(n16404_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16404_bdd_4_lut_LC_8_7_1.C_ON=1'b0;
    defparam n16404_bdd_4_lut_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam n16404_bdd_4_lut_LC_8_7_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16404_bdd_4_lut_LC_8_7_1 (
            .in0(N__33183),
            .in1(N__34560),
            .in2(N__19850),
            .in3(N__41105),
            .lcout(),
            .ltout(n16407_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i979126_i1_3_lut_LC_8_7_2.C_ON=1'b0;
    defparam i979126_i1_3_lut_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam i979126_i1_3_lut_LC_8_7_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 i979126_i1_3_lut_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__19976),
            .in2(N__20006),
            .in3(N__33524),
            .lcout(n7_adj_1240),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16512_bdd_4_lut_LC_8_7_3.C_ON=1'b0;
    defparam n16512_bdd_4_lut_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam n16512_bdd_4_lut_LC_8_7_3.LUT_INIT=16'b1110111001010000;
    LogicCell40 n16512_bdd_4_lut_LC_8_7_3 (
            .in0(N__33181),
            .in1(N__20003),
            .in2(N__19991),
            .in3(N__19970),
            .lcout(n16515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13284_LC_8_7_4.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13284_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13284_LC_8_7_4.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13284_LC_8_7_4 (
            .in0(N__23774),
            .in1(N__33180),
            .in2(N__22091),
            .in3(N__38838),
            .lcout(n16512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16422_bdd_4_lut_LC_8_7_5.C_ON=1'b0;
    defparam n16422_bdd_4_lut_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam n16422_bdd_4_lut_LC_8_7_5.LUT_INIT=16'b1111101001000100;
    LogicCell40 n16422_bdd_4_lut_LC_8_7_5 (
            .in0(N__33184),
            .in1(N__23645),
            .in2(N__24707),
            .in3(N__24980),
            .lcout(),
            .ltout(n16425_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i1_LC_8_7_6.C_ON=1'b0;
    defparam comm_tx_buf_i1_LC_8_7_6.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i1_LC_8_7_6.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_tx_buf_i1_LC_8_7_6 (
            .in0(N__33351),
            .in1(N__19964),
            .in2(N__19958),
            .in3(N__33525),
            .lcout(comm_tx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51139),
            .ce(N__43138),
            .sr(N__22392));
    defparam \comm_spi.data_tx_i7_7337_7338_set_LC_8_8_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_7337_7338_set_LC_8_8_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i7_7337_7338_set_LC_8_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_7337_7338_set_LC_8_8_0  (
            .in0(N__27668),
            .in1(N__27794),
            .in2(_gnd_net_),
            .in3(N__28994),
            .lcout(\comm_spi.n10448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42467),
            .ce(),
            .sr(N__30779));
    defparam i1_2_lut_adj_60_LC_8_8_1.C_ON=1'b0;
    defparam i1_2_lut_adj_60_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_60_LC_8_8_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_60_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__36587),
            .in2(_gnd_net_),
            .in3(N__33566),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1457_i5_4_lut_LC_8_9_0.C_ON=1'b0;
    defparam mux_1457_i5_4_lut_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam mux_1457_i5_4_lut_LC_8_9_0.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1457_i5_4_lut_LC_8_9_0 (
            .in0(N__19955),
            .in1(N__48035),
            .in2(N__20491),
            .in3(N__47291),
            .lcout(),
            .ltout(n4060_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i4_LC_8_9_1.C_ON=1'b0;
    defparam comm_buf_4__i4_LC_8_9_1.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i4_LC_8_9_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_4__i4_LC_8_9_1 (
            .in0(N__39932),
            .in1(_gnd_net_),
            .in2(N__19934),
            .in3(N__50325),
            .lcout(comm_buf_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51162),
            .ce(N__25449),
            .sr(N__20095));
    defparam comm_buf_4__i5_LC_8_9_3.C_ON=1'b0;
    defparam comm_buf_4__i5_LC_8_9_3.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i5_LC_8_9_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i5_LC_8_9_3 (
            .in0(N__39798),
            .in1(N__28595),
            .in2(_gnd_net_),
            .in3(N__50326),
            .lcout(comm_buf_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51162),
            .ce(N__25449),
            .sr(N__20095));
    defparam comm_buf_4__i6_LC_8_9_5.C_ON=1'b0;
    defparam comm_buf_4__i6_LC_8_9_5.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i6_LC_8_9_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i6_LC_8_9_5 (
            .in0(N__40732),
            .in1(N__20258),
            .in2(_gnd_net_),
            .in3(N__50327),
            .lcout(comm_buf_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51162),
            .ce(N__25449),
            .sr(N__20095));
    defparam mux_1457_i8_4_lut_LC_8_9_6.C_ON=1'b0;
    defparam mux_1457_i8_4_lut_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam mux_1457_i8_4_lut_LC_8_9_6.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1457_i8_4_lut_LC_8_9_6 (
            .in0(N__20126),
            .in1(N__48036),
            .in2(N__26003),
            .in3(N__47292),
            .lcout(),
            .ltout(n4057_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i7_LC_8_9_7.C_ON=1'b0;
    defparam comm_buf_4__i7_LC_8_9_7.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i7_LC_8_9_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_4__i7_LC_8_9_7 (
            .in0(N__39383),
            .in1(_gnd_net_),
            .in2(N__20105),
            .in3(N__50328),
            .lcout(comm_buf_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51162),
            .ce(N__25449),
            .sr(N__20095));
    defparam \ADC_VAC1.ADC_DATA_i17_LC_8_10_0 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i17_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i17_LC_8_10_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i17_LC_8_10_0  (
            .in0(N__53075),
            .in1(N__20056),
            .in2(N__20207),
            .in3(N__52888),
            .lcout(buf_adcdata1_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i18_LC_8_10_1 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i18_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i18_LC_8_10_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i18_LC_8_10_1  (
            .in0(N__52879),
            .in1(N__53076),
            .in2(N__20041),
            .in3(N__20020),
            .lcout(buf_adcdata1_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i26_LC_8_10_2 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i26_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i26_LC_8_10_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i26_LC_8_10_2  (
            .in0(N__20202),
            .in1(N__52883),
            .in2(N__20021),
            .in3(N__26158),
            .lcout(cmd_rdadctmp_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i27_LC_8_10_3 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i27_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i27_LC_8_10_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i27_LC_8_10_3  (
            .in0(N__26159),
            .in1(N__20247),
            .in2(N__52898),
            .in3(N__20019),
            .lcout(cmd_rdadctmp_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i28_LC_8_10_4 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i28_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i28_LC_8_10_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i28_LC_8_10_4  (
            .in0(N__20248),
            .in1(N__52884),
            .in2(N__20374),
            .in3(N__26160),
            .lcout(cmd_rdadctmp_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i19_LC_8_10_5 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i19_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i19_LC_8_10_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i19_LC_8_10_5  (
            .in0(N__52880),
            .in1(N__53077),
            .in2(N__20227),
            .in3(N__20249),
            .lcout(buf_adcdata1_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i25_LC_8_10_6 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i25_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i25_LC_8_10_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i25_LC_8_10_6  (
            .in0(N__48259),
            .in1(N__52882),
            .in2(N__20206),
            .in3(N__26157),
            .lcout(cmd_rdadctmp_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i20_LC_8_10_7 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i20_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i20_LC_8_10_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i20_LC_8_10_7  (
            .in0(N__52881),
            .in1(N__53078),
            .in2(N__20182),
            .in3(N__20370),
            .lcout(buf_adcdata1_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51180),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_140_LC_8_11_0.C_ON=1'b0;
    defparam i1_4_lut_adj_140_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_140_LC_8_11_0.LUT_INIT=16'b1111111100100001;
    LogicCell40 i1_4_lut_adj_140_LC_8_11_0 (
            .in0(N__45659),
            .in1(N__47077),
            .in2(N__39556),
            .in3(N__40884),
            .lcout(n84),
            .ltout(n84_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12632_2_lut_LC_8_11_1.C_ON=1'b0;
    defparam i12632_2_lut_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam i12632_2_lut_LC_8_11_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12632_2_lut_LC_8_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20162),
            .in3(N__34550),
            .lcout(),
            .ltout(n15593_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i1_LC_8_11_2.C_ON=1'b0;
    defparam comm_buf_0__i1_LC_8_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i1_LC_8_11_2.LUT_INIT=16'b1011101110111000;
    LogicCell40 comm_buf_0__i1_LC_8_11_2 (
            .in0(N__44178),
            .in1(N__50345),
            .in2(N__20159),
            .in3(N__26012),
            .lcout(comm_buf_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51198),
            .ce(N__25274),
            .sr(N__24209));
    defparam i1_4_lut_adj_150_LC_8_11_3.C_ON=1'b0;
    defparam i1_4_lut_adj_150_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_150_LC_8_11_3.LUT_INIT=16'b1010000010101000;
    LogicCell40 i1_4_lut_adj_150_LC_8_11_3 (
            .in0(N__40252),
            .in1(N__23867),
            .in2(N__27617),
            .in3(N__45220),
            .lcout(),
            .ltout(n8045_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i7_LC_8_11_4.C_ON=1'b0;
    defparam comm_buf_0__i7_LC_8_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i7_LC_8_11_4.LUT_INIT=16'b1111111001010100;
    LogicCell40 comm_buf_0__i7_LC_8_11_4 (
            .in0(N__50344),
            .in1(N__20153),
            .in2(N__20156),
            .in3(N__39396),
            .lcout(comm_buf_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51198),
            .ce(N__25274),
            .sr(N__24209));
    defparam i12650_2_lut_LC_8_11_5.C_ON=1'b0;
    defparam i12650_2_lut_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam i12650_2_lut_LC_8_11_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12650_2_lut_LC_8_11_5 (
            .in0(_gnd_net_),
            .in1(N__38904),
            .in2(_gnd_net_),
            .in3(N__32094),
            .lcout(n15573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i11_LC_8_12_0 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i11_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i11_LC_8_12_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i11_LC_8_12_0  (
            .in0(N__44464),
            .in1(N__52837),
            .in2(N__20518),
            .in3(N__26177),
            .lcout(cmd_rdadctmp_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51215),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i12_LC_8_12_1 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i12_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i12_LC_8_12_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i12_LC_8_12_1  (
            .in0(N__25920),
            .in1(N__20481),
            .in2(N__22666),
            .in3(N__27464),
            .lcout(buf_adcdata4_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51215),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i8_LC_8_12_2 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i8_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i8_LC_8_12_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i8_LC_8_12_2  (
            .in0(N__53697),
            .in1(N__20410),
            .in2(N__20459),
            .in3(N__53294),
            .lcout(buf_adcdata2_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51215),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i9_LC_8_12_3 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i9_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i9_LC_8_12_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i9_LC_8_12_3  (
            .in0(N__20391),
            .in1(N__49240),
            .in2(N__43840),
            .in3(N__48816),
            .lcout(cmd_rdadctmp_9_adj_1103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51215),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i29_LC_8_12_6 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i29_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i29_LC_8_12_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i29_LC_8_12_6  (
            .in0(N__20375),
            .in1(N__21288),
            .in2(N__52889),
            .in3(N__26178),
            .lcout(cmd_rdadctmp_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51215),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i9_LC_8_13_0 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i9_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i9_LC_8_13_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i9_LC_8_13_0  (
            .in0(N__24144),
            .in1(N__22476),
            .in2(N__52891),
            .in3(N__26161),
            .lcout(cmd_rdadctmp_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51232),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i17_LC_8_13_1 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i17_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i17_LC_8_13_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i17_LC_8_13_1  (
            .in0(N__53716),
            .in1(N__20344),
            .in2(N__43966),
            .in3(N__53276),
            .lcout(buf_adcdata2_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51232),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i15_LC_8_13_2 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i15_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i15_LC_8_13_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i15_LC_8_13_2  (
            .in0(N__48776),
            .in1(N__21663),
            .in2(N__49204),
            .in3(N__20292),
            .lcout(cmd_rdadctmp_15_adj_1097),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51232),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i14_LC_8_13_3 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i14_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i14_LC_8_13_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i14_LC_8_13_3  (
            .in0(N__20330),
            .in1(N__49124),
            .in2(N__20296),
            .in3(N__48777),
            .lcout(cmd_rdadctmp_14_adj_1098),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51232),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1457_i7_4_lut_LC_8_13_7.C_ON=1'b0;
    defparam mux_1457_i7_4_lut_LC_8_13_7.SEQ_MODE=4'b0000;
    defparam mux_1457_i7_4_lut_LC_8_13_7.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1457_i7_4_lut_LC_8_13_7 (
            .in0(N__20276),
            .in1(N__48074),
            .in2(N__24103),
            .in3(N__47311),
            .lcout(n4058),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_200_LC_8_14_3.C_ON=1'b0;
    defparam i1_4_lut_adj_200_LC_8_14_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_200_LC_8_14_3.LUT_INIT=16'b0000101100001110;
    LogicCell40 i1_4_lut_adj_200_LC_8_14_3 (
            .in0(N__23062),
            .in1(N__49107),
            .in2(N__20695),
            .in3(N__22978),
            .lcout(),
            .ltout(n14_adj_1031_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.CS_37_LC_8_14_4 .C_ON=1'b0;
    defparam \ADC_VAC3.CS_37_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.CS_37_LC_8_14_4 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \ADC_VAC3.CS_37_LC_8_14_4  (
            .in0(N__49108),
            .in1(N__23123),
            .in2(N__20711),
            .in3(N__20723),
            .lcout(M_CS3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51248),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i25_LC_8_14_5 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i25_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i25_LC_8_14_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i25_LC_8_14_5  (
            .in0(N__21327),
            .in1(N__46063),
            .in2(N__43962),
            .in3(N__53277),
            .lcout(cmd_rdadctmp_25_adj_1051),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51248),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i24_LC_8_15_0 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i24_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i24_LC_8_15_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i24_LC_8_15_0  (
            .in0(N__34475),
            .in1(N__46039),
            .in2(N__21331),
            .in3(N__53278),
            .lcout(cmd_rdadctmp_24_adj_1052),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51265),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.SCLK_35_LC_8_15_1 .C_ON=1'b0;
    defparam \ADC_VAC3.SCLK_35_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.SCLK_35_LC_8_15_1 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_VAC3.SCLK_35_LC_8_15_1  (
            .in0(N__49225),
            .in1(N__22979),
            .in2(N__20674),
            .in3(N__23058),
            .lcout(M_SCLK3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51265),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i2_LC_8_15_4 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i2_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i2_LC_8_15_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i2_LC_8_15_4  (
            .in0(N__20749),
            .in1(N__49226),
            .in2(N__21538),
            .in3(N__48734),
            .lcout(cmd_rdadctmp_2_adj_1110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51265),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i4_LC_8_15_5 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i4_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i4_LC_8_15_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i4_LC_8_15_5  (
            .in0(N__48733),
            .in1(N__21521),
            .in2(N__49256),
            .in3(N__20656),
            .lcout(cmd_rdadctmp_4_adj_1108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51265),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i5_LC_8_15_6 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i5_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i5_LC_8_15_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i5_LC_8_15_6  (
            .in0(N__20657),
            .in1(N__49227),
            .in2(N__24286),
            .in3(N__48735),
            .lcout(cmd_rdadctmp_5_adj_1107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51265),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.DTRIG_39_LC_8_16_0 .C_ON=1'b0;
    defparam \ADC_VAC1.DTRIG_39_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.DTRIG_39_LC_8_16_0 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \ADC_VAC1.DTRIG_39_LC_8_16_0  (
            .in0(N__20648),
            .in1(N__20585),
            .in2(N__52890),
            .in3(N__21482),
            .lcout(acadc_dtrig1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51279),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i0_LC_8_16_1 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i0_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i0_LC_8_16_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i0_LC_8_16_1  (
            .in0(N__20758),
            .in1(N__49129),
            .in2(N__20780),
            .in3(N__48678),
            .lcout(cmd_rdadctmp_0_adj_1112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51279),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i1_LC_8_16_3 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i1_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i1_LC_8_16_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i1_LC_8_16_3  (
            .in0(N__20759),
            .in1(N__49130),
            .in2(N__20750),
            .in3(N__48679),
            .lcout(cmd_rdadctmp_1_adj_1111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51279),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i13060_2_lut_LC_8_16_5 .C_ON=1'b0;
    defparam \ADC_VAC3.i13060_2_lut_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i13060_2_lut_LC_8_16_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_VAC3.i13060_2_lut_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__49128),
            .in2(_gnd_net_),
            .in3(N__22553),
            .lcout(\ADC_VAC3.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_32_LC_8_16_7.C_ON=1'b0;
    defparam i1_2_lut_adj_32_LC_8_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_32_LC_8_16_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_32_LC_8_16_7 (
            .in0(_gnd_net_),
            .in1(N__22956),
            .in2(_gnd_net_),
            .in3(N__23042),
            .lcout(n15147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.adc_state_i2_LC_8_17_1 .C_ON=1'b0;
    defparam \ADC_VAC3.adc_state_i2_LC_8_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.adc_state_i2_LC_8_17_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_VAC3.adc_state_i2_LC_8_17_1  (
            .in0(N__49122),
            .in1(N__22955),
            .in2(_gnd_net_),
            .in3(N__23040),
            .lcout(DTRIG_N_957_adj_1114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51292),
            .ce(N__20735),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.adc_state_i1_LC_8_17_3 .C_ON=1'b0;
    defparam \ADC_VAC3.adc_state_i1_LC_8_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.adc_state_i1_LC_8_17_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \ADC_VAC3.adc_state_i1_LC_8_17_3  (
            .in0(N__49121),
            .in1(N__22954),
            .in2(_gnd_net_),
            .in3(N__23041),
            .lcout(adc_state_1_adj_1079),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51292),
            .ce(N__20735),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_50_LC_8_17_5.C_ON=1'b0;
    defparam i1_2_lut_adj_50_LC_8_17_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_50_LC_8_17_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_50_LC_8_17_5 (
            .in0(_gnd_net_),
            .in1(N__22953),
            .in2(_gnd_net_),
            .in3(N__23039),
            .lcout(n15162),
            .ltout(n15162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i1_3_lut_LC_8_17_6 .C_ON=1'b0;
    defparam \ADC_VAC3.i1_3_lut_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i1_3_lut_LC_8_17_6 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \ADC_VAC3.i1_3_lut_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__23111),
            .in2(N__20714),
            .in3(N__49120),
            .lcout(n8332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_7322_7323_set_LC_9_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_7322_7323_set_LC_9_3_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i0_7322_7323_set_LC_9_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_7322_7323_set_LC_9_3_0  (
            .in0(N__28752),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n10433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42464),
            .ce(),
            .sr(N__20876));
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_9_4_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_9_4_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_98_2_lut_LC_9_4_0  (
            .in0(N__20869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46607),
            .lcout(\comm_spi.data_tx_7__N_811 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13117_4_lut_3_lut_LC_9_4_1 .C_ON=1'b0;
    defparam \comm_spi.i13117_4_lut_3_lut_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13117_4_lut_3_lut_LC_9_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.i13117_4_lut_3_lut_LC_9_4_1  (
            .in0(N__46610),
            .in1(N__20923),
            .in2(_gnd_net_),
            .in3(N__21598),
            .lcout(\comm_spi.n16911 ),
            .ltout(\comm_spi.n16911_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i1_7348_7349_set_LC_9_4_2 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_7348_7349_set_LC_9_4_2 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i1_7348_7349_set_LC_9_4_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.data_tx_i1_7348_7349_set_LC_9_4_2  (
            .in0(N__20911),
            .in1(_gnd_net_),
            .in2(N__20900),
            .in3(N__21610),
            .lcout(\comm_spi.n10459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42465),
            .ce(),
            .sr(N__20897));
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_9_4_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_9_4_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_106_2_lut_LC_9_4_3  (
            .in0(N__46606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20868),
            .lcout(\comm_spi.data_tx_7__N_831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_9_4_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_9_4_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_99_2_lut_LC_9_4_5  (
            .in0(N__46608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21597),
            .lcout(\comm_spi.data_tx_7__N_812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13082_4_lut_3_lut_LC_9_4_6 .C_ON=1'b0;
    defparam \comm_spi.i13082_4_lut_3_lut_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13082_4_lut_3_lut_LC_9_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i13082_4_lut_3_lut_LC_9_4_6  (
            .in0(N__20870),
            .in1(N__23235),
            .in2(_gnd_net_),
            .in3(N__46609),
            .lcout(\comm_spi.n16908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_13249_LC_9_5_1.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_13249_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_13249_LC_9_5_1.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_1__bdd_4_lut_13249_LC_9_5_1 (
            .in0(N__20852),
            .in1(N__33330),
            .in2(N__20969),
            .in3(N__33176),
            .lcout(),
            .ltout(n16446_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16446_bdd_4_lut_LC_9_5_2.C_ON=1'b0;
    defparam n16446_bdd_4_lut_LC_9_5_2.SEQ_MODE=4'b0000;
    defparam n16446_bdd_4_lut_LC_9_5_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16446_bdd_4_lut_LC_9_5_2 (
            .in0(N__33331),
            .in1(N__29102),
            .in2(N__20846),
            .in3(N__20843),
            .lcout(n16449),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1525_i4_4_lut_LC_9_5_3.C_ON=1'b0;
    defparam mux_1525_i4_4_lut_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam mux_1525_i4_4_lut_LC_9_5_3.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1525_i4_4_lut_LC_9_5_3 (
            .in0(N__20831),
            .in1(N__48012),
            .in2(N__20818),
            .in3(N__47337),
            .lcout(n4305),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16428_bdd_4_lut_LC_9_5_4.C_ON=1'b0;
    defparam n16428_bdd_4_lut_LC_9_5_4.SEQ_MODE=4'b0000;
    defparam n16428_bdd_4_lut_LC_9_5_4.LUT_INIT=16'b1110111001010000;
    LogicCell40 n16428_bdd_4_lut_LC_9_5_4 (
            .in0(N__33175),
            .in1(N__24737),
            .in2(N__23261),
            .in3(N__21572),
            .lcout(n16431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13279_LC_9_6_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13279_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13279_LC_9_6_0.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_0__bdd_4_lut_13279_LC_9_6_0 (
            .in0(N__38825),
            .in1(N__23801),
            .in2(N__21860),
            .in3(N__33173),
            .lcout(),
            .ltout(n16506_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16506_bdd_4_lut_LC_9_6_1.C_ON=1'b0;
    defparam n16506_bdd_4_lut_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam n16506_bdd_4_lut_LC_9_6_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16506_bdd_4_lut_LC_9_6_1 (
            .in0(N__33174),
            .in1(N__21017),
            .in2(N__21005),
            .in3(N__21002),
            .lcout(n16509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12214_3_lut_LC_9_6_2.C_ON=1'b0;
    defparam i12214_3_lut_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam i12214_3_lut_LC_9_6_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12214_3_lut_LC_9_6_2 (
            .in0(N__38823),
            .in1(N__22151),
            .in2(_gnd_net_),
            .in3(N__23486),
            .lcout(n15424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12202_3_lut_LC_9_6_3.C_ON=1'b0;
    defparam i12202_3_lut_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam i12202_3_lut_LC_9_6_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12202_3_lut_LC_9_6_3 (
            .in0(N__21914),
            .in1(N__23894),
            .in2(_gnd_net_),
            .in3(N__38821),
            .lcout(n15412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12240_3_lut_LC_9_6_4.C_ON=1'b0;
    defparam i12240_3_lut_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam i12240_3_lut_LC_9_6_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12240_3_lut_LC_9_6_4 (
            .in0(N__38822),
            .in1(N__20960),
            .in2(_gnd_net_),
            .in3(N__20951),
            .lcout(n15450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13259_LC_9_6_6.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13259_LC_9_6_6.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13259_LC_9_6_6.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_0__bdd_4_lut_13259_LC_9_6_6 (
            .in0(N__38824),
            .in1(N__25370),
            .in2(N__21983),
            .in3(N__33171),
            .lcout(),
            .ltout(n16482_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16482_bdd_4_lut_LC_9_6_7.C_ON=1'b0;
    defparam n16482_bdd_4_lut_LC_9_6_7.SEQ_MODE=4'b0000;
    defparam n16482_bdd_4_lut_LC_9_6_7.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16482_bdd_4_lut_LC_9_6_7 (
            .in0(N__33172),
            .in1(N__23342),
            .in2(N__20939),
            .in3(N__24824),
            .lcout(n16485),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imiso_83_7340_7341_reset_LC_9_7_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_7340_7341_reset_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imiso_83_7340_7341_reset_LC_9_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.imiso_83_7340_7341_reset_LC_9_7_0  (
            .in0(N__29128),
            .in1(N__29156),
            .in2(_gnd_net_),
            .in3(N__30845),
            .lcout(\comm_spi.n10452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_7340_7341_resetC_net ),
            .ce(),
            .sr(N__31007));
    defparam comm_buf_3__i2_LC_9_8_0.C_ON=1'b0;
    defparam comm_buf_3__i2_LC_9_8_0.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i2_LC_9_8_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i2_LC_9_8_0 (
            .in0(N__40121),
            .in1(N__21137),
            .in2(_gnd_net_),
            .in3(N__49896),
            .lcout(comm_buf_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51140),
            .ce(N__25175),
            .sr(N__30736));
    defparam comm_buf_3__i3_LC_9_8_1.C_ON=1'b0;
    defparam comm_buf_3__i3_LC_9_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i3_LC_9_8_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i3_LC_9_8_1 (
            .in0(N__49895),
            .in1(N__44909),
            .in2(_gnd_net_),
            .in3(N__43001),
            .lcout(comm_buf_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51140),
            .ce(N__25175),
            .sr(N__30736));
    defparam comm_buf_9__i3_LC_9_9_0.C_ON=1'b0;
    defparam comm_buf_9__i3_LC_9_9_0.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i3_LC_9_9_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_9__i3_LC_9_9_0 (
            .in0(N__44910),
            .in1(N__21104),
            .in2(_gnd_net_),
            .in3(N__50330),
            .lcout(comm_buf_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51150),
            .ce(N__27707),
            .sr(N__30743));
    defparam comm_buf_9__i4_LC_9_9_1.C_ON=1'b0;
    defparam comm_buf_9__i4_LC_9_9_1.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i4_LC_9_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_9__i4_LC_9_9_1 (
            .in0(N__50329),
            .in1(N__39940),
            .in2(_gnd_net_),
            .in3(N__21077),
            .lcout(comm_buf_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51150),
            .ce(N__27707),
            .sr(N__30743));
    defparam i132_4_lut_adj_100_LC_9_10_0.C_ON=1'b0;
    defparam i132_4_lut_adj_100_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam i132_4_lut_adj_100_LC_9_10_0.LUT_INIT=16'b0101100000001000;
    LogicCell40 i132_4_lut_adj_100_LC_9_10_0 (
            .in0(N__48041),
            .in1(N__41258),
            .in2(N__45317),
            .in3(N__29581),
            .lcout(),
            .ltout(n66_adj_1153_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i123_3_lut_adj_105_LC_9_10_1.C_ON=1'b0;
    defparam i123_3_lut_adj_105_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam i123_3_lut_adj_105_LC_9_10_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 i123_3_lut_adj_105_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(N__29300),
            .in2(N__21062),
            .in3(N__47268),
            .lcout(n96_adj_1159),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12672_2_lut_LC_9_10_2.C_ON=1'b0;
    defparam i12672_2_lut_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam i12672_2_lut_LC_9_10_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12672_2_lut_LC_9_10_2 (
            .in0(N__32104),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33752),
            .lcout(n15578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i20_LC_9_10_3 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i20_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i20_LC_9_10_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i20_LC_9_10_3  (
            .in0(N__44351),
            .in1(N__49123),
            .in2(N__24251),
            .in3(N__24060),
            .lcout(buf_adcdata3_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51163),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.SCLK_27_LC_9_10_4 .C_ON=1'b0;
    defparam \CLOCK_DDS.SCLK_27_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.SCLK_27_LC_9_10_4 .LUT_INIT=16'b0101010011010001;
    LogicCell40 \CLOCK_DDS.SCLK_27_LC_9_10_4  (
            .in0(N__35765),
            .in1(N__48363),
            .in2(N__21046),
            .in3(N__48544),
            .lcout(DDS_SCK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51163),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.MOSI_31_LC_9_10_6 .C_ON=1'b0;
    defparam \CLOCK_DDS.MOSI_31_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.MOSI_31_LC_9_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CLOCK_DDS.MOSI_31_LC_9_10_6  (
            .in0(N__31046),
            .in1(N__21214),
            .in2(_gnd_net_),
            .in3(N__48543),
            .lcout(DDS_MOSI1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51163),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.bit_cnt_i0_LC_9_10_7 .C_ON=1'b0;
    defparam \CLOCK_DDS.bit_cnt_i0_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.bit_cnt_i0_LC_9_10_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \CLOCK_DDS.bit_cnt_i0_LC_9_10_7  (
            .in0(N__48545),
            .in1(N__25495),
            .in2(_gnd_net_),
            .in3(N__31189),
            .lcout(bit_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51163),
            .ce(),
            .sr(_gnd_net_));
    defparam i12726_2_lut_LC_9_11_0.C_ON=1'b0;
    defparam i12726_2_lut_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam i12726_2_lut_LC_9_11_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12726_2_lut_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(N__48040),
            .in2(_gnd_net_),
            .in3(N__32216),
            .lcout(n15522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12666_2_lut_LC_9_11_1.C_ON=1'b0;
    defparam i12666_2_lut_LC_9_11_1.SEQ_MODE=4'b0000;
    defparam i12666_2_lut_LC_9_11_1.LUT_INIT=16'b0000000010101010;
    LogicCell40 i12666_2_lut_LC_9_11_1 (
            .in0(N__31430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48042),
            .lcout(n15523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_13215_LC_9_11_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_13215_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_13215_LC_9_11_2.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_13215_LC_9_11_2 (
            .in0(N__45219),
            .in1(N__21203),
            .in2(N__21197),
            .in3(N__47260),
            .lcout(),
            .ltout(n16398_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16398_bdd_4_lut_LC_9_11_3.C_ON=1'b0;
    defparam n16398_bdd_4_lut_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam n16398_bdd_4_lut_LC_9_11_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16398_bdd_4_lut_LC_9_11_3 (
            .in0(N__47261),
            .in1(N__34046),
            .in2(N__21188),
            .in3(N__27749),
            .lcout(),
            .ltout(n16401_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i108_4_lut_LC_9_11_4.C_ON=1'b0;
    defparam i108_4_lut_LC_9_11_4.SEQ_MODE=4'b0000;
    defparam i108_4_lut_LC_9_11_4.LUT_INIT=16'b1101100001010000;
    LogicCell40 i108_4_lut_LC_9_11_4 (
            .in0(N__45660),
            .in1(N__34253),
            .in2(N__21185),
            .in3(N__47262),
            .lcout(),
            .ltout(n109_adj_1155_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_123_LC_9_11_5.C_ON=1'b0;
    defparam i1_4_lut_adj_123_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_123_LC_9_11_5.LUT_INIT=16'b1111001000000000;
    LogicCell40 i1_4_lut_adj_123_LC_9_11_5 (
            .in0(N__31292),
            .in1(N__39543),
            .in2(N__21182),
            .in3(N__40251),
            .lcout(),
            .ltout(n8048_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i5_LC_9_11_6.C_ON=1'b0;
    defparam comm_buf_0__i5_LC_9_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i5_LC_9_11_6.LUT_INIT=16'b1011101110111000;
    LogicCell40 comm_buf_0__i5_LC_9_11_6 (
            .in0(N__39808),
            .in1(N__50323),
            .in2(N__21179),
            .in3(N__21176),
            .lcout(comm_buf_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51181),
            .ce(N__25269),
            .sr(N__24205));
    defparam \ADC_VAC1.ADC_DATA_i21_LC_9_12_0 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i21_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i21_LC_9_12_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i21_LC_9_12_0  (
            .in0(N__52831),
            .in1(N__53127),
            .in2(N__21157),
            .in3(N__21290),
            .lcout(buf_adcdata1_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51199),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i22_LC_9_12_1 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i22_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i22_LC_9_12_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i22_LC_9_12_1  (
            .in0(N__53126),
            .in1(N__52834),
            .in2(N__21355),
            .in3(N__21274),
            .lcout(buf_adcdata1_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51199),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i16_LC_9_12_2 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i16_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i16_LC_9_12_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i16_LC_9_12_2  (
            .in0(N__53698),
            .in1(N__21304),
            .in2(N__21335),
            .in3(N__53293),
            .lcout(buf_adcdata2_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51199),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i31_LC_9_12_3 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i31_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i31_LC_9_12_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i31_LC_9_12_3  (
            .in0(N__26180),
            .in1(N__21273),
            .in2(N__22753),
            .in3(N__52835),
            .lcout(cmd_rdadctmp_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51199),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i30_LC_9_12_4 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i30_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i30_LC_9_12_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i30_LC_9_12_4  (
            .in0(N__52832),
            .in1(N__21289),
            .in2(N__21275),
            .in3(N__26179),
            .lcout(cmd_rdadctmp_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51199),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i1_LC_9_12_7 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i1_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i1_LC_9_12_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i1_LC_9_12_7  (
            .in0(N__53125),
            .in1(N__21250),
            .in2(N__24154),
            .in3(N__52833),
            .lcout(buf_adcdata1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51199),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.bit_cnt_i0_LC_9_13_0 .C_ON=1'b1;
    defparam \ADC_VAC2.bit_cnt_i0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i0_LC_9_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i0_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__21383),
            .in2(_gnd_net_),
            .in3(N__21236),
            .lcout(\ADC_VAC2.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\ADC_VAC2.n13988 ),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.bit_cnt_i1_LC_9_13_1 .C_ON=1'b1;
    defparam \ADC_VAC2.bit_cnt_i1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i1_LC_9_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i1_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__21439),
            .in2(_gnd_net_),
            .in3(N__21233),
            .lcout(\ADC_VAC2.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC2.n13988 ),
            .carryout(\ADC_VAC2.n13989 ),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.bit_cnt_i2_LC_9_13_2 .C_ON=1'b1;
    defparam \ADC_VAC2.bit_cnt_i2_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i2_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i2_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__22601),
            .in2(_gnd_net_),
            .in3(N__21230),
            .lcout(\ADC_VAC2.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC2.n13989 ),
            .carryout(\ADC_VAC2.n13990 ),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.bit_cnt_i3_LC_9_13_3 .C_ON=1'b1;
    defparam \ADC_VAC2.bit_cnt_i3_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i3_LC_9_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i3_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__22628),
            .in2(_gnd_net_),
            .in3(N__21227),
            .lcout(\ADC_VAC2.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC2.n13990 ),
            .carryout(\ADC_VAC2.n13991 ),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.bit_cnt_i4_LC_9_13_4 .C_ON=1'b1;
    defparam \ADC_VAC2.bit_cnt_i4_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i4_LC_9_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i4_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__22640),
            .in2(_gnd_net_),
            .in3(N__21452),
            .lcout(\ADC_VAC2.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC2.n13991 ),
            .carryout(\ADC_VAC2.n13992 ),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.bit_cnt_i5_LC_9_13_5 .C_ON=1'b1;
    defparam \ADC_VAC2.bit_cnt_i5_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i5_LC_9_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i5_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__22615),
            .in2(_gnd_net_),
            .in3(N__21449),
            .lcout(\ADC_VAC2.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC2.n13992 ),
            .carryout(\ADC_VAC2.n13993 ),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.bit_cnt_i6_LC_9_13_6 .C_ON=1'b1;
    defparam \ADC_VAC2.bit_cnt_i6_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i6_LC_9_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i6_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__21397),
            .in2(_gnd_net_),
            .in3(N__21446),
            .lcout(\ADC_VAC2.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC2.n13993 ),
            .carryout(\ADC_VAC2.n13994 ),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.bit_cnt_i7_LC_9_13_7 .C_ON=1'b0;
    defparam \ADC_VAC2.bit_cnt_i7_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.bit_cnt_i7_LC_9_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC2.bit_cnt_i7_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__21427),
            .in2(_gnd_net_),
            .in3(N__21443),
            .lcout(\ADC_VAC2.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51216),
            .ce(N__36505),
            .sr(N__36377));
    defparam \ADC_VAC2.i12780_4_lut_LC_9_14_0 .C_ON=1'b0;
    defparam \ADC_VAC2.i12780_4_lut_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i12780_4_lut_LC_9_14_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \ADC_VAC2.i12780_4_lut_LC_9_14_0  (
            .in0(N__21440),
            .in1(N__21371),
            .in2(N__21428),
            .in3(N__22589),
            .lcout(\ADC_VAC2.n15595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i1_4_lut_adj_5_LC_9_14_1 .C_ON=1'b0;
    defparam \ADC_VAC2.i1_4_lut_adj_5_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i1_4_lut_adj_5_LC_9_14_1 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_VAC2.i1_4_lut_adj_5_LC_9_14_1  (
            .in0(N__36456),
            .in1(N__53222),
            .in2(N__30214),
            .in3(N__30656),
            .lcout(),
            .ltout(\ADC_VAC2.n15261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i1_2_lut_LC_9_14_2 .C_ON=1'b0;
    defparam \ADC_VAC2.i1_2_lut_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i1_2_lut_LC_9_14_2 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \ADC_VAC2.i1_2_lut_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21413),
            .in3(N__35598),
            .lcout(\ADC_VAC2.n15262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.adc_state_i0_LC_9_14_3 .C_ON=1'b0;
    defparam \ADC_VAC2.adc_state_i0_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.adc_state_i0_LC_9_14_3 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \ADC_VAC2.adc_state_i0_LC_9_14_3  (
            .in0(N__35599),
            .in1(N__53223),
            .in2(N__36470),
            .in3(N__21410),
            .lcout(adc_state_0_adj_1044),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51233),
            .ce(N__21404),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i6_4_lut_LC_9_14_4 .C_ON=1'b0;
    defparam \ADC_VAC2.i6_4_lut_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i6_4_lut_LC_9_14_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \ADC_VAC2.i6_4_lut_LC_9_14_4  (
            .in0(N__53221),
            .in1(N__35595),
            .in2(N__21398),
            .in3(N__21382),
            .lcout(\ADC_VAC2.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i30_4_lut_LC_9_14_5 .C_ON=1'b0;
    defparam \ADC_VAC2.i30_4_lut_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i30_4_lut_LC_9_14_5 .LUT_INIT=16'b1010100000110001;
    LogicCell40 \ADC_VAC2.i30_4_lut_LC_9_14_5  (
            .in0(N__35597),
            .in1(N__36434),
            .in2(N__30215),
            .in3(N__30657),
            .lcout(),
            .ltout(\ADC_VAC2.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i13058_2_lut_LC_9_14_6 .C_ON=1'b0;
    defparam \ADC_VAC2.i13058_2_lut_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i13058_2_lut_LC_9_14_6 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \ADC_VAC2.i13058_2_lut_LC_9_14_6  (
            .in0(N__53220),
            .in1(_gnd_net_),
            .in2(N__21542),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC2.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i1_4_lut_LC_9_14_7 .C_ON=1'b0;
    defparam \ADC_VAC2.i1_4_lut_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i1_4_lut_LC_9_14_7 .LUT_INIT=16'b0000000001000110;
    LogicCell40 \ADC_VAC2.i1_4_lut_LC_9_14_7  (
            .in0(N__35596),
            .in1(N__36433),
            .in2(N__30213),
            .in3(N__53219),
            .lcout(\ADC_VAC2.n9413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i1_2_lut_LC_9_15_1 .C_ON=1'b0;
    defparam \ADC_VAC3.i1_2_lut_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i1_2_lut_LC_9_15_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \ADC_VAC3.i1_2_lut_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__23057),
            .in2(_gnd_net_),
            .in3(N__22559),
            .lcout(\ADC_VAC3.n15260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.DTRIG_39_LC_9_15_4 .C_ON=1'b0;
    defparam \ADC_VAC2.DTRIG_39_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.DTRIG_39_LC_9_15_4 .LUT_INIT=16'b1111010011100000;
    LogicCell40 \ADC_VAC2.DTRIG_39_LC_9_15_4  (
            .in0(N__53275),
            .in1(N__35568),
            .in2(N__21502),
            .in3(N__36474),
            .lcout(acadc_dtrig2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51249),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i3_LC_9_15_7 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i3_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i3_LC_9_15_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i3_LC_9_15_7  (
            .in0(N__21539),
            .in1(N__49012),
            .in2(N__21520),
            .in3(N__48757),
            .lcout(cmd_rdadctmp_3_adj_1109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51249),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_127_LC_9_16_0.C_ON=1'b0;
    defparam i3_4_lut_adj_127_LC_9_16_0.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_127_LC_9_16_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i3_4_lut_adj_127_LC_9_16_0 (
            .in0(N__21460),
            .in1(N__21469),
            .in2(N__21503),
            .in3(N__21481),
            .lcout(n14087),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.DTRIG_39_LC_9_16_1 .C_ON=1'b0;
    defparam \ADC_VAC4.DTRIG_39_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.DTRIG_39_LC_9_16_1 .LUT_INIT=16'b1010111010101000;
    LogicCell40 \ADC_VAC4.DTRIG_39_LC_9_16_1  (
            .in0(N__21470),
            .in1(N__27115),
            .in2(N__27467),
            .in3(N__27034),
            .lcout(acadc_dtrig4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51266),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.DTRIG_39_LC_9_16_4 .C_ON=1'b0;
    defparam \ADC_VAC3.DTRIG_39_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.DTRIG_39_LC_9_16_4 .LUT_INIT=16'b1011101010101000;
    LogicCell40 \ADC_VAC3.DTRIG_39_LC_9_16_4  (
            .in0(N__21461),
            .in1(N__49231),
            .in2(N__22980),
            .in3(N__23049),
            .lcout(acadc_dtrig3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51266),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i6_LC_9_16_7 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i6_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i6_LC_9_16_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i6_LC_9_16_7  (
            .in0(N__53063),
            .in1(N__21694),
            .in2(N__21734),
            .in3(N__52846),
            .lcout(buf_adcdata1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51266),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i18_LC_9_17_0 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i18_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i18_LC_9_17_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i18_LC_9_17_0  (
            .in0(N__46228),
            .in1(N__46072),
            .in2(N__38283),
            .in3(N__53325),
            .lcout(cmd_rdadctmp_18_adj_1058),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51280),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i16_LC_9_17_3 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i16_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i16_LC_9_17_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i16_LC_9_17_3  (
            .in0(N__21676),
            .in1(N__49029),
            .in2(N__38193),
            .in3(N__48680),
            .lcout(cmd_rdadctmp_16_adj_1096),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51280),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.SCLK_35_LC_9_17_5 .C_ON=1'b0;
    defparam \ADC_VAC4.SCLK_35_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.SCLK_35_LC_9_17_5 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_VAC4.SCLK_35_LC_9_17_5  (
            .in0(N__27336),
            .in1(N__27116),
            .in2(N__21634),
            .in3(N__27035),
            .lcout(M_SCLK4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51280),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_7322_7323_reset_LC_10_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_7322_7323_reset_LC_10_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i0_7322_7323_reset_LC_10_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_7322_7323_reset_LC_10_3_0  (
            .in0(N__28751),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n10434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42463),
            .ce(),
            .sr(N__21581));
    defparam \comm_spi.data_tx_i2_7352_7353_set_LC_10_4_4 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_7352_7353_set_LC_10_4_4 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i2_7352_7353_set_LC_10_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_7352_7353_set_LC_10_4_4  (
            .in0(N__23236),
            .in1(N__23215),
            .in2(_gnd_net_),
            .in3(N__23200),
            .lcout(\comm_spi.n10463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42448),
            .ce(),
            .sr(N__24905));
    defparam \comm_spi.RESET_I_0_2_lut_LC_10_5_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_2_lut_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_2_lut_LC_10_5_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_2_lut_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__21599),
            .in2(_gnd_net_),
            .in3(N__46605),
            .lcout(\comm_spi.data_tx_7__N_834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13220_LC_10_5_1.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13220_LC_10_5_1.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13220_LC_10_5_1.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13220_LC_10_5_1 (
            .in0(N__23705),
            .in1(N__33170),
            .in2(N__21746),
            .in3(N__38837),
            .lcout(n16428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1469_i5_4_lut_LC_10_5_3.C_ON=1'b0;
    defparam mux_1469_i5_4_lut_LC_10_5_3.SEQ_MODE=4'b0000;
    defparam mux_1469_i5_4_lut_LC_10_5_3.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1469_i5_4_lut_LC_10_5_3 (
            .in0(N__21566),
            .in1(N__48083),
            .in2(N__24652),
            .in3(N__47293),
            .lcout(n4104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12172_3_lut_LC_10_6_0.C_ON=1'b0;
    defparam i12172_3_lut_LC_10_6_0.SEQ_MODE=4'b0000;
    defparam i12172_3_lut_LC_10_6_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12172_3_lut_LC_10_6_0 (
            .in0(N__21827),
            .in1(N__21818),
            .in2(_gnd_net_),
            .in3(N__38828),
            .lcout(),
            .ltout(n15382_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16380_bdd_4_lut_LC_10_6_1.C_ON=1'b0;
    defparam n16380_bdd_4_lut_LC_10_6_1.SEQ_MODE=4'b0000;
    defparam n16380_bdd_4_lut_LC_10_6_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 n16380_bdd_4_lut_LC_10_6_1 (
            .in0(N__38582),
            .in1(N__21782),
            .in2(N__21806),
            .in3(N__33490),
            .lcout(),
            .ltout(n16383_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i7_LC_10_6_2.C_ON=1'b0;
    defparam comm_tx_buf_i7_LC_10_6_2.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i7_LC_10_6_2.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_tx_buf_i7_LC_10_6_2 (
            .in0(N__33491),
            .in1(N__21797),
            .in2(N__21803),
            .in3(N__33346),
            .lcout(comm_tx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51114),
            .ce(N__43139),
            .sr(N__22384));
    defparam comm_index_0__bdd_4_lut_13274_LC_10_6_4.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13274_LC_10_6_4.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13274_LC_10_6_4.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13274_LC_10_6_4 (
            .in0(N__33130),
            .in1(N__23930),
            .in2(N__21944),
            .in3(N__38827),
            .lcout(),
            .ltout(n16494_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16494_bdd_4_lut_LC_10_6_5.C_ON=1'b0;
    defparam n16494_bdd_4_lut_LC_10_6_5.SEQ_MODE=4'b0000;
    defparam n16494_bdd_4_lut_LC_10_6_5.LUT_INIT=16'b1110001111100000;
    LogicCell40 n16494_bdd_4_lut_LC_10_6_5 (
            .in0(N__24764),
            .in1(N__33132),
            .in2(N__21800),
            .in3(N__23390),
            .lcout(n16497),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12241_3_lut_LC_10_6_6.C_ON=1'b0;
    defparam i12241_3_lut_LC_10_6_6.SEQ_MODE=4'b0000;
    defparam i12241_3_lut_LC_10_6_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12241_3_lut_LC_10_6_6 (
            .in0(N__21887),
            .in1(N__23588),
            .in2(_gnd_net_),
            .in3(N__38826),
            .lcout(),
            .ltout(n15451_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_13177_LC_10_6_7.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_13177_LC_10_6_7.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_13177_LC_10_6_7.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_1__bdd_4_lut_13177_LC_10_6_7 (
            .in0(N__21791),
            .in1(N__33131),
            .in2(N__21785),
            .in3(N__33489),
            .lcout(n16380),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_11__i1_LC_10_7_0.C_ON=1'b0;
    defparam comm_buf_11__i1_LC_10_7_0.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i1_LC_10_7_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_buf_11__i1_LC_10_7_0 (
            .in0(N__50258),
            .in1(N__21776),
            .in2(_gnd_net_),
            .in3(N__44159),
            .lcout(comm_buf_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_11__i2_LC_10_7_1.C_ON=1'b0;
    defparam comm_buf_11__i2_LC_10_7_1.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i2_LC_10_7_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_11__i2_LC_10_7_1 (
            .in0(N__40118),
            .in1(N__21764),
            .in2(_gnd_net_),
            .in3(N__50264),
            .lcout(comm_buf_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_11__i3_LC_10_7_2.C_ON=1'b0;
    defparam comm_buf_11__i3_LC_10_7_2.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i3_LC_10_7_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_11__i3_LC_10_7_2 (
            .in0(N__50259),
            .in1(N__44887),
            .in2(_gnd_net_),
            .in3(N__22043),
            .lcout(comm_buf_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_11__i4_LC_10_7_3.C_ON=1'b0;
    defparam comm_buf_11__i4_LC_10_7_3.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i4_LC_10_7_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_11__i4_LC_10_7_3 (
            .in0(N__39928),
            .in1(N__22010),
            .in2(_gnd_net_),
            .in3(N__50265),
            .lcout(comm_buf_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_11__i5_LC_10_7_4.C_ON=1'b0;
    defparam comm_buf_11__i5_LC_10_7_4.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i5_LC_10_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_11__i5_LC_10_7_4 (
            .in0(N__50260),
            .in1(N__39804),
            .in2(_gnd_net_),
            .in3(N__21995),
            .lcout(comm_buf_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_11__i6_LC_10_7_5.C_ON=1'b0;
    defparam comm_buf_11__i6_LC_10_7_5.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i6_LC_10_7_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_11__i6_LC_10_7_5 (
            .in0(N__21974),
            .in1(N__50263),
            .in2(_gnd_net_),
            .in3(N__40706),
            .lcout(comm_buf_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_11__i7_LC_10_7_6.C_ON=1'b0;
    defparam comm_buf_11__i7_LC_10_7_6.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i7_LC_10_7_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_11__i7_LC_10_7_6 (
            .in0(N__50261),
            .in1(N__39394),
            .in2(_gnd_net_),
            .in3(N__21959),
            .lcout(comm_buf_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_11__i0_LC_10_7_7.C_ON=1'b0;
    defparam comm_buf_11__i0_LC_10_7_7.SEQ_MODE=4'b1000;
    defparam comm_buf_11__i0_LC_10_7_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_11__i0_LC_10_7_7 (
            .in0(N__21932),
            .in1(N__50262),
            .in2(_gnd_net_),
            .in3(N__39188),
            .lcout(comm_buf_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51120),
            .ce(N__23837),
            .sr(N__23822));
    defparam comm_buf_7__i7_LC_10_8_0.C_ON=1'b0;
    defparam comm_buf_7__i7_LC_10_8_0.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i7_LC_10_8_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_7__i7_LC_10_8_0 (
            .in0(N__49892),
            .in1(N__39395),
            .in2(_gnd_net_),
            .in3(N__21908),
            .lcout(comm_buf_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam comm_buf_7__i0_LC_10_8_1.C_ON=1'b0;
    defparam comm_buf_7__i0_LC_10_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i0_LC_10_8_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_7__i0_LC_10_8_1 (
            .in0(N__21878),
            .in1(N__49893),
            .in2(_gnd_net_),
            .in3(N__39205),
            .lcout(comm_buf_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam comm_buf_7__i6_LC_10_8_2.C_ON=1'b0;
    defparam comm_buf_7__i6_LC_10_8_2.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i6_LC_10_8_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_7__i6_LC_10_8_2 (
            .in0(N__49891),
            .in1(N__40730),
            .in2(_gnd_net_),
            .in3(N__21848),
            .lcout(comm_buf_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam comm_buf_7__i5_LC_10_8_3.C_ON=1'b0;
    defparam comm_buf_7__i5_LC_10_8_3.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i5_LC_10_8_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_buf_7__i5_LC_10_8_3 (
            .in0(N__49898),
            .in1(N__22217),
            .in2(_gnd_net_),
            .in3(N__39803),
            .lcout(comm_buf_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam comm_buf_7__i4_LC_10_8_4.C_ON=1'b0;
    defparam comm_buf_7__i4_LC_10_8_4.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i4_LC_10_8_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_7__i4_LC_10_8_4 (
            .in0(N__49890),
            .in1(N__39915),
            .in2(_gnd_net_),
            .in3(N__22190),
            .lcout(comm_buf_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam comm_buf_7__i3_LC_10_8_5.C_ON=1'b0;
    defparam comm_buf_7__i3_LC_10_8_5.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i3_LC_10_8_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_buf_7__i3_LC_10_8_5 (
            .in0(N__49897),
            .in1(N__22169),
            .in2(_gnd_net_),
            .in3(N__44886),
            .lcout(comm_buf_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam comm_buf_7__i2_LC_10_8_6.C_ON=1'b0;
    defparam comm_buf_7__i2_LC_10_8_6.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i2_LC_10_8_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_7__i2_LC_10_8_6 (
            .in0(N__49889),
            .in1(N__40120),
            .in2(_gnd_net_),
            .in3(N__22142),
            .lcout(comm_buf_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam comm_buf_7__i1_LC_10_8_7.C_ON=1'b0;
    defparam comm_buf_7__i1_LC_10_8_7.SEQ_MODE=4'b1000;
    defparam comm_buf_7__i1_LC_10_8_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_7__i1_LC_10_8_7 (
            .in0(N__44157),
            .in1(N__22112),
            .in2(_gnd_net_),
            .in3(N__49894),
            .lcout(comm_buf_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51128),
            .ce(N__23855),
            .sr(N__23846));
    defparam i12193_3_lut_LC_10_9_0.C_ON=1'b0;
    defparam i12193_3_lut_LC_10_9_0.SEQ_MODE=4'b0000;
    defparam i12193_3_lut_LC_10_9_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12193_3_lut_LC_10_9_0 (
            .in0(N__38836),
            .in1(N__22076),
            .in2(_gnd_net_),
            .in3(N__22061),
            .lcout(),
            .ltout(n15403_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16476_bdd_4_lut_LC_10_9_1.C_ON=1'b0;
    defparam n16476_bdd_4_lut_LC_10_9_1.SEQ_MODE=4'b0000;
    defparam n16476_bdd_4_lut_LC_10_9_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 n16476_bdd_4_lut_LC_10_9_1 (
            .in0(N__29339),
            .in1(N__22244),
            .in2(N__22049),
            .in3(N__33484),
            .lcout(),
            .ltout(n16479_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i4_LC_10_9_2.C_ON=1'b0;
    defparam comm_tx_buf_i4_LC_10_9_2.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i4_LC_10_9_2.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_tx_buf_i4_LC_10_9_2 (
            .in0(N__33485),
            .in1(N__22283),
            .in2(N__22046),
            .in3(N__33321),
            .lcout(comm_tx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51141),
            .ce(N__43109),
            .sr(N__22385));
    defparam i12190_3_lut_LC_10_9_3.C_ON=1'b0;
    defparam i12190_3_lut_LC_10_9_3.SEQ_MODE=4'b0000;
    defparam i12190_3_lut_LC_10_9_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12190_3_lut_LC_10_9_3 (
            .in0(N__22307),
            .in1(N__23510),
            .in2(_gnd_net_),
            .in3(N__38833),
            .lcout(n15400),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13244_LC_10_9_4.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13244_LC_10_9_4.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13244_LC_10_9_4.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_index_0__bdd_4_lut_13244_LC_10_9_4 (
            .in0(N__38835),
            .in1(N__22301),
            .in2(N__23960),
            .in3(N__33177),
            .lcout(),
            .ltout(n16452_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16452_bdd_4_lut_LC_10_9_5.C_ON=1'b0;
    defparam n16452_bdd_4_lut_LC_10_9_5.SEQ_MODE=4'b0000;
    defparam n16452_bdd_4_lut_LC_10_9_5.LUT_INIT=16'b1111000011001010;
    LogicCell40 n16452_bdd_4_lut_LC_10_9_5 (
            .in0(N__23318),
            .in1(N__22292),
            .in2(N__22286),
            .in3(N__33179),
            .lcout(n16455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12189_3_lut_LC_10_9_6.C_ON=1'b0;
    defparam i12189_3_lut_LC_10_9_6.SEQ_MODE=4'b0000;
    defparam i12189_3_lut_LC_10_9_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12189_3_lut_LC_10_9_6 (
            .in0(N__38834),
            .in1(N__22277),
            .in2(_gnd_net_),
            .in3(N__22262),
            .lcout(),
            .ltout(n15399_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_LC_10_9_7.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_LC_10_9_7.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_LC_10_9_7.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_index_1__bdd_4_lut_LC_10_9_7 (
            .in0(N__22253),
            .in1(N__33483),
            .in2(N__22247),
            .in3(N__33178),
            .lcout(n16476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12674_2_lut_LC_10_10_0.C_ON=1'b0;
    defparam i12674_2_lut_LC_10_10_0.SEQ_MODE=4'b0000;
    defparam i12674_2_lut_LC_10_10_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 i12674_2_lut_LC_10_10_0 (
            .in0(_gnd_net_),
            .in1(N__48039),
            .in2(_gnd_net_),
            .in3(N__34037),
            .lcout(),
            .ltout(n15633_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_13269_LC_10_10_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_13269_LC_10_10_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_13269_LC_10_10_1.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_13269_LC_10_10_1 (
            .in0(N__22424),
            .in1(N__45309),
            .in2(N__22238),
            .in3(N__47272),
            .lcout(),
            .ltout(n16458_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16458_bdd_4_lut_LC_10_10_2.C_ON=1'b0;
    defparam n16458_bdd_4_lut_LC_10_10_2.SEQ_MODE=4'b0000;
    defparam n16458_bdd_4_lut_LC_10_10_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16458_bdd_4_lut_LC_10_10_2 (
            .in0(N__47273),
            .in1(N__29198),
            .in2(N__22235),
            .in3(N__28013),
            .lcout(),
            .ltout(n16461_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_117_LC_10_10_3.C_ON=1'b0;
    defparam i1_4_lut_adj_117_LC_10_10_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_117_LC_10_10_3.LUT_INIT=16'b0100010011110100;
    LogicCell40 i1_4_lut_adj_117_LC_10_10_3 (
            .in0(N__39568),
            .in1(N__24038),
            .in2(N__22232),
            .in3(N__45654),
            .lcout(),
            .ltout(n76_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_118_LC_10_10_4.C_ON=1'b0;
    defparam i1_4_lut_adj_118_LC_10_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_118_LC_10_10_4.LUT_INIT=16'b1111100010001000;
    LogicCell40 i1_4_lut_adj_118_LC_10_10_4 (
            .in0(N__36960),
            .in1(N__22541),
            .in2(N__22430),
            .in3(N__40253),
            .lcout(),
            .ltout(n4_adj_1195_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i4_LC_10_10_5.C_ON=1'b0;
    defparam comm_buf_0__i4_LC_10_10_5.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i4_LC_10_10_5.LUT_INIT=16'b1100110011111010;
    LogicCell40 comm_buf_0__i4_LC_10_10_5 (
            .in0(N__36887),
            .in1(N__39922),
            .in2(N__22427),
            .in3(N__50291),
            .lcout(comm_buf_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51151),
            .ce(N__25266),
            .sr(N__24192));
    defparam i12816_2_lut_LC_10_10_6.C_ON=1'b0;
    defparam i12816_2_lut_LC_10_10_6.SEQ_MODE=4'b0000;
    defparam i12816_2_lut_LC_10_10_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12816_2_lut_LC_10_10_6 (
            .in0(_gnd_net_),
            .in1(N__48038),
            .in2(_gnd_net_),
            .in3(N__30062),
            .lcout(n15632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i2_LC_10_11_0.C_ON=1'b0;
    defparam comm_buf_0__i2_LC_10_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i2_LC_10_11_0.LUT_INIT=16'b1100111111001010;
    LogicCell40 comm_buf_0__i2_LC_10_11_0 (
            .in0(N__22418),
            .in1(N__40053),
            .in2(N__50324),
            .in3(N__22400),
            .lcout(comm_buf_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51164),
            .ce(N__25268),
            .sr(N__24186));
    defparam i127_4_lut_adj_96_LC_10_11_2.C_ON=1'b0;
    defparam i127_4_lut_adj_96_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam i127_4_lut_adj_96_LC_10_11_2.LUT_INIT=16'b1010000011001100;
    LogicCell40 i127_4_lut_adj_96_LC_10_11_2 (
            .in0(N__47254),
            .in1(N__27887),
            .in2(N__36734),
            .in3(N__45647),
            .lcout(n130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12699_2_lut_LC_10_11_3.C_ON=1'b0;
    defparam i12699_2_lut_LC_10_11_3.SEQ_MODE=4'b0000;
    defparam i12699_2_lut_LC_10_11_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12699_2_lut_LC_10_11_3 (
            .in0(_gnd_net_),
            .in1(N__34373),
            .in2(_gnd_net_),
            .in3(N__32108),
            .lcout(n15589),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i131_3_lut_LC_10_11_5.C_ON=1'b0;
    defparam i131_3_lut_LC_10_11_5.SEQ_MODE=4'b0000;
    defparam i131_3_lut_LC_10_11_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 i131_3_lut_LC_10_11_5 (
            .in0(N__26458),
            .in1(N__34819),
            .in2(_gnd_net_),
            .in3(N__47255),
            .lcout(),
            .ltout(n87_adj_1165_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i124_4_lut_LC_10_11_6.C_ON=1'b0;
    defparam i124_4_lut_LC_10_11_6.SEQ_MODE=4'b0000;
    defparam i124_4_lut_LC_10_11_6.LUT_INIT=16'b1111000010001000;
    LogicCell40 i124_4_lut_LC_10_11_6 (
            .in0(N__47256),
            .in1(N__26257),
            .in2(N__22412),
            .in3(N__45648),
            .lcout(),
            .ltout(n69_adj_1161_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_97_LC_10_11_7.C_ON=1'b0;
    defparam i1_4_lut_adj_97_LC_10_11_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_97_LC_10_11_7.LUT_INIT=16'b1100110001000000;
    LogicCell40 i1_4_lut_adj_97_LC_10_11_7 (
            .in0(N__39542),
            .in1(N__40241),
            .in2(N__22409),
            .in3(N__22406),
            .lcout(n8050),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_116_LC_10_12_1.C_ON=1'b0;
    defparam i1_4_lut_adj_116_LC_10_12_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_116_LC_10_12_1.LUT_INIT=16'b1111111100000001;
    LogicCell40 i1_4_lut_adj_116_LC_10_12_1 (
            .in0(N__45661),
            .in1(N__39569),
            .in2(N__47315),
            .in3(N__40886),
            .lcout(n8089),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12691_2_lut_LC_10_12_2.C_ON=1'b0;
    defparam i12691_2_lut_LC_10_12_2.SEQ_MODE=4'b0000;
    defparam i12691_2_lut_LC_10_12_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12691_2_lut_LC_10_12_2 (
            .in0(_gnd_net_),
            .in1(N__43532),
            .in2(_gnd_net_),
            .in3(N__32118),
            .lcout(n15587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i127_4_lut_adj_107_LC_10_12_5.C_ON=1'b0;
    defparam i127_4_lut_adj_107_LC_10_12_5.SEQ_MODE=4'b0000;
    defparam i127_4_lut_adj_107_LC_10_12_5.LUT_INIT=16'b1101100001010000;
    LogicCell40 i127_4_lut_adj_107_LC_10_12_5 (
            .in0(N__45662),
            .in1(N__40565),
            .in2(N__22532),
            .in3(N__47274),
            .lcout(),
            .ltout(n130_adj_1156_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_110_LC_10_12_6.C_ON=1'b0;
    defparam i1_4_lut_adj_110_LC_10_12_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_110_LC_10_12_6.LUT_INIT=16'b1100010011000000;
    LogicCell40 i1_4_lut_adj_110_LC_10_12_6 (
            .in0(N__39570),
            .in1(N__40211),
            .in2(N__22520),
            .in3(N__24113),
            .lcout(),
            .ltout(n8051_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i3_LC_10_12_7.C_ON=1'b0;
    defparam comm_buf_0__i3_LC_10_12_7.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i3_LC_10_12_7.LUT_INIT=16'b1010101011111100;
    LogicCell40 comm_buf_0__i3_LC_10_12_7 (
            .in0(N__44917),
            .in1(N__22517),
            .in2(N__22511),
            .in3(N__50343),
            .lcout(comm_buf_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51182),
            .ce(N__25270),
            .sr(N__24193));
    defparam \ADC_VAC4.ADC_DATA_i11_LC_10_13_1 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i11_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i11_LC_10_13_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i11_LC_10_13_1  (
            .in0(N__25897),
            .in1(N__26541),
            .in2(N__22508),
            .in3(N__27380),
            .lcout(buf_adcdata4_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51200),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i22_LC_10_13_2 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i22_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i22_LC_10_13_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i22_LC_10_13_2  (
            .in0(N__37461),
            .in1(N__52875),
            .in2(N__44602),
            .in3(N__26162),
            .lcout(cmd_rdadctmp_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51200),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i23_LC_10_13_3 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i23_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i23_LC_10_13_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i23_LC_10_13_3  (
            .in0(N__26163),
            .in1(N__37462),
            .in2(N__22710),
            .in3(N__52877),
            .lcout(cmd_rdadctmp_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51200),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i0_LC_10_13_4 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i0_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i0_LC_10_13_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i0_LC_10_13_4  (
            .in0(N__53123),
            .in1(N__22444),
            .in2(N__22478),
            .in3(N__52876),
            .lcout(buf_adcdata1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51200),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i15_LC_10_13_5 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i15_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i15_LC_10_13_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i15_LC_10_13_5  (
            .in0(N__52874),
            .in1(N__53124),
            .in2(N__22711),
            .in3(N__22684),
            .lcout(buf_adcdata1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51200),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i21_LC_10_13_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i21_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i21_LC_10_13_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i21_LC_10_13_7  (
            .in0(N__26404),
            .in1(N__27379),
            .in2(N__22670),
            .in3(N__26850),
            .lcout(cmd_rdadctmp_21_adj_1128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51200),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i12926_4_lut_LC_10_14_0 .C_ON=1'b0;
    defparam \ADC_VAC2.i12926_4_lut_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i12926_4_lut_LC_10_14_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ADC_VAC2.i12926_4_lut_LC_10_14_0  (
            .in0(N__22639),
            .in1(N__22627),
            .in2(N__22616),
            .in3(N__22600),
            .lcout(\ADC_VAC2.n15596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i12127_4_lut_LC_10_14_1 .C_ON=1'b0;
    defparam \ADC_VAC3.i12127_4_lut_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i12127_4_lut_LC_10_14_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC3.i12127_4_lut_LC_10_14_1  (
            .in0(N__22819),
            .in1(N__22834),
            .in2(N__22868),
            .in3(N__22849),
            .lcout(),
            .ltout(\ADC_VAC3.n15334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i12149_4_lut_LC_10_14_2 .C_ON=1'b0;
    defparam \ADC_VAC3.i12149_4_lut_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i12149_4_lut_LC_10_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC3.i12149_4_lut_LC_10_14_2  (
            .in0(N__22789),
            .in1(N__22882),
            .in2(N__22583),
            .in3(N__22771),
            .lcout(),
            .ltout(\ADC_VAC3.n15358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i12787_4_lut_LC_10_14_3 .C_ON=1'b0;
    defparam \ADC_VAC3.i12787_4_lut_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i12787_4_lut_LC_10_14_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_VAC3.i12787_4_lut_LC_10_14_3  (
            .in0(N__23066),
            .in1(N__22804),
            .in2(N__22580),
            .in3(N__49007),
            .lcout(),
            .ltout(\ADC_VAC3.n15602_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.adc_state_i0_LC_10_14_4 .C_ON=1'b0;
    defparam \ADC_VAC3.adc_state_i0_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.adc_state_i0_LC_10_14_4 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \ADC_VAC3.adc_state_i0_LC_10_14_4  (
            .in0(N__22983),
            .in1(N__23067),
            .in2(N__22577),
            .in3(N__48943),
            .lcout(adc_state_0_adj_1080),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51217),
            .ce(N__22574),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i1_4_lut_adj_7_LC_10_14_6 .C_ON=1'b0;
    defparam \ADC_VAC3.i1_4_lut_adj_7_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i1_4_lut_adj_7_LC_10_14_6 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_VAC3.i1_4_lut_adj_7_LC_10_14_6  (
            .in0(N__22982),
            .in1(N__48942),
            .in2(N__23129),
            .in3(N__30654),
            .lcout(\ADC_VAC3.n15259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i30_4_lut_LC_10_14_7 .C_ON=1'b0;
    defparam \ADC_VAC3.i30_4_lut_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i30_4_lut_LC_10_14_7 .LUT_INIT=16'b1011000110000001;
    LogicCell40 \ADC_VAC3.i30_4_lut_LC_10_14_7  (
            .in0(N__30655),
            .in1(N__22981),
            .in2(N__23069),
            .in3(N__23128),
            .lcout(\ADC_VAC3.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.bit_cnt_i0_LC_10_15_0 .C_ON=1'b1;
    defparam \ADC_VAC3.bit_cnt_i0_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i0_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i0_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__22883),
            .in2(_gnd_net_),
            .in3(N__22871),
            .lcout(\ADC_VAC3.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\ADC_VAC3.n13995 ),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC3.bit_cnt_i1_LC_10_15_1 .C_ON=1'b1;
    defparam \ADC_VAC3.bit_cnt_i1_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i1_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i1_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__22867),
            .in2(_gnd_net_),
            .in3(N__22853),
            .lcout(\ADC_VAC3.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC3.n13995 ),
            .carryout(\ADC_VAC3.n13996 ),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC3.bit_cnt_i2_LC_10_15_2 .C_ON=1'b1;
    defparam \ADC_VAC3.bit_cnt_i2_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i2_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i2_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__22850),
            .in2(_gnd_net_),
            .in3(N__22838),
            .lcout(\ADC_VAC3.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC3.n13996 ),
            .carryout(\ADC_VAC3.n13997 ),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC3.bit_cnt_i3_LC_10_15_3 .C_ON=1'b1;
    defparam \ADC_VAC3.bit_cnt_i3_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i3_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i3_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__22835),
            .in2(_gnd_net_),
            .in3(N__22823),
            .lcout(\ADC_VAC3.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC3.n13997 ),
            .carryout(\ADC_VAC3.n13998 ),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC3.bit_cnt_i4_LC_10_15_4 .C_ON=1'b1;
    defparam \ADC_VAC3.bit_cnt_i4_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i4_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i4_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__22820),
            .in2(_gnd_net_),
            .in3(N__22808),
            .lcout(\ADC_VAC3.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC3.n13998 ),
            .carryout(\ADC_VAC3.n13999 ),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC3.bit_cnt_i5_LC_10_15_5 .C_ON=1'b1;
    defparam \ADC_VAC3.bit_cnt_i5_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i5_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i5_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__22805),
            .in2(_gnd_net_),
            .in3(N__22793),
            .lcout(\ADC_VAC3.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC3.n13999 ),
            .carryout(\ADC_VAC3.n14000 ),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC3.bit_cnt_i6_LC_10_15_6 .C_ON=1'b1;
    defparam \ADC_VAC3.bit_cnt_i6_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i6_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i6_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__22790),
            .in2(_gnd_net_),
            .in3(N__22778),
            .lcout(\ADC_VAC3.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC3.n14000 ),
            .carryout(\ADC_VAC3.n14001 ),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC3.bit_cnt_i7_LC_10_15_7 .C_ON=1'b0;
    defparam \ADC_VAC3.bit_cnt_i7_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.bit_cnt_i7_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC3.bit_cnt_i7_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__22772),
            .in2(_gnd_net_),
            .in3(N__22775),
            .lcout(\ADC_VAC3.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51234),
            .ce(N__22991),
            .sr(N__22913));
    defparam \ADC_VAC1.ADC_DATA_i23_LC_10_16_1 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i23_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i23_LC_10_16_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i23_LC_10_16_1  (
            .in0(N__53064),
            .in1(N__22729),
            .in2(N__22760),
            .in3(N__52844),
            .lcout(buf_adcdata1_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51250),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i1_4_lut_LC_10_16_2 .C_ON=1'b0;
    defparam \ADC_VAC3.i1_4_lut_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i1_4_lut_LC_10_16_2 .LUT_INIT=16'b0000000101000100;
    LogicCell40 \ADC_VAC3.i1_4_lut_LC_10_16_2  (
            .in0(N__49020),
            .in1(N__22984),
            .in2(N__23124),
            .in3(N__23068),
            .lcout(\ADC_VAC3.n9514 ),
            .ltout(\ADC_VAC3.n9514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.i7638_2_lut_LC_10_16_3 .C_ON=1'b0;
    defparam \ADC_VAC3.i7638_2_lut_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC3.i7638_2_lut_LC_10_16_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ADC_VAC3.i7638_2_lut_LC_10_16_3  (
            .in0(N__22985),
            .in1(_gnd_net_),
            .in2(N__22916),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC3.n10744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_67_LC_10_16_4.C_ON=1'b0;
    defparam i1_2_lut_adj_67_LC_10_16_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_67_LC_10_16_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_67_LC_10_16_4 (
            .in0(_gnd_net_),
            .in1(N__27105),
            .in2(_gnd_net_),
            .in3(N__27033),
            .lcout(n15144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.bit_cnt_i0_LC_10_17_0 .C_ON=1'b1;
    defparam \ADC_VAC4.bit_cnt_i0_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i0_LC_10_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i0_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__24413),
            .in2(_gnd_net_),
            .in3(N__22901),
            .lcout(\ADC_VAC4.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\ADC_VAC4.n14002 ),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.bit_cnt_i1_LC_10_17_1 .C_ON=1'b1;
    defparam \ADC_VAC4.bit_cnt_i1_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i1_LC_10_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i1_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__24454),
            .in2(_gnd_net_),
            .in3(N__22898),
            .lcout(\ADC_VAC4.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC4.n14002 ),
            .carryout(\ADC_VAC4.n14003 ),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.bit_cnt_i2_LC_10_17_2 .C_ON=1'b1;
    defparam \ADC_VAC4.bit_cnt_i2_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i2_LC_10_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i2_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__24440),
            .in2(_gnd_net_),
            .in3(N__22895),
            .lcout(\ADC_VAC4.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC4.n14003 ),
            .carryout(\ADC_VAC4.n14004 ),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.bit_cnt_i3_LC_10_17_3 .C_ON=1'b1;
    defparam \ADC_VAC4.bit_cnt_i3_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i3_LC_10_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i3_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__24467),
            .in2(_gnd_net_),
            .in3(N__22892),
            .lcout(\ADC_VAC4.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC4.n14004 ),
            .carryout(\ADC_VAC4.n14005 ),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.bit_cnt_i4_LC_10_17_4 .C_ON=1'b1;
    defparam \ADC_VAC4.bit_cnt_i4_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i4_LC_10_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i4_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__24479),
            .in2(_gnd_net_),
            .in3(N__22889),
            .lcout(\ADC_VAC4.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC4.n14005 ),
            .carryout(\ADC_VAC4.n14006 ),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.bit_cnt_i5_LC_10_17_5 .C_ON=1'b1;
    defparam \ADC_VAC4.bit_cnt_i5_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i5_LC_10_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i5_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__24691),
            .in2(_gnd_net_),
            .in3(N__22886),
            .lcout(\ADC_VAC4.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC4.n14006 ),
            .carryout(\ADC_VAC4.n14007 ),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.bit_cnt_i6_LC_10_17_6 .C_ON=1'b1;
    defparam \ADC_VAC4.bit_cnt_i6_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i6_LC_10_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i6_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__24427),
            .in2(_gnd_net_),
            .in3(N__23246),
            .lcout(\ADC_VAC4.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC4.n14007 ),
            .carryout(\ADC_VAC4.n14008 ),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.bit_cnt_i7_LC_10_17_7 .C_ON=1'b0;
    defparam \ADC_VAC4.bit_cnt_i7_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.bit_cnt_i7_LC_10_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC4.bit_cnt_i7_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__24398),
            .in2(_gnd_net_),
            .in3(N__23243),
            .lcout(\ADC_VAC4.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51267),
            .ce(N__24668),
            .sr(N__24659));
    defparam \ADC_VAC4.ADC_DATA_i22_LC_11_3_2 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i22_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i22_LC_11_3_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i22_LC_11_3_2  (
            .in0(N__25961),
            .in1(N__29061),
            .in2(N__23438),
            .in3(N__27352),
            .lcout(buf_adcdata4_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51107),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i2_7352_7353_reset_LC_11_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_7352_7353_reset_LC_11_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i2_7352_7353_reset_LC_11_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_7352_7353_reset_LC_11_4_0  (
            .in0(N__23240),
            .in1(N__23219),
            .in2(_gnd_net_),
            .in3(N__23204),
            .lcout(\comm_spi.n10464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42455),
            .ce(),
            .sr(N__23186));
    defparam \ADC_VAC4.ADC_DATA_i19_LC_11_5_0 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i19_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i19_LC_11_5_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i19_LC_11_5_0  (
            .in0(N__25942),
            .in1(N__43017),
            .in2(N__25655),
            .in3(N__27524),
            .lcout(buf_adcdata4_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51109),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_11_5_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_11_5_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.RESET_I_0_105_2_lut_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__46604),
            .in2(_gnd_net_),
            .in3(N__24928),
            .lcout(\comm_spi.data_tx_7__N_828 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i21_LC_11_5_2 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i21_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i21_LC_11_5_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i21_LC_11_5_2  (
            .in0(N__25943),
            .in1(N__23166),
            .in2(N__23144),
            .in3(N__27525),
            .lcout(buf_adcdata4_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51109),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i29_LC_11_5_3 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i29_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i29_LC_11_5_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i29_LC_11_5_3  (
            .in0(N__26851),
            .in1(N__23139),
            .in2(N__27529),
            .in3(N__25624),
            .lcout(cmd_rdadctmp_29_adj_1120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51109),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i30_LC_11_5_4 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i30_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i30_LC_11_5_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i30_LC_11_5_4  (
            .in0(N__23140),
            .in1(N__27517),
            .in2(N__23434),
            .in3(N__26853),
            .lcout(cmd_rdadctmp_30_adj_1119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51109),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i31_LC_11_5_5 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i31_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i31_LC_11_5_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i31_LC_11_5_5  (
            .in0(N__26852),
            .in1(N__23413),
            .in2(N__27530),
            .in3(N__23430),
            .lcout(cmd_rdadctmp_31_adj_1118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51109),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i23_LC_11_5_7 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i23_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i23_LC_11_5_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i23_LC_11_5_7  (
            .in0(N__27516),
            .in1(N__25944),
            .in2(N__45867),
            .in3(N__23414),
            .lcout(buf_adcdata4_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51109),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_8__i7_LC_11_6_0.C_ON=1'b0;
    defparam comm_buf_8__i7_LC_11_6_0.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i7_LC_11_6_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_8__i7_LC_11_6_0 (
            .in0(N__50316),
            .in1(N__39334),
            .in2(_gnd_net_),
            .in3(N__23405),
            .lcout(comm_buf_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_8__i6_LC_11_6_1.C_ON=1'b0;
    defparam comm_buf_8__i6_LC_11_6_1.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i6_LC_11_6_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_8__i6_LC_11_6_1 (
            .in0(N__23381),
            .in1(N__40691),
            .in2(_gnd_net_),
            .in3(N__50320),
            .lcout(comm_buf_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_8__i5_LC_11_6_2.C_ON=1'b0;
    defparam comm_buf_8__i5_LC_11_6_2.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i5_LC_11_6_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_8__i5_LC_11_6_2 (
            .in0(N__50315),
            .in1(_gnd_net_),
            .in2(N__39795),
            .in3(N__23357),
            .lcout(comm_buf_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_8__i4_LC_11_6_3.C_ON=1'b0;
    defparam comm_buf_8__i4_LC_11_6_3.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i4_LC_11_6_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_8__i4_LC_11_6_3 (
            .in0(N__39859),
            .in1(N__23333),
            .in2(_gnd_net_),
            .in3(N__50319),
            .lcout(comm_buf_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_8__i3_LC_11_6_4.C_ON=1'b0;
    defparam comm_buf_8__i3_LC_11_6_4.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i3_LC_11_6_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_8__i3_LC_11_6_4 (
            .in0(N__50314),
            .in1(N__44856),
            .in2(_gnd_net_),
            .in3(N__23306),
            .lcout(comm_buf_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_8__i2_LC_11_6_5.C_ON=1'b0;
    defparam comm_buf_8__i2_LC_11_6_5.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i2_LC_11_6_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_8__i2_LC_11_6_5 (
            .in0(N__23273),
            .in1(N__40076),
            .in2(_gnd_net_),
            .in3(N__50318),
            .lcout(comm_buf_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_8__i1_LC_11_6_6.C_ON=1'b0;
    defparam comm_buf_8__i1_LC_11_6_6.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i1_LC_11_6_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_8__i1_LC_11_6_6 (
            .in0(N__50313),
            .in1(N__44099),
            .in2(_gnd_net_),
            .in3(N__23660),
            .lcout(comm_buf_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_8__i0_LC_11_6_7.C_ON=1'b0;
    defparam comm_buf_8__i0_LC_11_6_7.SEQ_MODE=4'b1000;
    defparam comm_buf_8__i0_LC_11_6_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_8__i0_LC_11_6_7 (
            .in0(N__23633),
            .in1(N__50317),
            .in2(_gnd_net_),
            .in3(N__39177),
            .lcout(comm_buf_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51112),
            .ce(N__25082),
            .sr(N__25067));
    defparam comm_buf_6__i7_LC_11_7_0.C_ON=1'b0;
    defparam comm_buf_6__i7_LC_11_7_0.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i7_LC_11_7_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_6__i7_LC_11_7_0 (
            .in0(N__39390),
            .in1(N__23603),
            .in2(_gnd_net_),
            .in3(N__50257),
            .lcout(comm_buf_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51115),
            .ce(N__23762),
            .sr(N__23743));
    defparam comm_buf_6__i6_LC_11_7_1.C_ON=1'b0;
    defparam comm_buf_6__i6_LC_11_7_1.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i6_LC_11_7_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_6__i6_LC_11_7_1 (
            .in0(N__50254),
            .in1(_gnd_net_),
            .in2(N__40722),
            .in3(N__23582),
            .lcout(comm_buf_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51115),
            .ce(N__23762),
            .sr(N__23743));
    defparam comm_buf_6__i5_LC_11_7_2.C_ON=1'b0;
    defparam comm_buf_6__i5_LC_11_7_2.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i5_LC_11_7_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_6__i5_LC_11_7_2 (
            .in0(N__39785),
            .in1(N__23552),
            .in2(_gnd_net_),
            .in3(N__50256),
            .lcout(comm_buf_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51115),
            .ce(N__23762),
            .sr(N__23743));
    defparam comm_buf_6__i4_LC_11_7_3.C_ON=1'b0;
    defparam comm_buf_6__i4_LC_11_7_3.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i4_LC_11_7_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_6__i4_LC_11_7_3 (
            .in0(N__50253),
            .in1(N__39887),
            .in2(_gnd_net_),
            .in3(N__23525),
            .lcout(comm_buf_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51115),
            .ce(N__23762),
            .sr(N__23743));
    defparam comm_buf_6__i3_LC_11_7_4.C_ON=1'b0;
    defparam comm_buf_6__i3_LC_11_7_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i3_LC_11_7_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_6__i3_LC_11_7_4 (
            .in0(N__23501),
            .in1(N__44885),
            .in2(_gnd_net_),
            .in3(N__50255),
            .lcout(comm_buf_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51115),
            .ce(N__23762),
            .sr(N__23743));
    defparam comm_buf_6__i2_LC_11_7_5.C_ON=1'b0;
    defparam comm_buf_6__i2_LC_11_7_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i2_LC_11_7_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_6__i2_LC_11_7_5 (
            .in0(N__50252),
            .in1(N__40117),
            .in2(_gnd_net_),
            .in3(N__23474),
            .lcout(comm_buf_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51115),
            .ce(N__23762),
            .sr(N__23743));
    defparam i1_4_lut_adj_237_LC_11_8_0.C_ON=1'b0;
    defparam i1_4_lut_adj_237_LC_11_8_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_237_LC_11_8_0.LUT_INIT=16'b1100010011000000;
    LogicCell40 i1_4_lut_adj_237_LC_11_8_0 (
            .in0(N__38787),
            .in1(N__42798),
            .in2(N__38559),
            .in3(N__25399),
            .lcout(n8907),
            .ltout(n8907_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7512_2_lut_LC_11_8_1.C_ON=1'b0;
    defparam i7512_2_lut_LC_11_8_1.SEQ_MODE=4'b0000;
    defparam i7512_2_lut_LC_11_8_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 i7512_2_lut_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23858),
            .in3(N__52450),
            .lcout(n10618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_247_LC_11_8_2.C_ON=1'b0;
    defparam i1_4_lut_adj_247_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_247_LC_11_8_2.LUT_INIT=16'b1100100011000000;
    LogicCell40 i1_4_lut_adj_247_LC_11_8_2 (
            .in0(N__38788),
            .in1(N__42799),
            .in2(N__38560),
            .in3(N__25400),
            .lcout(n8943),
            .ltout(n8943_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7519_2_lut_LC_11_8_3.C_ON=1'b0;
    defparam i7519_2_lut_LC_11_8_3.SEQ_MODE=4'b0000;
    defparam i7519_2_lut_LC_11_8_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 i7519_2_lut_LC_11_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23849),
            .in3(N__52451),
            .lcout(n10625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_275_LC_11_8_4.C_ON=1'b0;
    defparam i1_4_lut_adj_275_LC_11_8_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_275_LC_11_8_4.LUT_INIT=16'b1100100011000000;
    LogicCell40 i1_4_lut_adj_275_LC_11_8_4 (
            .in0(N__38789),
            .in1(N__42800),
            .in2(N__38561),
            .in3(N__25154),
            .lcout(n9123),
            .ltout(n9123_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7547_2_lut_LC_11_8_5.C_ON=1'b0;
    defparam i7547_2_lut_LC_11_8_5.SEQ_MODE=4'b0000;
    defparam i7547_2_lut_LC_11_8_5.LUT_INIT=16'b1111000000000000;
    LogicCell40 i7547_2_lut_LC_11_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23825),
            .in3(N__52452),
            .lcout(n10653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i0_LC_11_8_6.C_ON=1'b0;
    defparam comm_buf_6__i0_LC_11_8_6.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i0_LC_11_8_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_6__i0_LC_11_8_6 (
            .in0(N__39179),
            .in1(N__23816),
            .in2(_gnd_net_),
            .in3(N__50312),
            .lcout(comm_buf_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51121),
            .ce(N__23761),
            .sr(N__23744));
    defparam comm_buf_6__i1_LC_11_8_7.C_ON=1'b0;
    defparam comm_buf_6__i1_LC_11_8_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i1_LC_11_8_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_6__i1_LC_11_8_7 (
            .in0(N__50311),
            .in1(N__44156),
            .in2(_gnd_net_),
            .in3(N__23789),
            .lcout(comm_buf_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51121),
            .ce(N__23761),
            .sr(N__23744));
    defparam comm_buf_10__i2_LC_11_9_0.C_ON=1'b0;
    defparam comm_buf_10__i2_LC_11_9_0.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i2_LC_11_9_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_10__i2_LC_11_9_0 (
            .in0(N__40119),
            .in1(N__23723),
            .in2(_gnd_net_),
            .in3(N__50303),
            .lcout(comm_buf_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51129),
            .ce(N__25356),
            .sr(N__25319));
    defparam comm_buf_10__i3_LC_11_9_1.C_ON=1'b0;
    defparam comm_buf_10__i3_LC_11_9_1.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i3_LC_11_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_10__i3_LC_11_9_1 (
            .in0(N__50300),
            .in1(N__44888),
            .in2(_gnd_net_),
            .in3(N__23693),
            .lcout(comm_buf_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51129),
            .ce(N__25356),
            .sr(N__25319));
    defparam comm_buf_10__i4_LC_11_9_2.C_ON=1'b0;
    defparam comm_buf_10__i4_LC_11_9_2.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i4_LC_11_9_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_10__i4_LC_11_9_2 (
            .in0(N__39914),
            .in1(N__23978),
            .in2(_gnd_net_),
            .in3(N__50304),
            .lcout(comm_buf_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51129),
            .ce(N__25356),
            .sr(N__25319));
    defparam comm_buf_10__i7_LC_11_9_3.C_ON=1'b0;
    defparam comm_buf_10__i7_LC_11_9_3.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i7_LC_11_9_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_10__i7_LC_11_9_3 (
            .in0(N__50301),
            .in1(_gnd_net_),
            .in2(N__39401),
            .in3(N__23951),
            .lcout(comm_buf_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51129),
            .ce(N__25356),
            .sr(N__25319));
    defparam comm_buf_10__i0_LC_11_9_4.C_ON=1'b0;
    defparam comm_buf_10__i0_LC_11_9_4.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i0_LC_11_9_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_10__i0_LC_11_9_4 (
            .in0(N__39180),
            .in1(N__23915),
            .in2(_gnd_net_),
            .in3(N__50302),
            .lcout(comm_buf_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51129),
            .ce(N__25356),
            .sr(N__25319));
    defparam comm_cmd_1__bdd_4_lut_13235_LC_11_10_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_13235_LC_11_10_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_13235_LC_11_10_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_13235_LC_11_10_0 (
            .in0(N__28052),
            .in1(N__45289),
            .in2(N__31307),
            .in3(N__47251),
            .lcout(),
            .ltout(n16434_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16434_bdd_4_lut_LC_11_10_1.C_ON=1'b0;
    defparam n16434_bdd_4_lut_LC_11_10_1.SEQ_MODE=4'b0000;
    defparam n16434_bdd_4_lut_LC_11_10_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16434_bdd_4_lut_LC_11_10_1 (
            .in0(N__47252),
            .in1(N__27980),
            .in2(N__23882),
            .in3(N__29168),
            .lcout(),
            .ltout(n16437_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i108_4_lut_adj_132_LC_11_10_2.C_ON=1'b0;
    defparam i108_4_lut_adj_132_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam i108_4_lut_adj_132_LC_11_10_2.LUT_INIT=16'b1011100000110000;
    LogicCell40 i108_4_lut_adj_132_LC_11_10_2 (
            .in0(N__30902),
            .in1(N__45538),
            .in2(N__23879),
            .in3(N__47253),
            .lcout(n109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_136_LC_11_10_5.C_ON=1'b0;
    defparam i1_4_lut_adj_136_LC_11_10_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_136_LC_11_10_5.LUT_INIT=16'b1010111000000000;
    LogicCell40 i1_4_lut_adj_136_LC_11_10_5 (
            .in0(N__23876),
            .in1(N__42968),
            .in2(N__39581),
            .in3(N__40240),
            .lcout(),
            .ltout(n8054_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i6_LC_11_10_6.C_ON=1'b0;
    defparam comm_buf_0__i6_LC_11_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i6_LC_11_10_6.LUT_INIT=16'b1010101011111100;
    LogicCell40 comm_buf_0__i6_LC_11_10_6 (
            .in0(N__40731),
            .in1(N__27758),
            .in2(N__23870),
            .in3(N__50305),
            .lcout(comm_buf_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51142),
            .ce(N__25265),
            .sr(N__24187));
    defparam i106_4_lut_LC_11_11_0.C_ON=1'b0;
    defparam i106_4_lut_LC_11_11_0.SEQ_MODE=4'b0000;
    defparam i106_4_lut_LC_11_11_0.LUT_INIT=16'b1110010010100000;
    LogicCell40 i106_4_lut_LC_11_11_0 (
            .in0(N__47921),
            .in1(N__25757),
            .in2(N__41633),
            .in3(N__45646),
            .lcout(n59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i16_LC_11_11_1 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i16_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i16_LC_11_11_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i16_LC_11_11_1  (
            .in0(N__44359),
            .in1(N__49110),
            .in2(N__28493),
            .in3(N__26355),
            .lcout(buf_adcdata3_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51152),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i17_LC_11_11_2 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i17_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i17_LC_11_11_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i17_LC_11_11_2  (
            .in0(N__49109),
            .in1(N__44360),
            .in2(N__24014),
            .in3(N__27954),
            .lcout(buf_adcdata3_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51152),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i25_LC_11_11_3 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i25_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i25_LC_11_11_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i25_LC_11_11_3  (
            .in0(N__28489),
            .in1(N__24009),
            .in2(N__48831),
            .in3(N__49111),
            .lcout(cmd_rdadctmp_25_adj_1087),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51152),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i26_LC_11_11_4 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i26_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i26_LC_11_11_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i26_LC_11_11_4  (
            .in0(N__24010),
            .in1(N__48805),
            .in2(N__49202),
            .in3(N__26481),
            .lcout(cmd_rdadctmp_26_adj_1086),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51152),
            .ce(),
            .sr(_gnd_net_));
    defparam i7470_2_lut_LC_11_11_5.C_ON=1'b0;
    defparam i7470_2_lut_LC_11_11_5.SEQ_MODE=4'b0000;
    defparam i7470_2_lut_LC_11_11_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i7470_2_lut_LC_11_11_5 (
            .in0(_gnd_net_),
            .in1(N__52453),
            .in2(_gnd_net_),
            .in3(N__25224),
            .lcout(n10576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i7_LC_11_11_6 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i7_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i7_LC_11_11_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i7_LC_11_11_6  (
            .in0(N__48824),
            .in1(N__24269),
            .in2(N__49203),
            .in3(N__23992),
            .lcout(cmd_rdadctmp_7_adj_1105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51152),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i27_LC_11_11_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i27_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i27_LC_11_11_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i27_LC_11_11_7  (
            .in0(N__26847),
            .in1(N__25741),
            .in2(N__25651),
            .in3(N__27466),
            .lcout(cmd_rdadctmp_27_adj_1122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51152),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_13289_LC_11_12_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_13289_LC_11_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_13289_LC_11_12_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_13289_LC_11_12_0 (
            .in0(N__26432),
            .in1(N__45308),
            .in2(N__31394),
            .in3(N__47247),
            .lcout(),
            .ltout(n16500_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16500_bdd_4_lut_LC_11_12_1.C_ON=1'b0;
    defparam n16500_bdd_4_lut_LC_11_12_1.SEQ_MODE=4'b0000;
    defparam n16500_bdd_4_lut_LC_11_12_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16500_bdd_4_lut_LC_11_12_1 (
            .in0(N__47248),
            .in1(N__27995),
            .in2(N__23981),
            .in3(N__27971),
            .lcout(),
            .ltout(n16503_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_293_LC_11_12_2.C_ON=1'b0;
    defparam i1_4_lut_adj_293_LC_11_12_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_293_LC_11_12_2.LUT_INIT=16'b1011101000110000;
    LogicCell40 i1_4_lut_adj_293_LC_11_12_2 (
            .in0(N__31349),
            .in1(N__45657),
            .in2(N__24221),
            .in3(N__47249),
            .lcout(n4_adj_1280),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_295_LC_11_12_5.C_ON=1'b0;
    defparam i1_4_lut_adj_295_LC_11_12_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_295_LC_11_12_5.LUT_INIT=16'b1000101010001000;
    LogicCell40 i1_4_lut_adj_295_LC_11_12_5 (
            .in0(N__40210),
            .in1(N__24218),
            .in2(N__39580),
            .in3(N__24386),
            .lcout(),
            .ltout(n8047_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i0_LC_11_12_6.C_ON=1'b0;
    defparam comm_buf_0__i0_LC_11_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i0_LC_11_12_6.LUT_INIT=16'b1010101011111100;
    LogicCell40 comm_buf_0__i0_LC_11_12_6 (
            .in0(N__39201),
            .in1(N__32069),
            .in2(N__24212),
            .in3(N__50342),
            .lcout(comm_buf_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51165),
            .ce(N__25267),
            .sr(N__24188));
    defparam \ADC_VAC1.cmd_rdadctmp_i10_LC_11_13_1 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i10_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i10_LC_11_13_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i10_LC_11_13_1  (
            .in0(N__24155),
            .in1(N__52813),
            .in2(N__44451),
            .in3(N__26182),
            .lcout(cmd_rdadctmp_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51183),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_3__358_LC_11_13_2.C_ON=1'b0;
    defparam buf_control_3__358_LC_11_13_2.SEQ_MODE=4'b1000;
    defparam buf_control_3__358_LC_11_13_2.LUT_INIT=16'b1111000011011000;
    LogicCell40 buf_control_3__358_LC_11_13_2 (
            .in0(N__39650),
            .in1(N__43533),
            .in2(N__24128),
            .in3(N__41169),
            .lcout(buf_control_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51183),
            .ce(),
            .sr(_gnd_net_));
    defparam i124_4_lut_adj_108_LC_11_13_4.C_ON=1'b0;
    defparam i124_4_lut_adj_108_LC_11_13_4.SEQ_MODE=4'b0000;
    defparam i124_4_lut_adj_108_LC_11_13_4.LUT_INIT=16'b1011100010001000;
    LogicCell40 i124_4_lut_adj_108_LC_11_13_4 (
            .in0(N__26192),
            .in1(N__45658),
            .in2(N__24127),
            .in3(N__47250),
            .lcout(n69_adj_1029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i14_LC_11_13_5 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i14_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i14_LC_11_13_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i14_LC_11_13_5  (
            .in0(N__25882),
            .in1(N__24096),
            .in2(N__27353),
            .in3(N__26392),
            .lcout(buf_adcdata4_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51183),
            .ce(),
            .sr(_gnd_net_));
    defparam i112_4_lut_LC_11_14_0.C_ON=1'b0;
    defparam i112_4_lut_LC_11_14_0.SEQ_MODE=4'b0000;
    defparam i112_4_lut_LC_11_14_0.LUT_INIT=16'b0011000010001000;
    LogicCell40 i112_4_lut_LC_11_14_0 (
            .in0(N__24074),
            .in1(N__45655),
            .in2(N__24026),
            .in3(N__47243),
            .lcout(n61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_4__357_LC_11_14_1.C_ON=1'b0;
    defparam buf_control_4__357_LC_11_14_1.SEQ_MODE=4'b1000;
    defparam buf_control_4__357_LC_11_14_1.LUT_INIT=16'b1111101101000000;
    LogicCell40 buf_control_4__357_LC_11_14_1 (
            .in0(N__41171),
            .in1(N__39655),
            .in2(N__36989),
            .in3(N__24025),
            .lcout(buf_control_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51201),
            .ce(),
            .sr(_gnd_net_));
    defparam i127_4_lut_adj_294_LC_11_14_2.C_ON=1'b0;
    defparam i127_4_lut_adj_294_LC_11_14_2.SEQ_MODE=4'b0000;
    defparam i127_4_lut_adj_294_LC_11_14_2.LUT_INIT=16'b1011100010001000;
    LogicCell40 i127_4_lut_adj_294_LC_11_14_2 (
            .in0(N__26333),
            .in1(N__45656),
            .in2(N__24376),
            .in3(N__47244),
            .lcout(n69),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_0__361_LC_11_14_4.C_ON=1'b0;
    defparam buf_control_0__361_LC_11_14_4.SEQ_MODE=4'b1000;
    defparam buf_control_0__361_LC_11_14_4.LUT_INIT=16'b1111000011011000;
    LogicCell40 buf_control_0__361_LC_11_14_4 (
            .in0(N__39654),
            .in1(N__34118),
            .in2(N__24377),
            .in3(N__41170),
            .lcout(buf_control_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51201),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i28_LC_11_14_5 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i28_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i28_LC_11_14_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i28_LC_11_14_5  (
            .in0(N__48978),
            .in1(N__24237),
            .in2(N__25708),
            .in3(N__48785),
            .lcout(cmd_rdadctmp_28_adj_1084),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51201),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i9_LC_11_14_6.C_ON=1'b0;
    defparam buf_dds_i9_LC_11_14_6.SEQ_MODE=4'b1000;
    defparam buf_dds_i9_LC_11_14_6.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i9_LC_11_14_6 (
            .in0(N__34590),
            .in1(N__29227),
            .in2(N__41527),
            .in3(N__41380),
            .lcout(buf_dds_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51201),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i27_LC_11_14_7 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i27_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i27_LC_11_14_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i27_LC_11_14_7  (
            .in0(N__48977),
            .in1(N__26488),
            .in2(N__25707),
            .in3(N__48784),
            .lcout(cmd_rdadctmp_27_adj_1085),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51201),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1457_i1_4_lut_LC_11_15_0.C_ON=1'b0;
    defparam mux_1457_i1_4_lut_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam mux_1457_i1_4_lut_LC_11_15_0.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1457_i1_4_lut_LC_11_15_0 (
            .in0(N__24362),
            .in1(N__48004),
            .in2(N__24346),
            .in3(N__47246),
            .lcout(n4064),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i6_LC_11_15_1 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i6_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i6_LC_11_15_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i6_LC_11_15_1  (
            .in0(N__48755),
            .in1(N__24262),
            .in2(N__24290),
            .in3(N__49011),
            .lcout(cmd_rdadctmp_6_adj_1106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51218),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i29_LC_11_15_2 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i29_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i29_LC_11_15_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i29_LC_11_15_2  (
            .in0(N__24244),
            .in1(N__36861),
            .in2(N__49119),
            .in3(N__48756),
            .lcout(cmd_rdadctmp_29_adj_1083),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51218),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i13_LC_11_15_4 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i13_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i13_LC_11_15_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i13_LC_11_15_4  (
            .in0(N__27288),
            .in1(N__25883),
            .in2(N__26420),
            .in3(N__28616),
            .lcout(buf_adcdata4_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51218),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i17_LC_11_15_6 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i17_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i17_LC_11_15_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i17_LC_11_15_6  (
            .in0(N__32173),
            .in1(N__52809),
            .in2(N__24575),
            .in3(N__26183),
            .lcout(cmd_rdadctmp_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51218),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i19_LC_11_15_7 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i19_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i19_LC_11_15_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i19_LC_11_15_7  (
            .in0(N__26184),
            .in1(N__24552),
            .in2(N__52878),
            .in3(N__52917),
            .lcout(cmd_rdadctmp_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51218),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i9_LC_11_16_0 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i9_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i9_LC_11_16_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i9_LC_11_16_0  (
            .in0(N__52795),
            .in1(N__53085),
            .in2(N__24595),
            .in3(N__24574),
            .lcout(buf_adcdata1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51235),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i18_LC_11_16_2 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i18_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i18_LC_11_16_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i18_LC_11_16_2  (
            .in0(N__52796),
            .in1(N__24573),
            .in2(N__52921),
            .in3(N__26185),
            .lcout(cmd_rdadctmp_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51235),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i20_LC_11_16_4 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i20_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i20_LC_11_16_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i20_LC_11_16_4  (
            .in0(N__52797),
            .in1(N__46272),
            .in2(N__24557),
            .in3(N__26186),
            .lcout(cmd_rdadctmp_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51235),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i11_LC_11_16_5 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i11_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i11_LC_11_16_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i11_LC_11_16_5  (
            .in0(N__53084),
            .in1(N__52798),
            .in2(N__24532),
            .in3(N__24556),
            .lcout(buf_adcdata1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51235),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i8_LC_11_16_6 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i8_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i8_LC_11_16_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i8_LC_11_16_6  (
            .in0(N__44302),
            .in1(N__49118),
            .in2(N__38207),
            .in3(N__24501),
            .lcout(buf_adcdata3_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51235),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i12123_4_lut_LC_11_17_0 .C_ON=1'b0;
    defparam \ADC_VAC4.i12123_4_lut_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i12123_4_lut_LC_11_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC4.i12123_4_lut_LC_11_17_0  (
            .in0(N__24478),
            .in1(N__24466),
            .in2(N__24455),
            .in3(N__24439),
            .lcout(),
            .ltout(\ADC_VAC4.n15330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i12146_4_lut_LC_11_17_1 .C_ON=1'b0;
    defparam \ADC_VAC4.i12146_4_lut_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i12146_4_lut_LC_11_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC4.i12146_4_lut_LC_11_17_1  (
            .in0(N__24428),
            .in1(N__24412),
            .in2(N__24401),
            .in3(N__24397),
            .lcout(\ADC_VAC4.n15354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i12804_4_lut_LC_11_17_4 .C_ON=1'b0;
    defparam \ADC_VAC4.i12804_4_lut_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i12804_4_lut_LC_11_17_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ADC_VAC4.i12804_4_lut_LC_11_17_4  (
            .in0(N__27250),
            .in1(N__27009),
            .in2(N__24692),
            .in3(N__24677),
            .lcout(),
            .ltout(\ADC_VAC4.n15619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.adc_state_i0_LC_11_17_5 .C_ON=1'b0;
    defparam \ADC_VAC4.adc_state_i0_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.adc_state_i0_LC_11_17_5 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \ADC_VAC4.adc_state_i0_LC_11_17_5  (
            .in0(N__27010),
            .in1(N__27251),
            .in2(N__24671),
            .in3(N__27110),
            .lcout(adc_state_0_adj_1117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51251),
            .ce(N__26681),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i30_4_lut_LC_11_17_6 .C_ON=1'b0;
    defparam \ADC_VAC4.i30_4_lut_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i30_4_lut_LC_11_17_6 .LUT_INIT=16'b1100100001010001;
    LogicCell40 \ADC_VAC4.i30_4_lut_LC_11_17_6  (
            .in0(N__27109),
            .in1(N__27008),
            .in2(N__26669),
            .in3(N__30647),
            .lcout(\ADC_VAC4.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i1_4_lut_LC_11_18_3 .C_ON=1'b0;
    defparam \ADC_VAC4.i1_4_lut_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i1_4_lut_LC_11_18_3 .LUT_INIT=16'b0000000101000100;
    LogicCell40 \ADC_VAC4.i1_4_lut_LC_11_18_3  (
            .in0(N__27238),
            .in1(N__27111),
            .in2(N__26665),
            .in3(N__27007),
            .lcout(\ADC_VAC4.n9631 ),
            .ltout(\ADC_VAC4.n9631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i7677_2_lut_LC_11_18_4 .C_ON=1'b0;
    defparam \ADC_VAC4.i7677_2_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i7677_2_lut_LC_11_18_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ADC_VAC4.i7677_2_lut_LC_11_18_4  (
            .in0(N__27112),
            .in1(_gnd_net_),
            .in2(N__24662),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC4.n10783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i20_LC_12_3_6 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i20_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i20_LC_12_3_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i20_LC_12_3_6  (
            .in0(N__25960),
            .in1(N__24639),
            .in2(N__25625),
            .in3(N__27489),
            .lcout(buf_adcdata4_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51106),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_4_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_12_4_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_96_2_lut_LC_12_4_0  (
            .in0(N__46601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30954),
            .lcout(\comm_spi.data_tx_7__N_809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13092_4_lut_3_lut_LC_12_4_1 .C_ON=1'b0;
    defparam \comm_spi.i13092_4_lut_3_lut_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13092_4_lut_3_lut_LC_12_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i13092_4_lut_3_lut_LC_12_4_1  (
            .in0(N__24935),
            .in1(N__24889),
            .in2(_gnd_net_),
            .in3(N__46603),
            .lcout(\comm_spi.n16905 ),
            .ltout(\comm_spi.n16905_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_7356_7357_set_LC_12_4_2 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_7356_7357_set_LC_12_4_2 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i3_7356_7357_set_LC_12_4_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.data_tx_i3_7356_7357_set_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(N__24871),
            .in2(N__24617),
            .in3(N__24853),
            .lcout(\comm_spi.n10467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42447),
            .ce(),
            .sr(N__24614));
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_12_4_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_12_4_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_97_2_lut_LC_12_4_5  (
            .in0(N__24934),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46602),
            .lcout(\comm_spi.data_tx_7__N_810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_12_4_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_12_4_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_103_2_lut_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(N__46640),
            .in2(_gnd_net_),
            .in3(N__46600),
            .lcout(\comm_spi.data_tx_7__N_822 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_7356_7357_reset_LC_12_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_7356_7357_reset_LC_12_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i3_7356_7357_reset_LC_12_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_7356_7357_reset_LC_12_5_0  (
            .in0(N__24890),
            .in1(N__24878),
            .in2(_gnd_net_),
            .in3(N__24854),
            .lcout(\comm_spi.n10468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42459),
            .ce(),
            .sr(N__30932));
    defparam comm_buf_9__i5_LC_12_6_0.C_ON=1'b0;
    defparam comm_buf_9__i5_LC_12_6_0.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i5_LC_12_6_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_9__i5_LC_12_6_0 (
            .in0(N__39766),
            .in1(N__24842),
            .in2(_gnd_net_),
            .in3(N__50309),
            .lcout(comm_buf_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51108),
            .ce(N__25031),
            .sr(N__25012));
    defparam comm_buf_9__i6_LC_12_6_1.C_ON=1'b0;
    defparam comm_buf_9__i6_LC_12_6_1.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i6_LC_12_6_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_9__i6_LC_12_6_1 (
            .in0(N__50307),
            .in1(N__40690),
            .in2(_gnd_net_),
            .in3(N__24812),
            .lcout(comm_buf_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51108),
            .ce(N__25031),
            .sr(N__25012));
    defparam comm_buf_9__i7_LC_12_6_2.C_ON=1'b0;
    defparam comm_buf_9__i7_LC_12_6_2.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i7_LC_12_6_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_9__i7_LC_12_6_2 (
            .in0(N__39333),
            .in1(N__24782),
            .in2(_gnd_net_),
            .in3(N__50310),
            .lcout(comm_buf_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51108),
            .ce(N__25031),
            .sr(N__25012));
    defparam comm_buf_9__i2_LC_12_6_3.C_ON=1'b0;
    defparam comm_buf_9__i2_LC_12_6_3.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i2_LC_12_6_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_9__i2_LC_12_6_3 (
            .in0(N__50306),
            .in1(N__40075),
            .in2(_gnd_net_),
            .in3(N__24755),
            .lcout(comm_buf_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51108),
            .ce(N__25031),
            .sr(N__25012));
    defparam comm_buf_9__i1_LC_12_6_4.C_ON=1'b0;
    defparam comm_buf_9__i1_LC_12_6_4.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i1_LC_12_6_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_9__i1_LC_12_6_4 (
            .in0(N__44098),
            .in1(N__24725),
            .in2(_gnd_net_),
            .in3(N__50308),
            .lcout(comm_buf_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51108),
            .ce(N__25031),
            .sr(N__25012));
    defparam i7533_2_lut_LC_12_7_0.C_ON=1'b0;
    defparam i7533_2_lut_LC_12_7_0.SEQ_MODE=4'b0000;
    defparam i7533_2_lut_LC_12_7_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 i7533_2_lut_LC_12_7_0 (
            .in0(_gnd_net_),
            .in1(N__52385),
            .in2(_gnd_net_),
            .in3(N__25029),
            .lcout(n10639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_231_LC_12_7_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_231_LC_12_7_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_231_LC_12_7_1.LUT_INIT=16'b0000010000000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_231_LC_12_7_1 (
            .in0(N__50601),
            .in1(N__33294),
            .in2(N__33488),
            .in3(N__27861),
            .lcout(n13470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_234_LC_12_7_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_234_LC_12_7_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_234_LC_12_7_2.LUT_INIT=16'b0000000000100000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_234_LC_12_7_2 (
            .in0(N__27862),
            .in1(N__25192),
            .in2(N__33328),
            .in3(N__33460),
            .lcout(),
            .ltout(n15161_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_268_LC_12_7_3.C_ON=1'b0;
    defparam i1_4_lut_adj_268_LC_12_7_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_268_LC_12_7_3.LUT_INIT=16'b1101110000000000;
    LogicCell40 i1_4_lut_adj_268_LC_12_7_3 (
            .in0(N__50602),
            .in1(N__38534),
            .in2(N__25085),
            .in3(N__42795),
            .lcout(n9027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_255_LC_12_7_4.C_ON=1'b0;
    defparam i1_4_lut_adj_255_LC_12_7_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_255_LC_12_7_4.LUT_INIT=16'b1010001010100000;
    LogicCell40 i1_4_lut_adj_255_LC_12_7_4 (
            .in0(N__42796),
            .in1(N__25421),
            .in2(N__38548),
            .in3(N__25166),
            .lcout(n8997),
            .ltout(n8997_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7526_2_lut_LC_12_7_5.C_ON=1'b0;
    defparam i7526_2_lut_LC_12_7_5.SEQ_MODE=4'b0000;
    defparam i7526_2_lut_LC_12_7_5.LUT_INIT=16'b1010000010100000;
    LogicCell40 i7526_2_lut_LC_12_7_5 (
            .in0(N__52386),
            .in1(_gnd_net_),
            .in2(N__25070),
            .in3(_gnd_net_),
            .lcout(n10632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_429_i6_2_lut_LC_12_7_6.C_ON=1'b0;
    defparam equal_429_i6_2_lut_LC_12_7_6.SEQ_MODE=4'b0000;
    defparam equal_429_i6_2_lut_LC_12_7_6.LUT_INIT=16'b1111111101010101;
    LogicCell40 equal_429_i6_2_lut_LC_12_7_6 (
            .in0(N__33295),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33459),
            .lcout(n6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_9__i0_LC_12_7_7.C_ON=1'b0;
    defparam comm_buf_9__i0_LC_12_7_7.SEQ_MODE=4'b1000;
    defparam comm_buf_9__i0_LC_12_7_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_9__i0_LC_12_7_7 (
            .in0(N__25061),
            .in1(N__50266),
            .in2(_gnd_net_),
            .in3(N__39178),
            .lcout(comm_buf_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51111),
            .ce(N__25030),
            .sr(N__25013));
    defparam comm_index_0__bdd_4_lut_13210_LC_12_8_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13210_LC_12_8_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13210_LC_12_8_0.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13210_LC_12_8_0 (
            .in0(N__33102),
            .in1(N__24941),
            .in2(N__24995),
            .in3(N__38785),
            .lcout(n16422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_10__i1_LC_12_8_1.C_ON=1'b0;
    defparam comm_buf_10__i1_LC_12_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i1_LC_12_8_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_10__i1_LC_12_8_1 (
            .in0(N__50215),
            .in1(N__44151),
            .in2(_gnd_net_),
            .in3(N__24965),
            .lcout(comm_buf_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51113),
            .ce(N__25357),
            .sr(N__25317));
    defparam i12638_2_lut_LC_12_8_2.C_ON=1'b0;
    defparam i12638_2_lut_LC_12_8_2.SEQ_MODE=4'b0000;
    defparam i12638_2_lut_LC_12_8_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12638_2_lut_LC_12_8_2 (
            .in0(N__33100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38784),
            .lcout(n15670),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_243_LC_12_8_4.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_243_LC_12_8_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_243_LC_12_8_4.LUT_INIT=16'b1110010010100000;
    LogicCell40 i1_4_lut_4_lut_adj_243_LC_12_8_4 (
            .in0(N__52449),
            .in1(N__31055),
            .in2(N__51928),
            .in3(N__31124),
            .lcout(n8763),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_273_LC_12_8_5.C_ON=1'b0;
    defparam i1_2_lut_adj_273_LC_12_8_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_273_LC_12_8_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_273_LC_12_8_5 (
            .in0(_gnd_net_),
            .in1(N__33101),
            .in2(_gnd_net_),
            .in3(N__25165),
            .lcout(n13497),
            .ltout(n13497_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_269_LC_12_8_6.C_ON=1'b0;
    defparam i1_4_lut_adj_269_LC_12_8_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_269_LC_12_8_6.LUT_INIT=16'b1011101000000000;
    LogicCell40 i1_4_lut_adj_269_LC_12_8_6 (
            .in0(N__38558),
            .in1(N__38786),
            .in2(N__25148),
            .in3(N__42797),
            .lcout(n9045),
            .ltout(n9045_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7540_2_lut_LC_12_8_7.C_ON=1'b0;
    defparam i7540_2_lut_LC_12_8_7.SEQ_MODE=4'b0000;
    defparam i7540_2_lut_LC_12_8_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i7540_2_lut_LC_12_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25145),
            .in3(N__52448),
            .lcout(n10646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_13264_LC_12_9_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_13264_LC_12_9_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_13264_LC_12_9_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_13264_LC_12_9_0 (
            .in0(N__25094),
            .in1(N__33097),
            .in2(N__25142),
            .in3(N__38781),
            .lcout(n16488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_10__i6_LC_12_9_1.C_ON=1'b0;
    defparam comm_buf_10__i6_LC_12_9_1.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i6_LC_12_9_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_10__i6_LC_12_9_1 (
            .in0(N__50201),
            .in1(_gnd_net_),
            .in2(N__25115),
            .in3(N__40723),
            .lcout(comm_buf_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51118),
            .ce(N__25355),
            .sr(N__25313));
    defparam i1_3_lut_4_lut_adj_260_LC_12_9_2.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_260_LC_12_9_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_260_LC_12_9_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 i1_3_lut_4_lut_adj_260_LC_12_9_2 (
            .in0(N__50597),
            .in1(N__33249),
            .in2(N__33449),
            .in3(N__27856),
            .lcout(n13457),
            .ltout(n13457_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12761_2_lut_LC_12_9_3.C_ON=1'b0;
    defparam i12761_2_lut_LC_12_9_3.SEQ_MODE=4'b0000;
    defparam i12761_2_lut_LC_12_9_3.LUT_INIT=16'b0000000011110000;
    LogicCell40 i12761_2_lut_LC_12_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25088),
            .in3(N__25417),
            .lcout(),
            .ltout(n15565_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20_4_lut_LC_12_9_4.C_ON=1'b0;
    defparam i20_4_lut_LC_12_9_4.SEQ_MODE=4'b0000;
    defparam i20_4_lut_LC_12_9_4.LUT_INIT=16'b1101000111000000;
    LogicCell40 i20_4_lut_LC_12_9_4 (
            .in0(N__50598),
            .in1(N__50200),
            .in2(N__25463),
            .in3(N__33626),
            .lcout(),
            .ltout(n13_adj_1257_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_219_LC_12_9_5.C_ON=1'b0;
    defparam i1_3_lut_adj_219_LC_12_9_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_219_LC_12_9_5.LUT_INIT=16'b1111110000000000;
    LogicCell40 i1_3_lut_adj_219_LC_12_9_5 (
            .in0(_gnd_net_),
            .in1(N__25581),
            .in2(N__25460),
            .in3(N__42856),
            .lcout(n8823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i61_2_lut_LC_12_9_6.C_ON=1'b0;
    defparam i61_2_lut_LC_12_9_6.SEQ_MODE=4'b0000;
    defparam i61_2_lut_LC_12_9_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i61_2_lut_LC_12_9_6 (
            .in0(_gnd_net_),
            .in1(N__33096),
            .in2(_gnd_net_),
            .in3(N__38780),
            .lcout(n41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_245_LC_12_9_7.C_ON=1'b0;
    defparam i1_2_lut_adj_245_LC_12_9_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_245_LC_12_9_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_adj_245_LC_12_9_7 (
            .in0(N__33098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25406),
            .lcout(n13458),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_10__i5_LC_12_10_1.C_ON=1'b0;
    defparam comm_buf_10__i5_LC_12_10_1.SEQ_MODE=4'b1000;
    defparam comm_buf_10__i5_LC_12_10_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_10__i5_LC_12_10_1 (
            .in0(N__50211),
            .in1(_gnd_net_),
            .in2(N__39802),
            .in3(N__25391),
            .lcout(comm_buf_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51125),
            .ce(N__25358),
            .sr(N__25318));
    defparam equal_436_i5_2_lut_LC_12_10_2.C_ON=1'b0;
    defparam equal_436_i5_2_lut_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam equal_436_i5_2_lut_LC_12_10_2.LUT_INIT=16'b1100110011111111;
    LogicCell40 equal_436_i5_2_lut_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(N__33099),
            .in2(_gnd_net_),
            .in3(N__38782),
            .lcout(n5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_256_LC_12_10_3.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_256_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_256_LC_12_10_3.LUT_INIT=16'b0001111100001111;
    LogicCell40 i1_3_lut_4_lut_adj_256_LC_12_10_3 (
            .in0(N__38783),
            .in1(N__33103),
            .in2(N__50322),
            .in3(N__31074),
            .lcout(),
            .ltout(n11_adj_1279_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_142_LC_12_10_4.C_ON=1'b0;
    defparam i1_4_lut_adj_142_LC_12_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_142_LC_12_10_4.LUT_INIT=16'b1000100010101000;
    LogicCell40 i1_4_lut_adj_142_LC_12_10_4 (
            .in0(N__42862),
            .in1(N__25582),
            .in2(N__25277),
            .in3(N__50599),
            .lcout(n8654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i36_4_lut_LC_12_10_5.C_ON=1'b0;
    defparam i36_4_lut_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam i36_4_lut_LC_12_10_5.LUT_INIT=16'b0100111001000100;
    LogicCell40 i36_4_lut_LC_12_10_5 (
            .in0(N__50210),
            .in1(N__37079),
            .in2(N__25196),
            .in3(N__31075),
            .lcout(),
            .ltout(n17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_179_LC_12_10_6.C_ON=1'b0;
    defparam i1_4_lut_adj_179_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_179_LC_12_10_6.LUT_INIT=16'b1000100010101000;
    LogicCell40 i1_4_lut_adj_179_LC_12_10_6 (
            .in0(N__42863),
            .in1(N__25583),
            .in2(N__25532),
            .in3(N__50600),
            .lcout(n8702),
            .ltout(n8702_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7477_2_lut_LC_12_10_7.C_ON=1'b0;
    defparam i7477_2_lut_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam i7477_2_lut_LC_12_10_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i7477_2_lut_LC_12_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25529),
            .in3(N__52376),
            .lcout(n10583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.i4_4_lut_LC_12_11_0 .C_ON=1'b0;
    defparam \CLOCK_DDS.i4_4_lut_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \CLOCK_DDS.i4_4_lut_LC_12_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CLOCK_DDS.i4_4_lut_LC_12_11_0  (
            .in0(N__25525),
            .in1(N__25515),
            .in2(N__25504),
            .in3(N__48381),
            .lcout(n10_adj_1172),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.bit_cnt_i3_LC_12_11_1 .C_ON=1'b0;
    defparam \CLOCK_DDS.bit_cnt_i3_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.bit_cnt_i3_LC_12_11_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \CLOCK_DDS.bit_cnt_i3_LC_12_11_1  (
            .in0(N__25517),
            .in1(N__25526),
            .in2(N__25505),
            .in3(N__31144),
            .lcout(bit_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51136),
            .ce(N__48548),
            .sr(N__31193));
    defparam \CLOCK_DDS.bit_cnt_i2_LC_12_11_2 .C_ON=1'b0;
    defparam \CLOCK_DDS.bit_cnt_i2_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.bit_cnt_i2_LC_12_11_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \CLOCK_DDS.bit_cnt_i2_LC_12_11_2  (
            .in0(N__31142),
            .in1(N__25500),
            .in2(_gnd_net_),
            .in3(N__25516),
            .lcout(bit_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51136),
            .ce(N__48548),
            .sr(N__31193));
    defparam \CLOCK_DDS.bit_cnt_i1_LC_12_11_3 .C_ON=1'b0;
    defparam \CLOCK_DDS.bit_cnt_i1_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.bit_cnt_i1_LC_12_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLOCK_DDS.bit_cnt_i1_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__25499),
            .in2(_gnd_net_),
            .in3(N__31143),
            .lcout(bit_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51136),
            .ce(N__48548),
            .sr(N__31193));
    defparam comm_cmd_1__bdd_4_lut_LC_12_11_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_LC_12_11_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_LC_12_11_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_LC_12_11_4 (
            .in0(N__31772),
            .in1(N__45218),
            .in2(N__28004),
            .in3(N__47140),
            .lcout(),
            .ltout(n16524_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16524_bdd_4_lut_LC_12_11_5.C_ON=1'b0;
    defparam n16524_bdd_4_lut_LC_12_11_5.SEQ_MODE=4'b0000;
    defparam n16524_bdd_4_lut_LC_12_11_5.LUT_INIT=16'b1111010010100100;
    LogicCell40 n16524_bdd_4_lut_LC_12_11_5 (
            .in0(N__47141),
            .in1(N__29183),
            .in2(N__25469),
            .in3(N__29405),
            .lcout(),
            .ltout(n16527_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_78_LC_12_11_6.C_ON=1'b0;
    defparam i1_4_lut_adj_78_LC_12_11_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_78_LC_12_11_6.LUT_INIT=16'b1011101000110000;
    LogicCell40 i1_4_lut_adj_78_LC_12_11_6 (
            .in0(N__33989),
            .in1(N__45645),
            .in2(N__25466),
            .in3(N__47142),
            .lcout(),
            .ltout(n4_adj_1264_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_82_LC_12_11_7.C_ON=1'b0;
    defparam i1_4_lut_adj_82_LC_12_11_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_82_LC_12_11_7.LUT_INIT=16'b1100010011000000;
    LogicCell40 i1_4_lut_adj_82_LC_12_11_7 (
            .in0(N__39541),
            .in1(N__40239),
            .in2(N__26015),
            .in3(N__27893),
            .lcout(n8055),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i15_LC_12_12_0 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i15_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i15_LC_12_12_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i15_LC_12_12_0  (
            .in0(N__25921),
            .in1(N__26326),
            .in2(N__25995),
            .in3(N__27398),
            .lcout(buf_adcdata4_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i16_LC_12_12_1 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i16_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i16_LC_12_12_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \ADC_VAC4.ADC_DATA_i16_LC_12_12_1  (
            .in0(N__27393),
            .in1(N__26309),
            .in2(N__47359),
            .in3(N__25923),
            .lcout(buf_adcdata4_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.ADC_DATA_i17_LC_12_12_2 .C_ON=1'b0;
    defparam \ADC_VAC4.ADC_DATA_i17_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.ADC_DATA_i17_LC_12_12_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC4.ADC_DATA_i17_LC_12_12_2  (
            .in0(N__25922),
            .in1(N__25779),
            .in2(N__26294),
            .in3(N__27399),
            .lcout(buf_adcdata4_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51147),
            .ce(),
            .sr(_gnd_net_));
    defparam i109_3_lut_LC_12_12_3.C_ON=1'b0;
    defparam i109_3_lut_LC_12_12_3.SEQ_MODE=4'b0000;
    defparam i109_3_lut_LC_12_12_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i109_3_lut_LC_12_12_3 (
            .in0(N__25668),
            .in1(N__28027),
            .in2(_gnd_net_),
            .in3(N__47238),
            .lcout(n71),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i26_LC_12_12_4 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i26_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i26_LC_12_12_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i26_LC_12_12_4  (
            .in0(N__26289),
            .in1(N__27394),
            .in2(N__25740),
            .in3(N__26849),
            .lcout(cmd_rdadctmp_26_adj_1123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i19_LC_12_12_5 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i19_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i19_LC_12_12_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i19_LC_12_12_5  (
            .in0(N__44367),
            .in1(N__49233),
            .in2(N__25715),
            .in3(N__26212),
            .lcout(buf_adcdata3_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i23_LC_12_12_6 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i23_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i23_LC_12_12_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i23_LC_12_12_6  (
            .in0(N__49232),
            .in1(N__44368),
            .in2(N__29396),
            .in3(N__25669),
            .lcout(buf_adcdata3_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i28_LC_12_12_7 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i28_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i28_LC_12_12_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i28_LC_12_12_7  (
            .in0(N__25647),
            .in1(N__25605),
            .in2(N__27465),
            .in3(N__26848),
            .lcout(cmd_rdadctmp_28_adj_1121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i24_LC_12_13_0 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i24_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i24_LC_12_13_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i24_LC_12_13_0  (
            .in0(N__26810),
            .in1(N__26325),
            .in2(N__27469),
            .in3(N__26307),
            .lcout(cmd_rdadctmp_24_adj_1125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51160),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i23_LC_12_13_1 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i23_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i23_LC_12_13_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i23_LC_12_13_1  (
            .in0(N__26393),
            .in1(N__27410),
            .in2(N__26327),
            .in3(N__26811),
            .lcout(cmd_rdadctmp_23_adj_1126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51160),
            .ce(),
            .sr(_gnd_net_));
    defparam i3181_3_lut_LC_12_13_2.C_ON=1'b0;
    defparam i3181_3_lut_LC_12_13_2.SEQ_MODE=4'b0000;
    defparam i3181_3_lut_LC_12_13_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 i3181_3_lut_LC_12_13_2 (
            .in0(N__31617),
            .in1(N__29904),
            .in2(_gnd_net_),
            .in3(N__40528),
            .lcout(n8_adj_1227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_279_LC_12_13_3.C_ON=1'b0;
    defparam i3_4_lut_adj_279_LC_12_13_3.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_279_LC_12_13_3.LUT_INIT=16'b0000001000000000;
    LogicCell40 i3_4_lut_adj_279_LC_12_13_3 (
            .in0(N__32812),
            .in1(N__28226),
            .in2(N__32912),
            .in3(N__28523),
            .lcout(n8_adj_1212),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i25_LC_12_13_5 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i25_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i25_LC_12_13_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i25_LC_12_13_5  (
            .in0(N__26308),
            .in1(N__27411),
            .in2(N__26293),
            .in3(N__26812),
            .lcout(cmd_rdadctmp_25_adj_1124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51160),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_2__359_LC_12_13_6.C_ON=1'b0;
    defparam buf_control_2__359_LC_12_13_6.SEQ_MODE=4'b1000;
    defparam buf_control_2__359_LC_12_13_6.LUT_INIT=16'b1111000011011000;
    LogicCell40 buf_control_2__359_LC_12_13_6 (
            .in0(N__39640),
            .in1(N__34408),
            .in2(N__26253),
            .in3(N__41167),
            .lcout(M_POW),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51160),
            .ce(),
            .sr(_gnd_net_));
    defparam i131_3_lut_adj_102_LC_12_13_7.C_ON=1'b0;
    defparam i131_3_lut_adj_102_LC_12_13_7.SEQ_MODE=4'b0000;
    defparam i131_3_lut_adj_102_LC_12_13_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 i131_3_lut_adj_102_LC_12_13_7 (
            .in0(N__26211),
            .in1(N__34787),
            .in2(_gnd_net_),
            .in3(N__47245),
            .lcout(n87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.cmd_rdadctmp_i21_LC_12_14_1 .C_ON=1'b0;
    defparam \ADC_VAC1.cmd_rdadctmp_i21_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.cmd_rdadctmp_i21_LC_12_14_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC1.cmd_rdadctmp_i21_LC_12_14_1  (
            .in0(N__44583),
            .in1(N__52793),
            .in2(N__46285),
            .in3(N__26181),
            .lcout(cmd_rdadctmp_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51177),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i6_LC_12_14_2.C_ON=1'b0;
    defparam buf_dds_i6_LC_12_14_2.SEQ_MODE=4'b1000;
    defparam buf_dds_i6_LC_12_14_2.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i6_LC_12_14_2 (
            .in0(N__33962),
            .in1(N__34617),
            .in2(N__41526),
            .in3(N__41373),
            .lcout(buf_dds_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51177),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_1__360_LC_12_14_3.C_ON=1'b0;
    defparam buf_control_1__360_LC_12_14_3.SEQ_MODE=4'b1000;
    defparam buf_control_1__360_LC_12_14_3.LUT_INIT=16'b1010101011001010;
    LogicCell40 buf_control_1__360_LC_12_14_3 (
            .in0(N__27915),
            .in1(N__34591),
            .in2(N__39663),
            .in3(N__41168),
            .lcout(M_DCSEL),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51177),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i18_LC_12_14_4 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i18_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i18_LC_12_14_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i18_LC_12_14_4  (
            .in0(N__44369),
            .in1(N__49189),
            .in2(N__26492),
            .in3(N__26451),
            .lcout(buf_adcdata3_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51177),
            .ce(),
            .sr(_gnd_net_));
    defparam i12630_2_lut_LC_12_14_6.C_ON=1'b0;
    defparam i12630_2_lut_LC_12_14_6.SEQ_MODE=4'b0000;
    defparam i12630_2_lut_LC_12_14_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12630_2_lut_LC_12_14_6 (
            .in0(N__32276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47917),
            .lcout(n15811),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i23_LC_12_15_2 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i23_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i23_LC_12_15_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i23_LC_12_15_2  (
            .in0(N__49237),
            .in1(N__41585),
            .in2(N__36793),
            .in3(N__48804),
            .lcout(cmd_rdadctmp_23_adj_1089),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51195),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i3_LC_12_15_3.C_ON=1'b0;
    defparam buf_device_acadc_i3_LC_12_15_3.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i3_LC_12_15_3.LUT_INIT=16'b0011101100001000;
    LogicCell40 buf_device_acadc_i3_LC_12_15_3 (
            .in0(N__34407),
            .in1(N__31869),
            .in2(N__51897),
            .in3(N__28554),
            .lcout(M_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51195),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i9_LC_12_15_5 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i9_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i9_LC_12_15_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i9_LC_12_15_5  (
            .in0(N__44331),
            .in1(N__49238),
            .in2(N__44549),
            .in3(N__42087),
            .lcout(buf_adcdata3_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51195),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.cmd_rdadctmp_i22_LC_12_15_6 .C_ON=1'b0;
    defparam \ADC_VAC4.cmd_rdadctmp_i22_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.cmd_rdadctmp_i22_LC_12_15_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC4.cmd_rdadctmp_i22_LC_12_15_6  (
            .in0(N__26416),
            .in1(N__27403),
            .in2(N__26388),
            .in3(N__26753),
            .lcout(cmd_rdadctmp_22_adj_1127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51195),
            .ce(),
            .sr(_gnd_net_));
    defparam i130_3_lut_adj_291_LC_12_15_7.C_ON=1'b0;
    defparam i130_3_lut_adj_291_LC_12_15_7.SEQ_MODE=4'b0000;
    defparam i130_3_lut_adj_291_LC_12_15_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 i130_3_lut_adj_291_LC_12_15_7 (
            .in0(N__26362),
            .in1(N__34888),
            .in2(_gnd_net_),
            .in3(N__47239),
            .lcout(n90),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.adc_state_i2_LC_12_16_1 .C_ON=1'b0;
    defparam \ADC_VAC4.adc_state_i2_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.adc_state_i2_LC_12_16_1 .LUT_INIT=16'b0110011000100010;
    LogicCell40 \ADC_VAC4.adc_state_i2_LC_12_16_1  (
            .in0(N__27023),
            .in1(N__27097),
            .in2(_gnd_net_),
            .in3(N__27230),
            .lcout(DTRIG_N_957_adj_1150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51212),
            .ce(N__26962),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_218_LC_12_16_2.C_ON=1'b0;
    defparam i1_2_lut_adj_218_LC_12_16_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_218_LC_12_16_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 i1_2_lut_adj_218_LC_12_16_2 (
            .in0(N__27096),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27022),
            .lcout(n15156),
            .ltout(n15156_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i1_3_lut_adj_9_LC_12_16_3 .C_ON=1'b0;
    defparam \ADC_VAC4.i1_3_lut_adj_9_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i1_3_lut_adj_9_LC_12_16_3 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \ADC_VAC4.i1_3_lut_adj_9_LC_12_16_3  (
            .in0(N__26657),
            .in1(_gnd_net_),
            .in2(N__26861),
            .in3(N__27229),
            .lcout(n9694),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i18_3_lut_LC_12_16_5 .C_ON=1'b0;
    defparam \ADC_VAC4.i18_3_lut_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i18_3_lut_LC_12_16_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ADC_VAC4.i18_3_lut_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__27095),
            .in2(N__26664),
            .in3(N__30636),
            .lcout(\ADC_VAC4.n15278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i1_4_lut_adj_8_LC_12_17_1 .C_ON=1'b0;
    defparam \ADC_VAC4.i1_4_lut_adj_8_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i1_4_lut_adj_8_LC_12_17_1 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \ADC_VAC4.i1_4_lut_adj_8_LC_12_17_1  (
            .in0(N__27235),
            .in1(N__26637),
            .in2(N__27114),
            .in3(N__30648),
            .lcout(),
            .ltout(\ADC_VAC4.n15257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i1_2_lut_LC_12_17_2 .C_ON=1'b0;
    defparam \ADC_VAC4.i1_2_lut_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i1_2_lut_LC_12_17_2 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \ADC_VAC4.i1_2_lut_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26684),
            .in3(N__27018),
            .lcout(\ADC_VAC4.n15258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i1_3_lut_LC_12_17_3 .C_ON=1'b0;
    defparam \ADC_VAC4.i1_3_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i1_3_lut_LC_12_17_3 .LUT_INIT=16'b1010000010101010;
    LogicCell40 \ADC_VAC4.i1_3_lut_LC_12_17_3  (
            .in0(N__27017),
            .in1(_gnd_net_),
            .in2(N__27322),
            .in3(N__26675),
            .lcout(\ADC_VAC4.n14930 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_198_LC_12_17_4.C_ON=1'b0;
    defparam i1_4_lut_adj_198_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_198_LC_12_17_4.LUT_INIT=16'b0000111100000110;
    LogicCell40 i1_4_lut_adj_198_LC_12_17_4 (
            .in0(N__27104),
            .in1(N__27236),
            .in2(N__26581),
            .in3(N__27016),
            .lcout(),
            .ltout(n14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.CS_37_LC_12_17_5 .C_ON=1'b0;
    defparam \ADC_VAC4.CS_37_LC_12_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.CS_37_LC_12_17_5 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \ADC_VAC4.CS_37_LC_12_17_5  (
            .in0(N__27237),
            .in1(N__26636),
            .in2(N__26606),
            .in3(N__26603),
            .lcout(M_CS4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51229),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1457_i4_4_lut_LC_12_17_6.C_ON=1'b0;
    defparam mux_1457_i4_4_lut_LC_12_17_6.SEQ_MODE=4'b0000;
    defparam mux_1457_i4_4_lut_LC_12_17_6.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1457_i4_4_lut_LC_12_17_6 (
            .in0(N__26564),
            .in1(N__47944),
            .in2(N__26548),
            .in3(N__47310),
            .lcout(n4061),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.i13062_2_lut_LC_12_17_7 .C_ON=1'b0;
    defparam \ADC_VAC4.i13062_2_lut_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC4.i13062_2_lut_LC_12_17_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \ADC_VAC4.i13062_2_lut_LC_12_17_7  (
            .in0(N__27234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26498),
            .lcout(\ADC_VAC4.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC4.adc_state_i1_LC_12_18_0 .C_ON=1'b0;
    defparam \ADC_VAC4.adc_state_i1_LC_12_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC4.adc_state_i1_LC_12_18_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \ADC_VAC4.adc_state_i1_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__27252),
            .in2(_gnd_net_),
            .in3(N__27113),
            .lcout(adc_state_1_adj_1116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51245),
            .ce(N__26963),
            .sr(N__26948));
    defparam CONSTANT_ONE_LUT4_LC_13_1_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_1_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_1_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i4_7360_7361_set_LC_13_3_3 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_7360_7361_set_LC_13_3_3 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i4_7360_7361_set_LC_13_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_7360_7361_set_LC_13_3_3  (
            .in0(N__29029),
            .in1(N__26939),
            .in2(_gnd_net_),
            .in3(N__26927),
            .lcout(\comm_spi.n10471 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42460),
            .ce(),
            .sr(N__46655));
    defparam \comm_spi.data_tx_i4_7360_7361_reset_LC_13_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_7360_7361_reset_LC_13_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i4_7360_7361_reset_LC_13_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_7360_7361_reset_LC_13_4_0  (
            .in0(N__29030),
            .in1(N__26938),
            .in2(_gnd_net_),
            .in3(N__26923),
            .lcout(\comm_spi.n10472 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42462),
            .ce(),
            .sr(N__26912));
    defparam \comm_spi.i13077_4_lut_3_lut_LC_13_5_0 .C_ON=1'b0;
    defparam \comm_spi.i13077_4_lut_3_lut_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13077_4_lut_3_lut_LC_13_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i13077_4_lut_3_lut_LC_13_5_0  (
            .in0(N__26877),
            .in1(N__30835),
            .in2(_gnd_net_),
            .in3(N__46575),
            .lcout(\comm_spi.n10444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.CS_28_LC_13_5_2 .C_ON=1'b0;
    defparam \CLOCK_DDS.CS_28_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.CS_28_LC_13_5_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \CLOCK_DDS.CS_28_LC_13_5_2  (
            .in0(N__35746),
            .in1(N__48388),
            .in2(_gnd_net_),
            .in3(N__48537),
            .lcout(DDS_CS1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51110),
            .ce(N__31166),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_13_5_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_13_5_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_100_2_lut_LC_13_5_3  (
            .in0(N__46576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26878),
            .lcout(\comm_spi.data_tx_7__N_813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_13_5_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_13_5_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_92_2_lut_LC_13_5_4  (
            .in0(N__26879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46574),
            .lcout(\comm_spi.data_tx_7__N_805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_5_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_5_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \comm_spi.RESET_I_0_101_2_lut_LC_13_5_5  (
            .in0(N__46577),
            .in1(N__27687),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_5_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_93_2_lut_LC_13_5_6  (
            .in0(N__27688),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46578),
            .lcout(\comm_spi.data_tx_7__N_806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13112_4_lut_3_lut_LC_13_5_7 .C_ON=1'b0;
    defparam \comm_spi.i13112_4_lut_3_lut_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13112_4_lut_3_lut_LC_13_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i13112_4_lut_3_lut_LC_13_5_7  (
            .in0(N__46579),
            .in1(N__27689),
            .in2(_gnd_net_),
            .in3(N__27657),
            .lcout(\comm_spi.n16884 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i7_7337_7338_reset_LC_13_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_7337_7338_reset_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i7_7337_7338_reset_LC_13_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_7337_7338_reset_LC_13_6_0  (
            .in0(N__27658),
            .in1(N__27787),
            .in2(_gnd_net_),
            .in3(N__28984),
            .lcout(\comm_spi.n10449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42461),
            .ce(),
            .sr(N__30996));
    defparam i1_2_lut_adj_289_LC_13_7_0.C_ON=1'b0;
    defparam i1_2_lut_adj_289_LC_13_7_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_289_LC_13_7_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_289_LC_13_7_0 (
            .in0(_gnd_net_),
            .in1(N__47989),
            .in2(_gnd_net_),
            .in3(N__45298),
            .lcout(),
            .ltout(n18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12648_4_lut_LC_13_7_1.C_ON=1'b0;
    defparam i12648_4_lut_LC_13_7_1.SEQ_MODE=4'b0000;
    defparam i12648_4_lut_LC_13_7_1.LUT_INIT=16'b1011000010000000;
    LogicCell40 i12648_4_lut_LC_13_7_1 (
            .in0(N__27641),
            .in1(N__45650),
            .in2(N__27623),
            .in3(N__29513),
            .lcout(),
            .ltout(n15466_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i103_4_lut_LC_13_7_2.C_ON=1'b0;
    defparam i103_4_lut_LC_13_7_2.SEQ_MODE=4'b0000;
    defparam i103_4_lut_LC_13_7_2.LUT_INIT=16'b1111000001000100;
    LogicCell40 i103_4_lut_LC_13_7_2 (
            .in0(N__45651),
            .in1(N__27599),
            .in2(N__27620),
            .in3(N__47085),
            .lcout(n104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i110_4_lut_LC_13_7_3.C_ON=1'b0;
    defparam i110_4_lut_LC_13_7_3.SEQ_MODE=4'b0000;
    defparam i110_4_lut_LC_13_7_3.LUT_INIT=16'b0101100000001000;
    LogicCell40 i110_4_lut_LC_13_7_3 (
            .in0(N__45297),
            .in1(N__29360),
            .in2(N__48046),
            .in3(N__31460),
            .lcout(n56),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1481_i2_4_lut_LC_13_7_5.C_ON=1'b0;
    defparam mux_1481_i2_4_lut_LC_13_7_5.SEQ_MODE=4'b0000;
    defparam mux_1481_i2_4_lut_LC_13_7_5.LUT_INIT=16'b1010111000000100;
    LogicCell40 mux_1481_i2_4_lut_LC_13_7_5 (
            .in0(N__47086),
            .in1(N__27586),
            .in2(N__48047),
            .in3(N__27557),
            .lcout(n4151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12765_2_lut_3_lut_4_lut_LC_13_7_6.C_ON=1'b0;
    defparam i12765_2_lut_3_lut_4_lut_LC_13_7_6.SEQ_MODE=4'b0000;
    defparam i12765_2_lut_3_lut_4_lut_LC_13_7_6.LUT_INIT=16'b0000010000000000;
    LogicCell40 i12765_2_lut_3_lut_4_lut_LC_13_7_6 (
            .in0(N__33116),
            .in1(N__38832),
            .in2(N__33329),
            .in3(N__27860),
            .lcout(),
            .ltout(n15567_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i22_4_lut_adj_232_LC_13_7_7.C_ON=1'b0;
    defparam i22_4_lut_adj_232_LC_13_7_7.SEQ_MODE=4'b0000;
    defparam i22_4_lut_adj_232_LC_13_7_7.LUT_INIT=16'b1101010110000000;
    LogicCell40 i22_4_lut_adj_232_LC_13_7_7 (
            .in0(N__50321),
            .in1(N__33487),
            .in2(N__27737),
            .in3(N__33632),
            .lcout(n7_adj_1255),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_196_LC_13_8_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_196_LC_13_8_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_196_LC_13_8_0.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_adj_196_LC_13_8_0 (
            .in0(N__43450),
            .in1(N__39256),
            .in2(_gnd_net_),
            .in3(N__43238),
            .lcout(n5_adj_1235),
            .ltout(n5_adj_1235_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12752_4_lut_LC_13_8_1.C_ON=1'b0;
    defparam i12752_4_lut_LC_13_8_1.SEQ_MODE=4'b0000;
    defparam i12752_4_lut_LC_13_8_1.LUT_INIT=16'b0001000000000000;
    LogicCell40 i12752_4_lut_LC_13_8_1 (
            .in0(N__27722),
            .in1(N__33117),
            .in2(N__27716),
            .in3(N__38763),
            .lcout(),
            .ltout(n15535_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i30_4_lut_adj_265_LC_13_8_2.C_ON=1'b0;
    defparam i30_4_lut_adj_265_LC_13_8_2.SEQ_MODE=4'b0000;
    defparam i30_4_lut_adj_265_LC_13_8_2.LUT_INIT=16'b1011000110100000;
    LogicCell40 i30_4_lut_adj_265_LC_13_8_2 (
            .in0(N__49880),
            .in1(N__43643),
            .in2(N__27713),
            .in3(N__41936),
            .lcout(),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_178_LC_13_8_3.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_178_LC_13_8_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_178_LC_13_8_3.LUT_INIT=16'b1110101001000000;
    LogicCell40 i1_4_lut_4_lut_adj_178_LC_13_8_3 (
            .in0(N__52380),
            .in1(N__31123),
            .in2(N__27710),
            .in3(N__51898),
            .lcout(n9021),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i6_LC_13_8_5.C_ON=1'b0;
    defparam data_index_i6_LC_13_8_5.SEQ_MODE=4'b1000;
    defparam data_index_i6_LC_13_8_5.LUT_INIT=16'b0111010100100000;
    LogicCell40 data_index_i6_LC_13_8_5 (
            .in0(N__52384),
            .in1(N__51899),
            .in2(N__30410),
            .in3(N__30431),
            .lcout(data_index_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51122),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_3_lut_4_lut_LC_13_8_7.C_ON=1'b0;
    defparam i1_3_lut_3_lut_4_lut_LC_13_8_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_3_lut_4_lut_LC_13_8_7.LUT_INIT=16'b1111010011000010;
    LogicCell40 i1_3_lut_3_lut_4_lut_LC_13_8_7 (
            .in0(N__50582),
            .in1(N__49479),
            .in2(N__52454),
            .in3(N__49881),
            .lcout(n8561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i2_LC_13_9_0.C_ON=1'b0;
    defparam comm_index_i2_LC_13_9_0.SEQ_MODE=4'b1000;
    defparam comm_index_i2_LC_13_9_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 comm_index_i2_LC_13_9_0 (
            .in0(N__33415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27695),
            .lcout(comm_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51130),
            .ce(N__32518),
            .sr(N__33704));
    defparam i1704_2_lut_3_lut_4_lut_LC_13_9_1.C_ON=1'b0;
    defparam i1704_2_lut_3_lut_4_lut_LC_13_9_1.SEQ_MODE=4'b0000;
    defparam i1704_2_lut_3_lut_4_lut_LC_13_9_1.LUT_INIT=16'b0010000000000000;
    LogicCell40 i1704_2_lut_3_lut_4_lut_LC_13_9_1 (
            .in0(N__38831),
            .in1(N__43454),
            .in2(N__33169),
            .in3(N__43281),
            .lcout(n4814),
            .ltout(n4814_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i3_LC_13_9_2.C_ON=1'b0;
    defparam comm_index_i3_LC_13_9_2.SEQ_MODE=4'b1000;
    defparam comm_index_i3_LC_13_9_2.LUT_INIT=16'b0101101010101010;
    LogicCell40 comm_index_i3_LC_13_9_2 (
            .in0(N__33251),
            .in1(_gnd_net_),
            .in2(N__27866),
            .in3(N__33448),
            .lcout(comm_index_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51130),
            .ce(N__32518),
            .sr(N__33704));
    defparam i1_2_lut_3_lut_adj_261_LC_13_9_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_261_LC_13_9_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_261_LC_13_9_3.LUT_INIT=16'b0000000000110000;
    LogicCell40 i1_2_lut_3_lut_adj_261_LC_13_9_3 (
            .in0(_gnd_net_),
            .in1(N__33414),
            .in2(N__27863),
            .in3(N__33250),
            .lcout(n13475),
            .ltout(n13475_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12972_2_lut_LC_13_9_4.C_ON=1'b0;
    defparam i12972_2_lut_LC_13_9_4.SEQ_MODE=4'b0000;
    defparam i12972_2_lut_LC_13_9_4.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12972_2_lut_LC_13_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27833),
            .in3(N__33111),
            .lcout(),
            .ltout(n15802_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i30_4_lut_LC_13_9_5.C_ON=1'b0;
    defparam i30_4_lut_LC_13_9_5.SEQ_MODE=4'b0000;
    defparam i30_4_lut_LC_13_9_5.LUT_INIT=16'b1011001110000000;
    LogicCell40 i30_4_lut_LC_13_9_5 (
            .in0(N__38830),
            .in1(N__50202),
            .in2(N__27830),
            .in3(N__33627),
            .lcout(n10_adj_1249),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12743_2_lut_LC_13_9_6.C_ON=1'b0;
    defparam i12743_2_lut_LC_13_9_6.SEQ_MODE=4'b0000;
    defparam i12743_2_lut_LC_13_9_6.LUT_INIT=16'b0011001100000000;
    LogicCell40 i12743_2_lut_LC_13_9_6 (
            .in0(_gnd_net_),
            .in1(N__38829),
            .in2(_gnd_net_),
            .in3(N__31073),
            .lcout(),
            .ltout(n15657_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i33_4_lut_LC_13_9_7.C_ON=1'b0;
    defparam i33_4_lut_LC_13_9_7.SEQ_MODE=4'b0000;
    defparam i33_4_lut_LC_13_9_7.LUT_INIT=16'b1011001110000000;
    LogicCell40 i33_4_lut_LC_13_9_7 (
            .in0(N__33112),
            .in1(N__50203),
            .in2(N__27812),
            .in3(N__33628),
            .lcout(n13_adj_1042),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_7368_7369_set_LC_13_10_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_7368_7369_set_LC_13_10_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i6_7368_7369_set_LC_13_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_7368_7369_set_LC_13_10_0  (
            .in0(N__28907),
            .in1(N__28934),
            .in2(_gnd_net_),
            .in3(N__29012),
            .lcout(\comm_spi.n10479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42438),
            .ce(),
            .sr(N__27770));
    defparam i12661_2_lut_LC_13_10_1.C_ON=1'b0;
    defparam i12661_2_lut_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam i12661_2_lut_LC_13_10_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12661_2_lut_LC_13_10_1 (
            .in0(_gnd_net_),
            .in1(N__41863),
            .in2(_gnd_net_),
            .in3(N__32126),
            .lcout(n15576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12670_2_lut_LC_13_10_2.C_ON=1'b0;
    defparam i12670_2_lut_LC_13_10_2.SEQ_MODE=4'b0000;
    defparam i12670_2_lut_LC_13_10_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 i12670_2_lut_LC_13_10_2 (
            .in0(N__47914),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31805),
            .lcout(n15691),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12678_2_lut_LC_13_10_3.C_ON=1'b0;
    defparam i12678_2_lut_LC_13_10_3.SEQ_MODE=4'b0000;
    defparam i12678_2_lut_LC_13_10_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i12678_2_lut_LC_13_10_3 (
            .in0(_gnd_net_),
            .in1(N__27877),
            .in2(_gnd_net_),
            .in3(N__47915),
            .lcout(n15475),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12701_2_lut_LC_13_10_4.C_ON=1'b0;
    defparam i12701_2_lut_LC_13_10_4.SEQ_MODE=4'b0000;
    defparam i12701_2_lut_LC_13_10_4.LUT_INIT=16'b0100010001000100;
    LogicCell40 i12701_2_lut_LC_13_10_4 (
            .in0(N__47912),
            .in1(N__29489),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n15835),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12746_2_lut_LC_13_10_5.C_ON=1'b0;
    defparam i12746_2_lut_LC_13_10_5.SEQ_MODE=4'b0000;
    defparam i12746_2_lut_LC_13_10_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12746_2_lut_LC_13_10_5 (
            .in0(_gnd_net_),
            .in1(N__33851),
            .in2(_gnd_net_),
            .in3(N__47911),
            .lcout(n15542),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12851_2_lut_LC_13_10_6.C_ON=1'b0;
    defparam i12851_2_lut_LC_13_10_6.SEQ_MODE=4'b0000;
    defparam i12851_2_lut_LC_13_10_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12851_2_lut_LC_13_10_6 (
            .in0(N__47913),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29545),
            .lcout(n15679),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12713_2_lut_LC_13_11_0.C_ON=1'b0;
    defparam i12713_2_lut_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam i12713_2_lut_LC_13_11_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 i12713_2_lut_LC_13_11_0 (
            .in0(_gnd_net_),
            .in1(N__28065),
            .in2(_gnd_net_),
            .in3(N__47916),
            .lcout(n15543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i130_3_lut_LC_13_11_1.C_ON=1'b0;
    defparam i130_3_lut_LC_13_11_1.SEQ_MODE=4'b0000;
    defparam i130_3_lut_LC_13_11_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i130_3_lut_LC_13_11_1 (
            .in0(N__27955),
            .in1(N__34856),
            .in2(_gnd_net_),
            .in3(N__47138),
            .lcout(),
            .ltout(n90_adj_1023_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i127_4_lut_LC_13_11_2.C_ON=1'b0;
    defparam i127_4_lut_LC_13_11_2.SEQ_MODE=4'b0000;
    defparam i127_4_lut_LC_13_11_2.LUT_INIT=16'b1111000010001000;
    LogicCell40 i127_4_lut_LC_13_11_2 (
            .in0(N__47139),
            .in1(N__27925),
            .in2(N__27896),
            .in3(N__45639),
            .lcout(n69_adj_1113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i123_3_lut_LC_13_11_3.C_ON=1'b0;
    defparam i123_3_lut_LC_13_11_3.SEQ_MODE=4'b0000;
    defparam i123_3_lut_LC_13_11_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i123_3_lut_LC_13_11_3 (
            .in0(N__28535),
            .in1(N__34154),
            .in2(_gnd_net_),
            .in3(N__47137),
            .lcout(n96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i5_LC_13_11_4.C_ON=1'b0;
    defparam buf_device_acadc_i5_LC_13_11_4.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i5_LC_13_11_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_device_acadc_i5_LC_13_11_4 (
            .in0(N__31846),
            .in1(N__36994),
            .in2(N__51770),
            .in3(N__27878),
            .lcout(buf_device_acadc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51153),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i1_LC_13_11_5.C_ON=1'b0;
    defparam buf_device_acadc_i1_LC_13_11_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i1_LC_13_11_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 buf_device_acadc_i1_LC_13_11_5 (
            .in0(N__28066),
            .in1(N__37272),
            .in2(_gnd_net_),
            .in3(N__31847),
            .lcout(M_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51153),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i15_LC_13_11_7.C_ON=1'b0;
    defparam req_data_cnt_i15_LC_13_11_7.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i15_LC_13_11_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i15_LC_13_11_7 (
            .in0(N__37583),
            .in1(N__40457),
            .in2(_gnd_net_),
            .in3(N__29511),
            .lcout(req_data_cnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51153),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_13_12_0.C_ON=1'b0;
    defparam i1_2_lut_LC_13_12_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_13_12_0.LUT_INIT=16'b0000000010101010;
    LogicCell40 i1_2_lut_LC_13_12_0 (
            .in0(N__52345),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50596),
            .lcout(n8062),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12984_2_lut_LC_13_12_1.C_ON=1'b0;
    defparam i12984_2_lut_LC_13_12_1.SEQ_MODE=4'b0000;
    defparam i12984_2_lut_LC_13_12_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12984_2_lut_LC_13_12_1 (
            .in0(_gnd_net_),
            .in1(N__47909),
            .in2(_gnd_net_),
            .in3(N__41708),
            .lcout(n15555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_49_LC_13_12_2.C_ON=1'b0;
    defparam i1_2_lut_adj_49_LC_13_12_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_49_LC_13_12_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_49_LC_13_12_2 (
            .in0(_gnd_net_),
            .in1(N__32877),
            .in2(_gnd_net_),
            .in3(N__38090),
            .lcout(n3),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_280_LC_13_12_3.C_ON=1'b0;
    defparam i1_4_lut_adj_280_LC_13_12_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_280_LC_13_12_3.LUT_INIT=16'b1111111000000000;
    LogicCell40 i1_4_lut_adj_280_LC_13_12_3 (
            .in0(N__32809),
            .in1(N__32736),
            .in2(N__28040),
            .in3(N__28028),
            .lcout(),
            .ltout(n10_adj_1242_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_end_328_LC_13_12_4.C_ON=1'b0;
    defparam eis_end_328_LC_13_12_4.SEQ_MODE=4'b1000;
    defparam eis_end_328_LC_13_12_4.LUT_INIT=16'b1111010011110000;
    LogicCell40 eis_end_328_LC_13_12_4 (
            .in0(N__32735),
            .in1(N__38092),
            .in2(N__28037),
            .in3(N__28034),
            .lcout(eis_end),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_end_328C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i3_3_lut_LC_13_12_5.C_ON=1'b0;
    defparam mux_1502_i3_3_lut_LC_13_12_5.SEQ_MODE=4'b0000;
    defparam mux_1502_i3_3_lut_LC_13_12_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_1502_i3_3_lut_LC_13_12_5 (
            .in0(N__31946),
            .in1(N__40325),
            .in2(_gnd_net_),
            .in3(N__47910),
            .lcout(n4219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_149_LC_13_12_6.C_ON=1'b0;
    defparam i1_2_lut_adj_149_LC_13_12_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_149_LC_13_12_6.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_149_LC_13_12_6 (
            .in0(_gnd_net_),
            .in1(N__32808),
            .in2(_gnd_net_),
            .in3(N__38091),
            .lcout(n15171),
            .ltout(n15171_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_3_lut_LC_13_12_7.C_ON=1'b0;
    defparam i2_3_lut_3_lut_LC_13_12_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_3_lut_LC_13_12_7.LUT_INIT=16'b0000000010100000;
    LogicCell40 i2_3_lut_3_lut_LC_13_12_7 (
            .in0(N__32878),
            .in1(_gnd_net_),
            .in2(N__28016),
            .in3(N__32737),
            .lcout(raw_buf1_N_775),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i0_LC_13_13_0.C_ON=1'b0;
    defparam eis_state_i0_LC_13_13_0.SEQ_MODE=4'b1010;
    defparam eis_state_i0_LC_13_13_0.LUT_INIT=16'b1000100010001101;
    LogicCell40 eis_state_i0_LC_13_13_0 (
            .in0(N__32813),
            .in1(N__28508),
            .in2(N__32916),
            .in3(N__29699),
            .lcout(eis_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__28187),
            .sr(N__32753));
    defparam i17_4_lut_LC_13_13_1.C_ON=1'b0;
    defparam i17_4_lut_LC_13_13_1.SEQ_MODE=4'b0000;
    defparam i17_4_lut_LC_13_13_1.LUT_INIT=16'b1110111111100000;
    LogicCell40 i17_4_lut_LC_13_13_1 (
            .in0(N__41037),
            .in1(N__34508),
            .in2(N__32923),
            .in3(N__28225),
            .lcout(),
            .ltout(n15356_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13047_3_lut_LC_13_13_2.C_ON=1'b0;
    defparam i13047_3_lut_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam i13047_3_lut_LC_13_13_2.LUT_INIT=16'b0011111111111111;
    LogicCell40 i13047_3_lut_LC_13_13_2 (
            .in0(_gnd_net_),
            .in1(N__32810),
            .in2(N__28208),
            .in3(N__38095),
            .lcout(n8459),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12862_2_lut_LC_13_13_3.C_ON=1'b0;
    defparam i12862_2_lut_LC_13_13_3.SEQ_MODE=4'b0000;
    defparam i12862_2_lut_LC_13_13_3.LUT_INIT=16'b0101010100000000;
    LogicCell40 i12862_2_lut_LC_13_13_3 (
            .in0(N__32911),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28522),
            .lcout(),
            .ltout(n15695_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i2_LC_13_13_4.C_ON=1'b0;
    defparam eis_state_i2_LC_13_13_4.SEQ_MODE=4'b1010;
    defparam eis_state_i2_LC_13_13_4.LUT_INIT=16'b1110011010100010;
    LogicCell40 eis_state_i2_LC_13_13_4 (
            .in0(N__32814),
            .in1(N__38096),
            .in2(N__28205),
            .in3(N__28202),
            .lcout(eis_end_N_770),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__28187),
            .sr(N__32753));
    defparam i12861_3_lut_LC_13_13_5.C_ON=1'b0;
    defparam i12861_3_lut_LC_13_13_5.SEQ_MODE=4'b0000;
    defparam i12861_3_lut_LC_13_13_5.LUT_INIT=16'b1111111111110101;
    LogicCell40 i12861_3_lut_LC_13_13_5 (
            .in0(N__41038),
            .in1(_gnd_net_),
            .in2(N__32924),
            .in3(N__29710),
            .lcout(n15696),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12776_2_lut_3_lut_LC_13_13_6.C_ON=1'b0;
    defparam i12776_2_lut_3_lut_LC_13_13_6.SEQ_MODE=4'b0000;
    defparam i12776_2_lut_3_lut_LC_13_13_6.LUT_INIT=16'b0100010000000000;
    LogicCell40 i12776_2_lut_3_lut_LC_13_13_6 (
            .in0(N__29711),
            .in1(N__38094),
            .in2(_gnd_net_),
            .in3(N__41039),
            .lcout(),
            .ltout(n15700_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i1_LC_13_13_7.C_ON=1'b0;
    defparam eis_state_i1_LC_13_13_7.SEQ_MODE=4'b1010;
    defparam eis_state_i1_LC_13_13_7.LUT_INIT=16'b0101010011111110;
    LogicCell40 eis_state_i1_LC_13_13_7 (
            .in0(N__32811),
            .in1(N__32899),
            .in2(N__28196),
            .in3(N__28193),
            .lcout(eis_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__28187),
            .sr(N__32753));
    defparam comm_state_3__I_0_394_Mux_4_i15_4_lut_LC_13_14_0.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_4_i15_4_lut_LC_13_14_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_4_i15_4_lut_LC_13_14_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_394_Mux_4_i15_4_lut_LC_13_14_0 (
            .in0(N__52430),
            .in1(N__28501),
            .in2(N__51766),
            .in3(N__29887),
            .lcout(data_index_9_N_258_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_end_I_3_3_lut_LC_13_14_1.C_ON=1'b0;
    defparam eis_end_I_3_3_lut_LC_13_14_1.SEQ_MODE=4'b0000;
    defparam eis_end_I_3_3_lut_LC_13_14_1.LUT_INIT=16'b1010101010111011;
    LogicCell40 eis_end_I_3_3_lut_LC_13_14_1 (
            .in0(N__34502),
            .in1(N__29459),
            .in2(_gnd_net_),
            .in3(N__31742),
            .lcout(eis_end_N_773),
            .ltout(eis_end_N_773_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12717_3_lut_LC_13_14_2.C_ON=1'b0;
    defparam i12717_3_lut_LC_13_14_2.SEQ_MODE=4'b0000;
    defparam i12717_3_lut_LC_13_14_2.LUT_INIT=16'b1010101010100000;
    LogicCell40 i12717_3_lut_LC_13_14_2 (
            .in0(N__38097),
            .in1(_gnd_net_),
            .in2(N__28511),
            .in3(N__32889),
            .lcout(n15510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i4_LC_13_14_3.C_ON=1'b0;
    defparam acadc_skipCount_i4_LC_13_14_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i4_LC_13_14_3.LUT_INIT=16'b0111010100100000;
    LogicCell40 acadc_skipCount_i4_LC_13_14_3 (
            .in0(N__41826),
            .in1(N__51668),
            .in2(N__31625),
            .in3(N__31885),
            .lcout(acadc_skipCount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51202),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i2_LC_13_14_4.C_ON=1'b0;
    defparam buf_device_acadc_i2_LC_13_14_4.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i2_LC_13_14_4.LUT_INIT=16'b0011101100001000;
    LogicCell40 buf_device_acadc_i2_LC_13_14_4 (
            .in0(N__34593),
            .in1(N__31862),
            .in2(N__51767),
            .in3(N__29424),
            .lcout(M_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51202),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i1_LC_13_14_5.C_ON=1'b0;
    defparam acadc_skipCount_i1_LC_13_14_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i1_LC_13_14_5.LUT_INIT=16'b0101000011011000;
    LogicCell40 acadc_skipCount_i1_LC_13_14_5 (
            .in0(N__41825),
            .in1(N__41101),
            .in2(N__42187),
            .in3(N__51675),
            .lcout(acadc_skipCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51202),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i4_LC_13_14_6.C_ON=1'b0;
    defparam data_index_i4_LC_13_14_6.SEQ_MODE=4'b1000;
    defparam data_index_i4_LC_13_14_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i4_LC_13_14_6 (
            .in0(N__52431),
            .in1(N__28502),
            .in2(N__51768),
            .in3(N__29888),
            .lcout(data_index_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51202),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_69_LC_13_14_7.C_ON=1'b0;
    defparam i2_4_lut_adj_69_LC_13_14_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_69_LC_13_14_7.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_69_LC_13_14_7 (
            .in0(N__28679),
            .in1(N__31884),
            .in2(N__28655),
            .in3(N__42177),
            .lcout(n18_adj_1276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i24_LC_13_15_1 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i24_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i24_LC_13_15_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i24_LC_13_15_1  (
            .in0(N__36789),
            .in1(N__49239),
            .in2(N__28483),
            .in3(N__48803),
            .lcout(cmd_rdadctmp_24_adj_1088),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51219),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_1_i15_4_lut_LC_13_15_3.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_1_i15_4_lut_LC_13_15_3.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_1_i15_4_lut_LC_13_15_3.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_394_Mux_1_i15_4_lut_LC_13_15_3 (
            .in0(N__52434),
            .in1(N__28577),
            .in2(N__51829),
            .in3(N__29959),
            .lcout(data_index_9_N_258_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1457_i6_4_lut_LC_13_15_4.C_ON=1'b0;
    defparam mux_1457_i6_4_lut_LC_13_15_4.SEQ_MODE=4'b0000;
    defparam mux_1457_i6_4_lut_LC_13_15_4.LUT_INIT=16'b1100010111000000;
    LogicCell40 mux_1457_i6_4_lut_LC_13_15_4 (
            .in0(N__47860),
            .in1(N__28628),
            .in2(N__47307),
            .in3(N__28614),
            .lcout(n4059),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3209_3_lut_LC_13_15_5.C_ON=1'b0;
    defparam i3209_3_lut_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam i3209_3_lut_LC_13_15_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 i3209_3_lut_LC_13_15_5 (
            .in0(N__41092),
            .in1(N__29978),
            .in2(_gnd_net_),
            .in3(N__40544),
            .lcout(n8_adj_1233),
            .ltout(n8_adj_1233_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i1_LC_13_15_6.C_ON=1'b0;
    defparam data_index_i1_LC_13_15_6.SEQ_MODE=4'b1000;
    defparam data_index_i1_LC_13_15_6.LUT_INIT=16'b0010001011100010;
    LogicCell40 data_index_i1_LC_13_15_6 (
            .in0(N__29960),
            .in1(N__52435),
            .in2(N__28571),
            .in3(N__51725),
            .lcout(data_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51219),
            .ce(),
            .sr(_gnd_net_));
    defparam i132_4_lut_LC_13_15_7.C_ON=1'b0;
    defparam i132_4_lut_LC_13_15_7.SEQ_MODE=4'b0000;
    defparam i132_4_lut_LC_13_15_7.LUT_INIT=16'b0011000010001000;
    LogicCell40 i132_4_lut_LC_13_15_7 (
            .in0(N__34348),
            .in1(N__47859),
            .in2(N__28558),
            .in3(N__45294),
            .lcout(n66_adj_1166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i0_LC_13_16_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i0_LC_13_16_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i0_LC_13_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i0_LC_13_16_0 (
            .in0(_gnd_net_),
            .in1(N__29755),
            .in2(_gnd_net_),
            .in3(N__28526),
            .lcout(acadc_skipcnt_0),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(n13966),
            .clk(INVacadc_skipcnt_i0_i0C_net),
            .ce(N__32367),
            .sr(N__30686));
    defparam add_58_2_THRU_CRY_0_LC_13_16_1.C_ON=1'b1;
    defparam add_58_2_THRU_CRY_0_LC_13_16_1.SEQ_MODE=4'b0000;
    defparam add_58_2_THRU_CRY_0_LC_13_16_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_58_2_THRU_CRY_0_LC_13_16_1 (
            .in0(_gnd_net_),
            .in1(N__28767),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n13966),
            .carryout(n13966_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_58_2_THRU_CRY_1_LC_13_16_2.C_ON=1'b1;
    defparam add_58_2_THRU_CRY_1_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam add_58_2_THRU_CRY_1_LC_13_16_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_58_2_THRU_CRY_1_LC_13_16_2 (
            .in0(_gnd_net_),
            .in1(N__28771),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n13966_THRU_CRY_0_THRU_CO),
            .carryout(n13966_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_58_2_THRU_CRY_2_LC_13_16_3.C_ON=1'b1;
    defparam add_58_2_THRU_CRY_2_LC_13_16_3.SEQ_MODE=4'b0000;
    defparam add_58_2_THRU_CRY_2_LC_13_16_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_58_2_THRU_CRY_2_LC_13_16_3 (
            .in0(_gnd_net_),
            .in1(N__28768),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n13966_THRU_CRY_1_THRU_CO),
            .carryout(n13966_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_58_2_THRU_CRY_3_LC_13_16_4.C_ON=1'b1;
    defparam add_58_2_THRU_CRY_3_LC_13_16_4.SEQ_MODE=4'b0000;
    defparam add_58_2_THRU_CRY_3_LC_13_16_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_58_2_THRU_CRY_3_LC_13_16_4 (
            .in0(_gnd_net_),
            .in1(N__28772),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n13966_THRU_CRY_2_THRU_CO),
            .carryout(n13966_THRU_CRY_3_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_58_2_THRU_CRY_4_LC_13_16_5.C_ON=1'b1;
    defparam add_58_2_THRU_CRY_4_LC_13_16_5.SEQ_MODE=4'b0000;
    defparam add_58_2_THRU_CRY_4_LC_13_16_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_58_2_THRU_CRY_4_LC_13_16_5 (
            .in0(_gnd_net_),
            .in1(N__28769),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n13966_THRU_CRY_3_THRU_CO),
            .carryout(n13966_THRU_CRY_4_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_58_2_THRU_CRY_5_LC_13_16_6.C_ON=1'b1;
    defparam add_58_2_THRU_CRY_5_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam add_58_2_THRU_CRY_5_LC_13_16_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_58_2_THRU_CRY_5_LC_13_16_6 (
            .in0(_gnd_net_),
            .in1(N__28773),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n13966_THRU_CRY_4_THRU_CO),
            .carryout(n13966_THRU_CRY_5_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_58_2_THRU_CRY_6_LC_13_16_7.C_ON=1'b1;
    defparam add_58_2_THRU_CRY_6_LC_13_16_7.SEQ_MODE=4'b0000;
    defparam add_58_2_THRU_CRY_6_LC_13_16_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_58_2_THRU_CRY_6_LC_13_16_7 (
            .in0(_gnd_net_),
            .in1(N__28770),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n13966_THRU_CRY_5_THRU_CO),
            .carryout(n13966_THRU_CRY_6_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i1_LC_13_17_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i1_LC_13_17_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i1_LC_13_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i1_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(N__28678),
            .in2(_gnd_net_),
            .in3(N__28664),
            .lcout(acadc_skipcnt_1),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(n13967),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i2_LC_13_17_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i2_LC_13_17_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i2_LC_13_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i2_LC_13_17_1 (
            .in0(_gnd_net_),
            .in1(N__32005),
            .in2(_gnd_net_),
            .in3(N__28661),
            .lcout(acadc_skipcnt_2),
            .ltout(),
            .carryin(n13967),
            .carryout(n13968),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i3_LC_13_17_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i3_LC_13_17_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i3_LC_13_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i3_LC_13_17_2 (
            .in0(_gnd_net_),
            .in1(N__32324),
            .in2(_gnd_net_),
            .in3(N__28658),
            .lcout(acadc_skipcnt_3),
            .ltout(),
            .carryin(n13968),
            .carryout(n13969),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i4_LC_13_17_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i4_LC_13_17_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i4_LC_13_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i4_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(N__28651),
            .in2(_gnd_net_),
            .in3(N__28637),
            .lcout(acadc_skipcnt_4),
            .ltout(),
            .carryin(n13969),
            .carryout(n13970),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i5_LC_13_17_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i5_LC_13_17_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i5_LC_13_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i5_LC_13_17_4 (
            .in0(_gnd_net_),
            .in1(N__32305),
            .in2(_gnd_net_),
            .in3(N__28634),
            .lcout(acadc_skipcnt_5),
            .ltout(),
            .carryin(n13970),
            .carryout(n13971),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i6_LC_13_17_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i6_LC_13_17_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i6_LC_13_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i6_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(N__29737),
            .in2(_gnd_net_),
            .in3(N__28631),
            .lcout(acadc_skipcnt_6),
            .ltout(),
            .carryin(n13971),
            .carryout(n13972),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i7_LC_13_17_6.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i7_LC_13_17_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i7_LC_13_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i7_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(N__31960),
            .in2(_gnd_net_),
            .in3(N__28880),
            .lcout(acadc_skipcnt_7),
            .ltout(),
            .carryin(n13972),
            .carryout(n13973),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i8_LC_13_17_7.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i8_LC_13_17_7.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i8_LC_13_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i8_LC_13_17_7 (
            .in0(_gnd_net_),
            .in1(N__32290),
            .in2(_gnd_net_),
            .in3(N__28877),
            .lcout(acadc_skipcnt_8),
            .ltout(),
            .carryin(n13973),
            .carryout(n13974),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__32371),
            .sr(N__30707));
    defparam acadc_skipcnt_i0_i9_LC_13_18_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i9_LC_13_18_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i9_LC_13_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i9_LC_13_18_0 (
            .in0(_gnd_net_),
            .in1(N__31507),
            .in2(_gnd_net_),
            .in3(N__28874),
            .lcout(acadc_skipcnt_9),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(n13975),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32375),
            .sr(N__30703));
    defparam acadc_skipcnt_i0_i10_LC_13_18_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i10_LC_13_18_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i10_LC_13_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i10_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(N__30076),
            .in2(_gnd_net_),
            .in3(N__28871),
            .lcout(acadc_skipcnt_10),
            .ltout(),
            .carryin(n13975),
            .carryout(n13976),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32375),
            .sr(N__30703));
    defparam acadc_skipcnt_i0_i11_LC_13_18_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i11_LC_13_18_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i11_LC_13_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i11_LC_13_18_2 (
            .in0(_gnd_net_),
            .in1(N__30121),
            .in2(_gnd_net_),
            .in3(N__28868),
            .lcout(acadc_skipcnt_11),
            .ltout(),
            .carryin(n13976),
            .carryout(n13977),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32375),
            .sr(N__30703));
    defparam acadc_skipcnt_i0_i12_LC_13_18_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i12_LC_13_18_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i12_LC_13_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i12_LC_13_18_3 (
            .in0(_gnd_net_),
            .in1(N__30028),
            .in2(_gnd_net_),
            .in3(N__28865),
            .lcout(acadc_skipcnt_12),
            .ltout(),
            .carryin(n13977),
            .carryout(n13978),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32375),
            .sr(N__30703));
    defparam acadc_skipcnt_i0_i13_LC_13_18_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i13_LC_13_18_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i13_LC_13_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i13_LC_13_18_4 (
            .in0(_gnd_net_),
            .in1(N__32230),
            .in2(_gnd_net_),
            .in3(N__28862),
            .lcout(acadc_skipcnt_13),
            .ltout(),
            .carryin(n13978),
            .carryout(n13979),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32375),
            .sr(N__30703));
    defparam acadc_skipcnt_i0_i14_LC_13_18_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i14_LC_13_18_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i14_LC_13_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i14_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(N__30139),
            .in2(_gnd_net_),
            .in3(N__28859),
            .lcout(acadc_skipcnt_14),
            .ltout(),
            .carryin(n13979),
            .carryout(n13980),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32375),
            .sr(N__30703));
    defparam acadc_skipcnt_i0_i15_LC_13_18_6.C_ON=1'b0;
    defparam acadc_skipcnt_i0_i15_LC_13_18_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i15_LC_13_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i15_LC_13_18_6 (
            .in0(_gnd_net_),
            .in1(N__31486),
            .in2(_gnd_net_),
            .in3(N__28856),
            .lcout(acadc_skipcnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__32375),
            .sr(N__30703));
    defparam mux_1469_i7_4_lut_LC_14_2_4.C_ON=1'b0;
    defparam mux_1469_i7_4_lut_LC_14_2_4.SEQ_MODE=4'b0000;
    defparam mux_1469_i7_4_lut_LC_14_2_4.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1469_i7_4_lut_LC_14_2_4 (
            .in0(N__29087),
            .in1(N__48084),
            .in2(N__29074),
            .in3(N__47084),
            .lcout(n4102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13097_4_lut_3_lut_LC_14_3_4 .C_ON=1'b0;
    defparam \comm_spi.i13097_4_lut_3_lut_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13097_4_lut_3_lut_LC_14_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i13097_4_lut_3_lut_LC_14_3_4  (
            .in0(N__29028),
            .in1(N__30971),
            .in2(_gnd_net_),
            .in3(N__46599),
            .lcout(\comm_spi.n16902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i5_7364_7365_reset_LC_14_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_7364_7365_reset_LC_14_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i5_7364_7365_reset_LC_14_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_7364_7365_reset_LC_14_4_0  (
            .in0(N__46397),
            .in1(N__28945),
            .in2(_gnd_net_),
            .in3(N__28963),
            .lcout(\comm_spi.n10476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42404),
            .ce(),
            .sr(N__32537));
    defparam \comm_spi.data_tx_i6_7368_7369_reset_LC_14_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_7368_7369_reset_LC_14_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i6_7368_7369_reset_LC_14_5_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_tx_i6_7368_7369_reset_LC_14_5_0  (
            .in0(N__28927),
            .in1(N__28897),
            .in2(_gnd_net_),
            .in3(N__29005),
            .lcout(\comm_spi.n10480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42439),
            .ce(),
            .sr(N__28973));
    defparam \comm_spi.data_tx_i5_7364_7365_set_LC_14_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_7364_7365_set_LC_14_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i5_7364_7365_set_LC_14_6_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.data_tx_i5_7364_7365_set_LC_14_6_0  (
            .in0(N__28967),
            .in1(N__46396),
            .in2(_gnd_net_),
            .in3(N__28949),
            .lcout(\comm_spi.n10475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42431),
            .ce(),
            .sr(N__28916));
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_14_6_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_14_6_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \comm_spi.RESET_I_0_94_2_lut_LC_14_6_2  (
            .in0(N__32562),
            .in1(N__46582),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13107_4_lut_3_lut_LC_14_6_3 .C_ON=1'b0;
    defparam \comm_spi.i13107_4_lut_3_lut_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13107_4_lut_3_lut_LC_14_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i13107_4_lut_3_lut_LC_14_6_3  (
            .in0(N__46583),
            .in1(N__32563),
            .in2(_gnd_net_),
            .in3(N__28896),
            .lcout(\comm_spi.n16896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_14_6_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_14_6_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \comm_spi.RESET_I_0_91_2_lut_LC_14_6_4  (
            .in0(N__51404),
            .in1(N__46581),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.iclk_N_802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12653_2_lut_LC_14_6_5.C_ON=1'b0;
    defparam i12653_2_lut_LC_14_6_5.SEQ_MODE=4'b0000;
    defparam i12653_2_lut_LC_14_6_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12653_2_lut_LC_14_6_5 (
            .in0(N__47985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32038),
            .lcout(n15474),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12656_2_lut_LC_14_6_6.C_ON=1'b0;
    defparam i12656_2_lut_LC_14_6_6.SEQ_MODE=4'b0000;
    defparam i12656_2_lut_LC_14_6_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12656_2_lut_LC_14_6_6 (
            .in0(_gnd_net_),
            .in1(N__47983),
            .in2(_gnd_net_),
            .in3(N__29239),
            .lcout(n15478),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12659_2_lut_LC_14_6_7.C_ON=1'b0;
    defparam i12659_2_lut_LC_14_6_7.SEQ_MODE=4'b0000;
    defparam i12659_2_lut_LC_14_6_7.LUT_INIT=16'b0100010001000100;
    LogicCell40 i12659_2_lut_LC_14_6_7 (
            .in0(N__47984),
            .in1(N__31382),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n15680),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_valid_85_LC_14_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_valid_85_LC_14_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_valid_85_LC_14_7_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.data_valid_85_LC_14_7_0  (
            .in0(N__38384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38423),
            .lcout(comm_data_vld),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.data_valid_85C_net ),
            .ce(),
            .sr(N__46580));
    defparam \comm_spi.imiso_83_7340_7341_set_LC_14_8_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_7340_7341_set_LC_14_8_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imiso_83_7340_7341_set_LC_14_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.imiso_83_7340_7341_set_LC_14_8_0  (
            .in0(N__30843),
            .in1(N__29152),
            .in2(_gnd_net_),
            .in3(N__29135),
            .lcout(\comm_spi.n10451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_7340_7341_setC_net ),
            .ce(),
            .sr(N__30768));
    defparam i12177_3_lut_LC_14_8_1.C_ON=1'b0;
    defparam i12177_3_lut_LC_14_8_1.SEQ_MODE=4'b0000;
    defparam i12177_3_lut_LC_14_8_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12177_3_lut_LC_14_8_1 (
            .in0(N__38765),
            .in1(N__39995),
            .in2(_gnd_net_),
            .in3(N__34396),
            .lcout(n15387),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12180_3_lut_LC_14_8_2.C_ON=1'b0;
    defparam i12180_3_lut_LC_14_8_2.SEQ_MODE=4'b0000;
    defparam i12180_3_lut_LC_14_8_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12180_3_lut_LC_14_8_2 (
            .in0(N__36712),
            .in1(N__34119),
            .in2(_gnd_net_),
            .in3(N__38764),
            .lcout(n15390),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9624_2_lut_3_lut_LC_14_8_3.C_ON=1'b0;
    defparam i9624_2_lut_3_lut_LC_14_8_3.SEQ_MODE=4'b0000;
    defparam i9624_2_lut_3_lut_LC_14_8_3.LUT_INIT=16'b0000000000100010;
    LogicCell40 i9624_2_lut_3_lut_LC_14_8_3 (
            .in0(N__34120),
            .in1(N__49875),
            .in2(_gnd_net_),
            .in3(N__49543),
            .lcout(n14_adj_1211),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9632_2_lut_3_lut_LC_14_8_5.C_ON=1'b0;
    defparam i9632_2_lut_3_lut_LC_14_8_5.SEQ_MODE=4'b0000;
    defparam i9632_2_lut_3_lut_LC_14_8_5.LUT_INIT=16'b0000000000100010;
    LogicCell40 i9632_2_lut_3_lut_LC_14_8_5 (
            .in0(N__38924),
            .in1(N__49879),
            .in2(_gnd_net_),
            .in3(N__49545),
            .lcout(n14_adj_1205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9637_2_lut_3_lut_LC_14_8_6.C_ON=1'b0;
    defparam i9637_2_lut_3_lut_LC_14_8_6.SEQ_MODE=4'b0000;
    defparam i9637_2_lut_3_lut_LC_14_8_6.LUT_INIT=16'b0000010100000000;
    LogicCell40 i9637_2_lut_3_lut_LC_14_8_6 (
            .in0(N__49544),
            .in1(_gnd_net_),
            .in2(N__50111),
            .in3(N__41096),
            .lcout(n14_adj_1198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i10_LC_14_9_0 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i10_LC_14_9_0 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i10_LC_14_9_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i10_LC_14_9_0  (
            .in0(N__35747),
            .in1(N__48525),
            .in2(N__29213),
            .in3(N__34352),
            .lcout(\CLOCK_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i11_LC_14_9_1 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i11_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i11_LC_14_9_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i11_LC_14_9_1  (
            .in0(N__48526),
            .in1(N__35748),
            .in2(N__29285),
            .in3(N__41257),
            .lcout(\CLOCK_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i12_LC_14_9_2 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i12_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i12_LC_14_9_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \CLOCK_DDS.tmp_buf_i12_LC_14_9_2  (
            .in0(N__32039),
            .in1(N__29276),
            .in2(N__35763),
            .in3(N__48527),
            .lcout(\CLOCK_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i13_LC_14_9_3 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i13_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i13_LC_14_9_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i13_LC_14_9_3  (
            .in0(N__48528),
            .in1(N__35752),
            .in2(N__29270),
            .in3(N__34067),
            .lcout(\CLOCK_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i14_LC_14_9_4 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i14_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i14_LC_14_9_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i14_LC_14_9_4  (
            .in0(N__35753),
            .in1(N__48529),
            .in2(N__29258),
            .in3(N__29546),
            .lcout(\CLOCK_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i15_LC_14_9_5 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i15_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i15_LC_14_9_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \CLOCK_DDS.tmp_buf_i15_LC_14_9_5  (
            .in0(N__31456),
            .in1(N__29249),
            .in2(N__48546),
            .in3(N__35754),
            .lcout(tmp_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i9_LC_14_9_6 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i9_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i9_LC_14_9_6 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \CLOCK_DDS.tmp_buf_i9_LC_14_9_6  (
            .in0(N__29243),
            .in1(N__29204),
            .in2(N__35764),
            .in3(N__48536),
            .lcout(\CLOCK_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i8_LC_14_9_7 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i8_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i8_LC_14_9_7 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \CLOCK_DDS.tmp_buf_i8_LC_14_9_7  (
            .in0(N__33849),
            .in1(N__31217),
            .in2(N__48547),
            .in3(N__35755),
            .lcout(\CLOCK_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51143),
            .ce(N__31210),
            .sr(_gnd_net_));
    defparam mux_1513_i5_4_lut_LC_14_10_0.C_ON=1'b0;
    defparam mux_1513_i5_4_lut_LC_14_10_0.SEQ_MODE=4'b0000;
    defparam mux_1513_i5_4_lut_LC_14_10_0.LUT_INIT=16'b1101110000010000;
    LogicCell40 mux_1513_i5_4_lut_LC_14_10_0 (
            .in0(N__45293),
            .in1(N__47308),
            .in2(N__29372),
            .in3(N__41600),
            .lcout(),
            .ltout(n4260_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i4_LC_14_10_1.C_ON=1'b0;
    defparam comm_buf_1__i4_LC_14_10_1.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i4_LC_14_10_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i4_LC_14_10_1 (
            .in0(N__39904),
            .in1(_gnd_net_),
            .in2(N__29342),
            .in3(N__50131),
            .lcout(comm_buf_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51154),
            .ce(N__44698),
            .sr(N__44645));
    defparam i9633_2_lut_3_lut_LC_14_10_2.C_ON=1'b0;
    defparam i9633_2_lut_3_lut_LC_14_10_2.SEQ_MODE=4'b0000;
    defparam i9633_2_lut_3_lut_LC_14_10_2.LUT_INIT=16'b0000010000000100;
    LogicCell40 i9633_2_lut_3_lut_LC_14_10_2 (
            .in0(N__49542),
            .in1(N__31598),
            .in2(N__50290),
            .in3(_gnd_net_),
            .lcout(n14_adj_1196),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9630_2_lut_3_lut_LC_14_10_5.C_ON=1'b0;
    defparam i9630_2_lut_3_lut_LC_14_10_5.SEQ_MODE=4'b0000;
    defparam i9630_2_lut_3_lut_LC_14_10_5.LUT_INIT=16'b0000000000100010;
    LogicCell40 i9630_2_lut_3_lut_LC_14_10_5 (
            .in0(N__36967),
            .in1(N__50127),
            .in2(_gnd_net_),
            .in3(N__49541),
            .lcout(n14_adj_1207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12192_3_lut_LC_14_10_6.C_ON=1'b0;
    defparam i12192_3_lut_LC_14_10_6.SEQ_MODE=4'b0000;
    defparam i12192_3_lut_LC_14_10_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12192_3_lut_LC_14_10_6 (
            .in0(N__38779),
            .in1(N__31597),
            .in2(_gnd_net_),
            .in3(N__36968),
            .lcout(n15402),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i11_LC_14_11_0.C_ON=1'b0;
    defparam acadc_skipCount_i11_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i11_LC_14_11_0.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i11_LC_14_11_0 (
            .in0(N__30106),
            .in1(N__51679),
            .in2(N__43561),
            .in3(N__41827),
            .lcout(acadc_skipCount_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51167),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_28_LC_14_11_1.C_ON=1'b0;
    defparam i1_4_lut_adj_28_LC_14_11_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_28_LC_14_11_1.LUT_INIT=16'b1100000011000100;
    LogicCell40 i1_4_lut_adj_28_LC_14_11_1 (
            .in0(N__34010),
            .in1(N__52349),
            .in2(N__51769),
            .in3(N__50609),
            .lcout(n9224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i8_LC_14_11_2.C_ON=1'b0;
    defparam req_data_cnt_i8_LC_14_11_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i8_LC_14_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i8_LC_14_11_2 (
            .in0(N__40464),
            .in1(N__37273),
            .in2(_gnd_net_),
            .in3(N__31409),
            .lcout(req_data_cnt_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51167),
            .ce(),
            .sr(_gnd_net_));
    defparam i130_3_lut_adj_98_LC_14_11_3.C_ON=1'b0;
    defparam i130_3_lut_adj_98_LC_14_11_3.SEQ_MODE=4'b0000;
    defparam i130_3_lut_adj_98_LC_14_11_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 i130_3_lut_adj_98_LC_14_11_3 (
            .in0(N__29327),
            .in1(N__45216),
            .in2(_gnd_net_),
            .in3(N__30105),
            .lcout(),
            .ltout(n90_adj_1154_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i125_4_lut_adj_99_LC_14_11_4.C_ON=1'b0;
    defparam i125_4_lut_adj_99_LC_14_11_4.SEQ_MODE=4'b0000;
    defparam i125_4_lut_adj_99_LC_14_11_4.LUT_INIT=16'b1110001011000000;
    LogicCell40 i125_4_lut_adj_99_LC_14_11_4 (
            .in0(N__45217),
            .in1(N__47864),
            .in2(N__29303),
            .in3(N__37427),
            .lcout(n72),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12629_2_lut_LC_14_11_5.C_ON=1'b0;
    defparam i12629_2_lut_LC_14_11_5.SEQ_MODE=4'b0000;
    defparam i12629_2_lut_LC_14_11_5.LUT_INIT=16'b0100010001000100;
    LogicCell40 i12629_2_lut_LC_14_11_5 (
            .in0(N__47865),
            .in1(N__29428),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n15479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i30_LC_14_11_6 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i30_LC_14_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i30_LC_14_11_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i30_LC_14_11_6  (
            .in0(N__36878),
            .in1(N__49205),
            .in2(N__43738),
            .in3(N__48818),
            .lcout(cmd_rdadctmp_30_adj_1082),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51167),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i31_LC_14_11_7 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i31_LC_14_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i31_LC_14_11_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i31_LC_14_11_7  (
            .in0(N__48817),
            .in1(N__29386),
            .in2(N__49241),
            .in3(N__43734),
            .lcout(cmd_rdadctmp_31_adj_1081),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51167),
            .ce(),
            .sr(_gnd_net_));
    defparam i3157_3_lut_LC_14_12_0.C_ON=1'b0;
    defparam i3157_3_lut_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam i3157_3_lut_LC_14_12_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 i3157_3_lut_LC_14_12_0 (
            .in0(N__38977),
            .in1(N__30258),
            .in2(_gnd_net_),
            .in3(N__40505),
            .lcout(n8_adj_1221),
            .ltout(n8_adj_1221_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i7_LC_14_12_1.C_ON=1'b0;
    defparam data_index_i7_LC_14_12_1.SEQ_MODE=4'b1000;
    defparam data_index_i7_LC_14_12_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 data_index_i7_LC_14_12_1 (
            .in0(N__51636),
            .in1(N__52350),
            .in2(N__29375),
            .in3(N__30542),
            .lcout(data_index_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51185),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_90_LC_14_12_2.C_ON=1'b0;
    defparam i6_4_lut_adj_90_LC_14_12_2.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_90_LC_14_12_2.LUT_INIT=16'b0111101111011110;
    LogicCell40 i6_4_lut_adj_90_LC_14_12_2 (
            .in0(N__34925),
            .in1(N__40324),
            .in2(N__31337),
            .in3(N__34688),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i5_3_lut_LC_14_12_4.C_ON=1'b0;
    defparam mux_1498_i5_3_lut_LC_14_12_4.SEQ_MODE=4'b0000;
    defparam mux_1498_i5_3_lut_LC_14_12_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_1498_i5_3_lut_LC_14_12_4 (
            .in0(N__31576),
            .in1(N__40784),
            .in2(_gnd_net_),
            .in3(N__47822),
            .lcout(n4205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i9_LC_14_12_5.C_ON=1'b0;
    defparam req_data_cnt_i9_LC_14_12_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i9_LC_14_12_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i9_LC_14_12_5 (
            .in0(N__37238),
            .in1(N__40455),
            .in2(_gnd_net_),
            .in3(N__29488),
            .lcout(req_data_cnt_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51185),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i8_LC_14_12_7.C_ON=1'b0;
    defparam buf_device_acadc_i8_LC_14_12_7.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i8_LC_14_12_7.LUT_INIT=16'b0000101011001100;
    LogicCell40 buf_device_acadc_i8_LC_14_12_7 (
            .in0(N__38925),
            .in1(N__29356),
            .in2(N__51738),
            .in3(N__31849),
            .lcout(buf_device_acadc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51185),
            .ce(),
            .sr(_gnd_net_));
    defparam i9631_2_lut_3_lut_LC_14_13_0.C_ON=1'b0;
    defparam i9631_2_lut_3_lut_LC_14_13_0.SEQ_MODE=4'b0000;
    defparam i9631_2_lut_3_lut_LC_14_13_0.LUT_INIT=16'b0000000001000100;
    LogicCell40 i9631_2_lut_3_lut_LC_14_13_0 (
            .in0(N__49540),
            .in1(N__41886),
            .in2(_gnd_net_),
            .in3(N__50288),
            .lcout(n14_adj_1206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i14_LC_14_13_1.C_ON=1'b0;
    defparam buf_dds_i14_LC_14_13_1.SEQ_MODE=4'b1000;
    defparam buf_dds_i14_LC_14_13_1.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i14_LC_14_13_1 (
            .in0(N__41887),
            .in1(N__29544),
            .in2(N__41518),
            .in3(N__41369),
            .lcout(buf_dds_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51203),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i3_3_lut_LC_14_13_2.C_ON=1'b0;
    defparam mux_1511_i3_3_lut_LC_14_13_2.SEQ_MODE=4'b0000;
    defparam mux_1511_i3_3_lut_LC_14_13_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_1511_i3_3_lut_LC_14_13_2 (
            .in0(N__29522),
            .in1(N__45652),
            .in2(_gnd_net_),
            .in3(N__31517),
            .lcout(n4252),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_75_LC_14_13_4.C_ON=1'b0;
    defparam i8_4_lut_adj_75_LC_14_13_4.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_75_LC_14_13_4.LUT_INIT=16'b0111110110111110;
    LogicCell40 i8_4_lut_adj_75_LC_14_13_4 (
            .in0(N__34855),
            .in1(N__29512),
            .in2(N__35402),
            .in3(N__29484),
            .lcout(),
            .ltout(n24_adj_1216_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_113_LC_14_13_5.C_ON=1'b0;
    defparam i14_4_lut_adj_113_LC_14_13_5.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_113_LC_14_13_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_113_LC_14_13_5 (
            .in0(N__29468),
            .in1(N__31895),
            .in2(N__29462),
            .in3(N__31631),
            .lcout(n30_adj_1278),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3754_2_lut_LC_14_13_6.C_ON=1'b0;
    defparam i3754_2_lut_LC_14_13_6.SEQ_MODE=4'b0000;
    defparam i3754_2_lut_LC_14_13_6.LUT_INIT=16'b1111111110101010;
    LogicCell40 i3754_2_lut_LC_14_13_6 (
            .in0(N__49539),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50287),
            .lcout(n6791),
            .ltout(n6791_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i0_LC_14_13_7.C_ON=1'b0;
    defparam acadc_skipCount_i0_LC_14_13_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i0_LC_14_13_7.LUT_INIT=16'b0011101100001000;
    LogicCell40 acadc_skipCount_i0_LC_14_13_7 (
            .in0(N__36715),
            .in1(N__41785),
            .in2(N__29453),
            .in3(N__34318),
            .lcout(acadc_skipCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51203),
            .ce(),
            .sr(_gnd_net_));
    defparam i2358_3_lut_LC_14_14_0.C_ON=1'b0;
    defparam i2358_3_lut_LC_14_14_0.SEQ_MODE=4'b0000;
    defparam i2358_3_lut_LC_14_14_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i2358_3_lut_LC_14_14_0 (
            .in0(N__30004),
            .in1(N__36714),
            .in2(_gnd_net_),
            .in3(N__40532),
            .lcout(n8_adj_1178),
            .ltout(n8_adj_1178_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i0_LC_14_14_1.C_ON=1'b0;
    defparam data_index_i0_LC_14_14_1.SEQ_MODE=4'b1000;
    defparam data_index_i0_LC_14_14_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 data_index_i0_LC_14_14_1 (
            .in0(N__51664),
            .in1(N__52426),
            .in2(N__29450),
            .in3(N__29447),
            .lcout(data_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51220),
            .ce(),
            .sr(_gnd_net_));
    defparam i2356_3_lut_LC_14_14_2.C_ON=1'b0;
    defparam i2356_3_lut_LC_14_14_2.SEQ_MODE=4'b0000;
    defparam i2356_3_lut_LC_14_14_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 i2356_3_lut_LC_14_14_2 (
            .in0(N__30003),
            .in1(N__31673),
            .in2(_gnd_net_),
            .in3(N__29987),
            .lcout(n7_adj_1177),
            .ltout(n7_adj_1177_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_0_i15_4_lut_LC_14_14_3.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_0_i15_4_lut_LC_14_14_3.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_0_i15_4_lut_LC_14_14_3.LUT_INIT=16'b0111010000110000;
    LogicCell40 comm_state_3__I_0_394_Mux_0_i15_4_lut_LC_14_14_3 (
            .in0(N__51663),
            .in1(N__52425),
            .in2(N__29873),
            .in3(N__29870),
            .lcout(data_index_9_N_258_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3201_3_lut_LC_14_14_4.C_ON=1'b0;
    defparam i3201_3_lut_LC_14_14_4.SEQ_MODE=4'b0000;
    defparam i3201_3_lut_LC_14_14_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i3201_3_lut_LC_14_14_4 (
            .in0(N__39997),
            .in1(N__29946),
            .in2(_gnd_net_),
            .in3(N__40533),
            .lcout(n8_adj_1231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_70_LC_14_14_5.C_ON=1'b0;
    defparam i1_4_lut_adj_70_LC_14_14_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_70_LC_14_14_5.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_70_LC_14_14_5 (
            .in0(N__29759),
            .in1(N__34760),
            .in2(N__29741),
            .in3(N__34314),
            .lcout(),
            .ltout(n17_adj_1277_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_LC_14_14_6.C_ON=1'b0;
    defparam i15_4_lut_LC_14_14_6.SEQ_MODE=4'b0000;
    defparam i15_4_lut_LC_14_14_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_LC_14_14_6 (
            .in0(N__29723),
            .in1(N__32246),
            .in2(N__29714),
            .in3(N__30086),
            .lcout(n31),
            .ltout(n31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_304_LC_14_14_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_304_LC_14_14_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_304_LC_14_14_7.LUT_INIT=16'b1010000000000000;
    LogicCell40 i1_2_lut_3_lut_adj_304_LC_14_14_7 (
            .in0(N__38093),
            .in1(_gnd_net_),
            .in2(N__29702),
            .in3(N__41045),
            .lcout(n15187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i2_LC_14_15_0.C_ON=1'b0;
    defparam data_index_i2_LC_14_15_0.SEQ_MODE=4'b1000;
    defparam data_index_i2_LC_14_15_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i2_LC_14_15_0 (
            .in0(N__52433),
            .in1(N__29693),
            .in2(N__51844),
            .in3(N__29927),
            .lcout(data_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51237),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_2_i15_4_lut_LC_14_15_2.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_2_i15_4_lut_LC_14_15_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_2_i15_4_lut_LC_14_15_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_394_Mux_2_i15_4_lut_LC_14_15_2 (
            .in0(N__52432),
            .in1(N__29692),
            .in2(N__51842),
            .in3(N__29926),
            .lcout(data_index_9_N_258_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i12_LC_14_15_3.C_ON=1'b0;
    defparam acadc_skipCount_i12_LC_14_15_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i12_LC_14_15_3.LUT_INIT=16'b0011000010111000;
    LogicCell40 acadc_skipCount_i12_LC_14_15_3 (
            .in0(N__36990),
            .in1(N__41824),
            .in2(N__30058),
            .in3(N__51749),
            .lcout(acadc_skipCount_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51237),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i4_LC_14_15_4.C_ON=1'b0;
    defparam buf_device_acadc_i4_LC_14_15_4.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i4_LC_14_15_4.LUT_INIT=16'b0000110010101010;
    LogicCell40 buf_device_acadc_i4_LC_14_15_4 (
            .in0(N__29565),
            .in1(N__43558),
            .in2(N__51843),
            .in3(N__31871),
            .lcout(M_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51237),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_14_15_5.C_ON=1'b0;
    defparam i7_4_lut_LC_14_15_5.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_14_15_5.LUT_INIT=16'b0110111111110110;
    LogicCell40 i7_4_lut_LC_14_15_5 (
            .in0(N__41704),
            .in1(N__30143),
            .in2(N__30125),
            .in3(N__30107),
            .lcout(),
            .ltout(n23_adj_1199_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_14_15_6.C_ON=1'b0;
    defparam i14_4_lut_LC_14_15_6.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_14_15_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_LC_14_15_6 (
            .in0(N__31472),
            .in1(N__31919),
            .in2(N__30089),
            .in3(N__30014),
            .lcout(n30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_14_15_7.C_ON=1'b0;
    defparam i5_4_lut_LC_14_15_7.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_14_15_7.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_LC_14_15_7 (
            .in0(N__30080),
            .in1(N__30048),
            .in2(N__30032),
            .in3(N__34206),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_2_lut_LC_14_16_0.C_ON=1'b1;
    defparam add_1443_2_lut_LC_14_16_0.SEQ_MODE=4'b0000;
    defparam add_1443_2_lut_LC_14_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_1443_2_lut_LC_14_16_0 (
            .in0(_gnd_net_),
            .in1(N__43616),
            .in2(N__30008),
            .in3(_gnd_net_),
            .lcout(data_index_9_N_647_0),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(n14031),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_3_lut_LC_14_16_1.C_ON=1'b1;
    defparam add_1443_3_lut_LC_14_16_1.SEQ_MODE=4'b0000;
    defparam add_1443_3_lut_LC_14_16_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_3_lut_LC_14_16_1 (
            .in0(N__29977),
            .in1(N__29976),
            .in2(N__31699),
            .in3(N__29951),
            .lcout(n7_adj_1232),
            .ltout(),
            .carryin(n14031),
            .carryout(n14032),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_4_lut_LC_14_16_2.C_ON=1'b1;
    defparam add_1443_4_lut_LC_14_16_2.SEQ_MODE=4'b0000;
    defparam add_1443_4_lut_LC_14_16_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_4_lut_LC_14_16_2 (
            .in0(N__29948),
            .in1(N__29947),
            .in2(N__31703),
            .in3(N__29918),
            .lcout(n7_adj_1230),
            .ltout(),
            .carryin(n14032),
            .carryout(n14033),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_5_lut_LC_14_16_3.C_ON=1'b1;
    defparam add_1443_5_lut_LC_14_16_3.SEQ_MODE=4'b0000;
    defparam add_1443_5_lut_LC_14_16_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_5_lut_LC_14_16_3 (
            .in0(N__30232),
            .in1(N__30231),
            .in2(N__31700),
            .in3(N__29915),
            .lcout(n7_adj_1228),
            .ltout(),
            .carryin(n14033),
            .carryout(n14034),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_6_lut_LC_14_16_4.C_ON=1'b1;
    defparam add_1443_6_lut_LC_14_16_4.SEQ_MODE=4'b0000;
    defparam add_1443_6_lut_LC_14_16_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_6_lut_LC_14_16_4 (
            .in0(N__29912),
            .in1(N__29911),
            .in2(N__31704),
            .in3(N__29876),
            .lcout(n7_adj_1226),
            .ltout(),
            .carryin(n14034),
            .carryout(n14035),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_7_lut_LC_14_16_5.C_ON=1'b1;
    defparam add_1443_7_lut_LC_14_16_5.SEQ_MODE=4'b0000;
    defparam add_1443_7_lut_LC_14_16_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_7_lut_LC_14_16_5 (
            .in0(N__32056),
            .in1(N__32055),
            .in2(N__31701),
            .in3(N__30266),
            .lcout(n7_adj_1224),
            .ltout(),
            .carryin(n14035),
            .carryout(n14036),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_8_lut_LC_14_16_6.C_ON=1'b1;
    defparam add_1443_8_lut_LC_14_16_6.SEQ_MODE=4'b0000;
    defparam add_1443_8_lut_LC_14_16_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_8_lut_LC_14_16_6 (
            .in0(N__30577),
            .in1(N__30576),
            .in2(N__31705),
            .in3(N__30263),
            .lcout(n7_adj_1222),
            .ltout(),
            .carryin(n14036),
            .carryout(n14037),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_9_lut_LC_14_16_7.C_ON=1'b1;
    defparam add_1443_9_lut_LC_14_16_7.SEQ_MODE=4'b0000;
    defparam add_1443_9_lut_LC_14_16_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_9_lut_LC_14_16_7 (
            .in0(N__30260),
            .in1(N__30259),
            .in2(N__31702),
            .in3(N__30239),
            .lcout(n7_adj_1220),
            .ltout(),
            .carryin(n14037),
            .carryout(n14038),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1443_10_lut_LC_14_17_0.C_ON=1'b0;
    defparam add_1443_10_lut_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam add_1443_10_lut_LC_14_17_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_1443_10_lut_LC_14_17_0 (
            .in0(N__32657),
            .in1(N__32656),
            .in2(N__31712),
            .in3(N__30236),
            .lcout(n7_adj_1218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i19_LC_14_17_2 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i19_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i19_LC_14_17_2 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i19_LC_14_17_2  (
            .in0(N__38284),
            .in1(N__46089),
            .in2(N__46164),
            .in3(N__53474),
            .lcout(cmd_rdadctmp_19_adj_1057),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51269),
            .ce(),
            .sr(_gnd_net_));
    defparam i3145_3_lut_LC_14_17_3.C_ON=1'b0;
    defparam i3145_3_lut_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam i3145_3_lut_LC_14_17_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i3145_3_lut_LC_14_17_3 (
            .in0(N__32655),
            .in1(N__34124),
            .in2(_gnd_net_),
            .in3(N__40545),
            .lcout(n8_adj_1219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3193_3_lut_LC_14_17_4.C_ON=1'b0;
    defparam i3193_3_lut_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam i3193_3_lut_LC_14_17_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 i3193_3_lut_LC_14_17_4 (
            .in0(N__40546),
            .in1(N__44776),
            .in2(_gnd_net_),
            .in3(N__30233),
            .lcout(n8_adj_1229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i3_LC_14_17_6.C_ON=1'b0;
    defparam data_index_i3_LC_14_17_6.SEQ_MODE=4'b1000;
    defparam data_index_i3_LC_14_17_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i3_LC_14_17_6 (
            .in0(N__52442),
            .in1(N__32501),
            .in2(N__51918),
            .in3(N__32489),
            .lcout(data_index_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51269),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.i18_3_lut_LC_14_17_7 .C_ON=1'b0;
    defparam \ADC_VAC2.i18_3_lut_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i18_3_lut_LC_14_17_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ADC_VAC2.i18_3_lut_LC_14_17_7  (
            .in0(N__30212),
            .in1(N__36475),
            .in2(_gnd_net_),
            .in3(N__30604),
            .lcout(\ADC_VAC2.n15280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13029_2_lut_LC_14_18_1.C_ON=1'b0;
    defparam i13029_2_lut_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam i13029_2_lut_LC_14_18_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 i13029_2_lut_LC_14_18_1 (
            .in0(N__32835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32345),
            .lcout(n10532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13050_2_lut_3_lut_LC_14_18_4.C_ON=1'b0;
    defparam i13050_2_lut_3_lut_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam i13050_2_lut_3_lut_LC_14_18_4.LUT_INIT=16'b0000000000010001;
    LogicCell40 i13050_2_lut_3_lut_LC_14_18_4 (
            .in0(N__32729),
            .in1(N__32836),
            .in2(_gnd_net_),
            .in3(N__38122),
            .lcout(n15344),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i17_3_lut_LC_14_18_5.C_ON=1'b0;
    defparam i17_3_lut_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam i17_3_lut_LC_14_18_5.LUT_INIT=16'b1101100011011000;
    LogicCell40 i17_3_lut_LC_14_18_5 (
            .in0(N__38123),
            .in1(N__32925),
            .in2(N__32840),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n15328_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_trig_329_LC_14_18_6.C_ON=1'b0;
    defparam acadc_trig_329_LC_14_18_6.SEQ_MODE=4'b1000;
    defparam acadc_trig_329_LC_14_18_6.LUT_INIT=16'b1111111000000100;
    LogicCell40 acadc_trig_329_LC_14_18_6 (
            .in0(N__32728),
            .in1(N__30674),
            .in2(N__30662),
            .in3(N__30618),
            .lcout(acadc_trig),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_trig_329C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i3165_3_lut_LC_14_18_7.C_ON=1'b0;
    defparam i3165_3_lut_LC_14_18_7.SEQ_MODE=4'b0000;
    defparam i3165_3_lut_LC_14_18_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 i3165_3_lut_LC_14_18_7 (
            .in0(N__33969),
            .in1(N__30578),
            .in2(_gnd_net_),
            .in3(N__40547),
            .lcout(n8_adj_1223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_7_i15_4_lut_LC_14_19_1.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_7_i15_4_lut_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_7_i15_4_lut_LC_14_19_1.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_394_Mux_7_i15_4_lut_LC_14_19_1 (
            .in0(N__52467),
            .in1(N__30551),
            .in2(N__51909),
            .in3(N__30541),
            .lcout(data_index_9_N_258_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_6_i15_4_lut_LC_14_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_6_i15_4_lut_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_6_i15_4_lut_LC_14_19_4.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_state_3__I_0_394_Mux_6_i15_4_lut_LC_14_19_4 (
            .in0(N__52468),
            .in1(N__30424),
            .in2(N__30397),
            .in3(N__51851),
            .lcout(data_index_9_N_258_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i7336_3_lut_LC_15_4_6 .C_ON=1'b0;
    defparam \comm_spi.i7336_3_lut_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i7336_3_lut_LC_15_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i7336_3_lut_LC_15_4_6  (
            .in0(N__30788),
            .in1(N__30272),
            .in2(_gnd_net_),
            .in3(N__30844),
            .lcout(ICE_SPI_MISO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.MISO_48_7334_7335_reset_LC_15_5_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_7334_7335_reset_LC_15_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.MISO_48_7334_7335_reset_LC_15_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.MISO_48_7334_7335_reset_LC_15_5_0  (
            .in0(N__30890),
            .in1(N__30863),
            .in2(_gnd_net_),
            .in3(N__30834),
            .lcout(\comm_spi.n10446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_7334_7335_resetC_net ),
            .ce(),
            .sr(N__31000));
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_15_6_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_15_6_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_104_2_lut_LC_15_6_1  (
            .in0(N__46556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30967),
            .lcout(\comm_spi.data_tx_7__N_825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i105_4_lut_adj_131_LC_15_6_4.C_ON=1'b0;
    defparam i105_4_lut_adj_131_LC_15_6_4.SEQ_MODE=4'b0000;
    defparam i105_4_lut_adj_131_LC_15_6_4.LUT_INIT=16'b0101000010001000;
    LogicCell40 i105_4_lut_adj_131_LC_15_6_4 (
            .in0(N__45285),
            .in1(N__30917),
            .in2(N__37610),
            .in3(N__47855),
            .lcout(n66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.MISO_48_7334_7335_set_LC_15_7_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_7334_7335_set_LC_15_7_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.MISO_48_7334_7335_set_LC_15_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.MISO_48_7334_7335_set_LC_15_7_0  (
            .in0(N__30886),
            .in1(N__30856),
            .in2(_gnd_net_),
            .in3(N__30842),
            .lcout(\comm_spi.n10445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_7334_7335_setC_net ),
            .ce(),
            .sr(N__30778));
    defparam i1_2_lut_3_lut_adj_176_LC_15_7_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_176_LC_15_7_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_176_LC_15_7_2.LUT_INIT=16'b1011101111111111;
    LogicCell40 i1_2_lut_3_lut_adj_176_LC_15_7_2 (
            .in0(N__52238),
            .in1(N__49996),
            .in2(_gnd_net_),
            .in3(N__49504),
            .lcout(n15204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_181_LC_15_7_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_181_LC_15_7_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_181_LC_15_7_3.LUT_INIT=16'b1111101000000000;
    LogicCell40 i1_2_lut_3_lut_adj_181_LC_15_7_3 (
            .in0(N__49505),
            .in1(_gnd_net_),
            .in2(N__50219),
            .in3(N__52239),
            .lcout(n10640),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_216_LC_15_7_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_216_LC_15_7_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_216_LC_15_7_4.LUT_INIT=16'b0000000000100010;
    LogicCell40 i1_2_lut_3_lut_adj_216_LC_15_7_4 (
            .in0(N__52240),
            .in1(N__50000),
            .in2(_gnd_net_),
            .in3(N__49507),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9642_2_lut_3_lut_LC_15_7_6.C_ON=1'b0;
    defparam i9642_2_lut_3_lut_LC_15_7_6.SEQ_MODE=4'b0000;
    defparam i9642_2_lut_3_lut_LC_15_7_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i9642_2_lut_3_lut_LC_15_7_6 (
            .in0(N__37883),
            .in1(N__50004),
            .in2(_gnd_net_),
            .in3(N__49508),
            .lcout(n14_adj_1213),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9697_2_lut_3_lut_LC_15_7_7.C_ON=1'b0;
    defparam i9697_2_lut_3_lut_LC_15_7_7.SEQ_MODE=4'b0000;
    defparam i9697_2_lut_3_lut_LC_15_7_7.LUT_INIT=16'b0000010100000000;
    LogicCell40 i9697_2_lut_3_lut_LC_15_7_7 (
            .in0(N__49506),
            .in1(_gnd_net_),
            .in2(N__50220),
            .in3(N__38976),
            .lcout(n14_adj_1168),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_262_LC_15_8_1.C_ON=1'b0;
    defparam i1_2_lut_adj_262_LC_15_8_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_262_LC_15_8_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_262_LC_15_8_1 (
            .in0(_gnd_net_),
            .in1(N__49471),
            .in2(_gnd_net_),
            .in3(N__50580),
            .lcout(n15176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12186_3_lut_LC_15_8_2.C_ON=1'b0;
    defparam i12186_3_lut_LC_15_8_2.SEQ_MODE=4'b0000;
    defparam i12186_3_lut_LC_15_8_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12186_3_lut_LC_15_8_2 (
            .in0(N__38766),
            .in1(N__44774),
            .in2(_gnd_net_),
            .in3(N__43560),
            .lcout(n15396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12817_4_lut_4_lut_LC_15_8_3.C_ON=1'b0;
    defparam i12817_4_lut_4_lut_LC_15_8_3.SEQ_MODE=4'b0000;
    defparam i12817_4_lut_4_lut_LC_15_8_3.LUT_INIT=16'b0001010000010000;
    LogicCell40 i12817_4_lut_4_lut_LC_15_8_3 (
            .in0(N__49868),
            .in1(N__49470),
            .in2(N__43439),
            .in3(N__43255),
            .lcout(n15527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_15_8_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_15_8_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_15_8_4.LUT_INIT=16'b1100110011011101;
    LogicCell40 i1_2_lut_3_lut_LC_15_8_4 (
            .in0(N__49473),
            .in1(N__52360),
            .in2(_gnd_net_),
            .in3(N__49870),
            .lcout(n8133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i34_4_lut_LC_15_8_6.C_ON=1'b0;
    defparam i34_4_lut_LC_15_8_6.SEQ_MODE=4'b0000;
    defparam i34_4_lut_LC_15_8_6.LUT_INIT=16'b1110010001000100;
    LogicCell40 i34_4_lut_LC_15_8_6 (
            .in0(N__49874),
            .in1(N__33625),
            .in2(N__31094),
            .in3(N__31082),
            .lcout(n15_adj_1203),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_3_lut_4_lut_LC_15_8_7.C_ON=1'b0;
    defparam i1_4_lut_3_lut_4_lut_LC_15_8_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_3_lut_4_lut_LC_15_8_7.LUT_INIT=16'b1110000111100000;
    LogicCell40 i1_4_lut_3_lut_4_lut_LC_15_8_7 (
            .in0(N__49869),
            .in1(N__49472),
            .in2(N__52446),
            .in3(N__50581),
            .lcout(n10566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i0_LC_15_9_0 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i0_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i0_LC_15_9_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i0_LC_15_9_0  (
            .in0(N__48518),
            .in1(N__35734),
            .in2(N__33875),
            .in3(N__31036),
            .lcout(\CLOCK_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51155),
            .ce(N__31209),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i1_LC_15_9_1 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i1_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i1_LC_15_9_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i1_LC_15_9_1  (
            .in0(N__35735),
            .in1(N__48519),
            .in2(N__31025),
            .in3(N__42125),
            .lcout(\CLOCK_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51155),
            .ce(N__31209),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i2_LC_15_9_2 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i2_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i2_LC_15_9_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i2_LC_15_9_2  (
            .in0(N__48520),
            .in1(N__35736),
            .in2(N__31016),
            .in3(N__43685),
            .lcout(\CLOCK_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51155),
            .ce(N__31209),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.i1_4_lut_LC_15_9_3 .C_ON=1'b0;
    defparam \CLOCK_DDS.i1_4_lut_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \CLOCK_DDS.i1_4_lut_LC_15_9_3 .LUT_INIT=16'b1010101000100110;
    LogicCell40 \CLOCK_DDS.i1_4_lut_LC_15_9_3  (
            .in0(N__35733),
            .in1(N__48387),
            .in2(N__33908),
            .in3(N__48517),
            .lcout(\CLOCK_DDS.n9759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i3_LC_15_9_4 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i3_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i3_LC_15_9_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i3_LC_15_9_4  (
            .in0(N__48521),
            .in1(N__35737),
            .in2(N__31262),
            .in3(N__40969),
            .lcout(\CLOCK_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51155),
            .ce(N__31209),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i4_LC_15_9_5 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i4_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i4_LC_15_9_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \CLOCK_DDS.tmp_buf_i4_LC_15_9_5  (
            .in0(N__31577),
            .in1(N__31253),
            .in2(N__35759),
            .in3(N__48522),
            .lcout(\CLOCK_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51155),
            .ce(N__31209),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i5_LC_15_9_6 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i5_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i5_LC_15_9_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i5_LC_15_9_6  (
            .in0(N__48523),
            .in1(N__35741),
            .in2(N__31244),
            .in3(N__34233),
            .lcout(\CLOCK_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51155),
            .ce(N__31209),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i6_LC_15_9_7 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i6_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i6_LC_15_9_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i6_LC_15_9_7  (
            .in0(N__35742),
            .in1(N__48524),
            .in2(N__31235),
            .in3(N__34628),
            .lcout(\CLOCK_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51155),
            .ce(N__31209),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.tmp_buf_i7_LC_15_10_0 .C_ON=1'b0;
    defparam \CLOCK_DDS.tmp_buf_i7_LC_15_10_0 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.tmp_buf_i7_LC_15_10_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLOCK_DDS.tmp_buf_i7_LC_15_10_0  (
            .in0(N__48506),
            .in1(N__35732),
            .in2(N__31226),
            .in3(N__31730),
            .lcout(\CLOCK_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51168),
            .ce(N__31211),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.i7713_3_lut_LC_15_10_1 .C_ON=1'b0;
    defparam \CLOCK_DDS.i7713_3_lut_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \CLOCK_DDS.i7713_3_lut_LC_15_10_1 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \CLOCK_DDS.i7713_3_lut_LC_15_10_1  (
            .in0(N__35728),
            .in1(N__48383),
            .in2(_gnd_net_),
            .in3(N__48503),
            .lcout(n10823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.i23_4_lut_LC_15_10_2 .C_ON=1'b0;
    defparam \CLOCK_DDS.i23_4_lut_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \CLOCK_DDS.i23_4_lut_LC_15_10_2 .LUT_INIT=16'b1111101000010101;
    LogicCell40 \CLOCK_DDS.i23_4_lut_LC_15_10_2  (
            .in0(N__48505),
            .in1(N__33896),
            .in2(N__48389),
            .in3(N__35731),
            .lcout(\CLOCK_DDS.n9_adj_1021 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.i13064_4_lut_LC_15_10_3 .C_ON=1'b0;
    defparam \CLOCK_DDS.i13064_4_lut_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \CLOCK_DDS.i13064_4_lut_LC_15_10_3 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \CLOCK_DDS.i13064_4_lut_LC_15_10_3  (
            .in0(N__35730),
            .in1(N__48382),
            .in2(N__33903),
            .in3(N__48504),
            .lcout(\CLOCK_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12766_2_lut_LC_15_10_4.C_ON=1'b0;
    defparam i12766_2_lut_LC_15_10_4.SEQ_MODE=4'b0000;
    defparam i12766_2_lut_LC_15_10_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 i12766_2_lut_LC_15_10_4 (
            .in0(_gnd_net_),
            .in1(N__31151),
            .in2(_gnd_net_),
            .in3(N__35729),
            .lcout(n15640),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i8_3_lut_LC_15_10_5.C_ON=1'b0;
    defparam mux_1498_i8_3_lut_LC_15_10_5.SEQ_MODE=4'b0000;
    defparam mux_1498_i8_3_lut_LC_15_10_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_1498_i8_3_lut_LC_15_10_5 (
            .in0(N__31729),
            .in1(N__36763),
            .in2(_gnd_net_),
            .in3(N__47702),
            .lcout(n4202),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i8_3_lut_LC_15_10_7.C_ON=1'b0;
    defparam mux_1511_i8_3_lut_LC_15_10_7.SEQ_MODE=4'b0000;
    defparam mux_1511_i8_3_lut_LC_15_10_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 mux_1511_i8_3_lut_LC_15_10_7 (
            .in0(N__31316),
            .in1(_gnd_net_),
            .in2(N__45653),
            .in3(N__33806),
            .lcout(n4247),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i7_LC_15_11_0.C_ON=1'b0;
    defparam req_data_cnt_i7_LC_15_11_0.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i7_LC_15_11_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i7_LC_15_11_0 (
            .in0(N__37318),
            .in1(N__40434),
            .in2(_gnd_net_),
            .in3(N__31336),
            .lcout(req_data_cnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51186),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i7_LC_15_11_1.C_ON=1'b0;
    defparam acadc_skipCount_i7_LC_15_11_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i7_LC_15_11_1.LUT_INIT=16'b0111010100100000;
    LogicCell40 acadc_skipCount_i7_LC_15_11_1 (
            .in0(N__41818),
            .in1(N__51915),
            .in2(N__38971),
            .in3(N__31986),
            .lcout(acadc_skipCount_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51186),
            .ce(),
            .sr(_gnd_net_));
    defparam i12655_2_lut_LC_15_11_2.C_ON=1'b0;
    defparam i12655_2_lut_LC_15_11_2.SEQ_MODE=4'b0000;
    defparam i12655_2_lut_LC_15_11_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i12655_2_lut_LC_15_11_2 (
            .in0(_gnd_net_),
            .in1(N__47810),
            .in2(_gnd_net_),
            .in3(N__31911),
            .lcout(n15556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i14_LC_15_11_3.C_ON=1'b0;
    defparam req_data_cnt_i14_LC_15_11_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i14_LC_15_11_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 req_data_cnt_i14_LC_15_11_3 (
            .in0(N__31912),
            .in1(_gnd_net_),
            .in2(N__40460),
            .in3(N__37630),
            .lcout(req_data_cnt_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51186),
            .ce(),
            .sr(_gnd_net_));
    defparam i111_4_lut_LC_15_11_4.C_ON=1'b0;
    defparam i111_4_lut_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam i111_4_lut_LC_15_11_4.LUT_INIT=16'b0011000010001000;
    LogicCell40 i111_4_lut_LC_15_11_4 (
            .in0(N__36843),
            .in1(N__45598),
            .in2(N__31553),
            .in3(N__47150),
            .lcout(n60_adj_1157),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1513_i3_4_lut_LC_15_11_5.C_ON=1'b0;
    defparam mux_1513_i3_4_lut_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam mux_1513_i3_4_lut_LC_15_11_5.LUT_INIT=16'b1011101000010000;
    LogicCell40 mux_1513_i3_4_lut_LC_15_11_5 (
            .in0(N__47151),
            .in1(N__45306),
            .in2(N__43661),
            .in3(N__31280),
            .lcout(n4262),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_299_LC_15_11_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_299_LC_15_11_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_299_LC_15_11_6.LUT_INIT=16'b1111111110101111;
    LogicCell40 i1_2_lut_3_lut_adj_299_LC_15_11_6 (
            .in0(N__50561),
            .in1(_gnd_net_),
            .in2(N__49538),
            .in3(N__49966),
            .lcout(n7567),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1513_i8_4_lut_LC_15_11_7.C_ON=1'b0;
    defparam mux_1513_i8_4_lut_LC_15_11_7.SEQ_MODE=4'b0000;
    defparam mux_1513_i8_4_lut_LC_15_11_7.LUT_INIT=16'b1011101000010000;
    LogicCell40 mux_1513_i8_4_lut_LC_15_11_7 (
            .in0(N__47152),
            .in1(N__45307),
            .in2(N__31271),
            .in3(N__31466),
            .lcout(n4257),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_15_12_0.C_ON=1'b0;
    defparam i3_4_lut_LC_15_12_0.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_15_12_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i3_4_lut_LC_15_12_0 (
            .in0(N__34889),
            .in1(N__31422),
            .in2(N__35453),
            .in3(N__31407),
            .lcout(n19_adj_1234),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i15_LC_15_12_1.C_ON=1'b0;
    defparam buf_dds_i15_LC_15_12_1.SEQ_MODE=4'b1000;
    defparam buf_dds_i15_LC_15_12_1.LUT_INIT=16'b1100000010101010;
    LogicCell40 buf_dds_i15_LC_15_12_1 (
            .in0(N__31452),
            .in1(N__38926),
            .in2(N__41511),
            .in3(N__41356),
            .lcout(buf_dds_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51204),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i13_LC_15_12_2.C_ON=1'b0;
    defparam req_data_cnt_i13_LC_15_12_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i13_LC_15_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i13_LC_15_12_2 (
            .in0(N__37663),
            .in1(N__40454),
            .in2(_gnd_net_),
            .in3(N__31423),
            .lcout(req_data_cnt_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51204),
            .ce(),
            .sr(_gnd_net_));
    defparam i12710_2_lut_LC_15_12_3.C_ON=1'b0;
    defparam i12710_2_lut_LC_15_12_3.SEQ_MODE=4'b0000;
    defparam i12710_2_lut_LC_15_12_3.LUT_INIT=16'b0000101000001010;
    LogicCell40 i12710_2_lut_LC_15_12_3 (
            .in0(N__31408),
            .in1(_gnd_net_),
            .in2(N__47918),
            .in3(_gnd_net_),
            .lcout(n15812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i7_LC_15_12_4.C_ON=1'b0;
    defparam buf_device_acadc_i7_LC_15_12_4.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i7_LC_15_12_4.LUT_INIT=16'b0011101100001000;
    LogicCell40 buf_device_acadc_i7_LC_15_12_4 (
            .in0(N__41896),
            .in1(N__31848),
            .in2(N__51739),
            .in3(N__31378),
            .lcout(buf_device_acadc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51204),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_292_LC_15_12_5.C_ON=1'b0;
    defparam i1_4_lut_adj_292_LC_15_12_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_292_LC_15_12_5.LUT_INIT=16'b1111101010001000;
    LogicCell40 i1_4_lut_adj_292_LC_15_12_5 (
            .in0(N__47816),
            .in1(N__40982),
            .in2(N__31364),
            .in3(N__41935),
            .lcout(n99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i8_3_lut_LC_15_12_7.C_ON=1'b0;
    defparam mux_1502_i8_3_lut_LC_15_12_7.SEQ_MODE=4'b0000;
    defparam mux_1502_i8_3_lut_LC_15_12_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_1502_i8_3_lut_LC_15_12_7 (
            .in0(N__47815),
            .in1(N__31335),
            .in2(_gnd_net_),
            .in3(N__31991),
            .lcout(n4214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i4_LC_15_13_0.C_ON=1'b0;
    defparam req_data_cnt_i4_LC_15_13_0.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i4_LC_15_13_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i4_LC_15_13_0 (
            .in0(N__40471),
            .in1(N__37400),
            .in2(_gnd_net_),
            .in3(N__34658),
            .lcout(req_data_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51221),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i10_LC_15_13_1.C_ON=1'b0;
    defparam req_data_cnt_i10_LC_15_13_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i10_LC_15_13_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i10_LC_15_13_1 (
            .in0(N__37190),
            .in1(N__40472),
            .in2(_gnd_net_),
            .in3(N__34177),
            .lcout(req_data_cnt_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51221),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i7_LC_15_13_2.C_ON=1'b0;
    defparam buf_dds_i7_LC_15_13_2.SEQ_MODE=4'b1000;
    defparam buf_dds_i7_LC_15_13_2.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i7_LC_15_13_2 (
            .in0(N__38972),
            .in1(N__31728),
            .in2(N__41506),
            .in3(N__41361),
            .lcout(buf_dds_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51221),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_288_LC_15_13_3.C_ON=1'b0;
    defparam i15_4_lut_adj_288_LC_15_13_3.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_288_LC_15_13_3.LUT_INIT=16'b1011000110111011;
    LogicCell40 i15_4_lut_adj_288_LC_15_13_3 (
            .in0(N__52443),
            .in1(N__31674),
            .in2(N__51737),
            .in3(N__40543),
            .lcout(n9187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_94_LC_15_13_5.C_ON=1'b0;
    defparam i5_4_lut_adj_94_LC_15_13_5.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_94_LC_15_13_5.LUT_INIT=16'b0111101111011110;
    LogicCell40 i5_4_lut_adj_94_LC_15_13_5 (
            .in0(N__34030),
            .in1(N__34820),
            .in2(N__35477),
            .in3(N__34176),
            .lcout(n21_adj_1204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i4_LC_15_13_6.C_ON=1'b0;
    defparam buf_dds_i4_LC_15_13_6.SEQ_MODE=4'b1000;
    defparam buf_dds_i4_LC_15_13_6.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i4_LC_15_13_6 (
            .in0(N__31624),
            .in1(N__31575),
            .in2(N__41505),
            .in3(N__41360),
            .lcout(buf_dds_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51221),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_5__356_LC_15_13_7.C_ON=1'b0;
    defparam buf_control_5__356_LC_15_13_7.SEQ_MODE=4'b1000;
    defparam buf_control_5__356_LC_15_13_7.LUT_INIT=16'b1100110011100100;
    LogicCell40 buf_control_5__356_LC_15_13_7 (
            .in0(N__39662),
            .in1(N__31549),
            .in2(N__33794),
            .in3(N__41151),
            .lcout(buf_control_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51221),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1494_i3_3_lut_LC_15_14_0.C_ON=1'b0;
    defparam mux_1494_i3_3_lut_LC_15_14_0.SEQ_MODE=4'b0000;
    defparam mux_1494_i3_3_lut_LC_15_14_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_1494_i3_3_lut_LC_15_14_0 (
            .in0(N__47805),
            .in1(N__37039),
            .in2(_gnd_net_),
            .in3(N__34684),
            .lcout(),
            .ltout(n4195_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i3_4_lut_LC_15_14_1.C_ON=1'b0;
    defparam mux_1507_i3_4_lut_LC_15_14_1.SEQ_MODE=4'b0000;
    defparam mux_1507_i3_4_lut_LC_15_14_1.LUT_INIT=16'b1110111011110000;
    LogicCell40 mux_1507_i3_4_lut_LC_15_14_1 (
            .in0(N__31535),
            .in1(N__47806),
            .in2(N__31520),
            .in3(N__45239),
            .lcout(n4232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_15_14_2.C_ON=1'b0;
    defparam i8_4_lut_LC_15_14_2.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_15_14_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i8_4_lut_LC_15_14_2 (
            .in0(N__31511),
            .in1(N__41656),
            .in2(N__31493),
            .in3(N__31782),
            .lcout(n24_adj_1174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i9_LC_15_14_3.C_ON=1'b0;
    defparam acadc_skipCount_i9_LC_15_14_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i9_LC_15_14_3.LUT_INIT=16'b0000101011001010;
    LogicCell40 acadc_skipCount_i9_LC_15_14_3 (
            .in0(N__31784),
            .in1(N__34594),
            .in2(N__41828),
            .in3(N__51853),
            .lcout(acadc_skipCount_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51238),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_92_LC_15_14_4.C_ON=1'b0;
    defparam i7_4_lut_adj_92_LC_15_14_4.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_92_LC_15_14_4.LUT_INIT=16'b0111110110111110;
    LogicCell40 i7_4_lut_adj_92_LC_15_14_4 (
            .in0(N__34786),
            .in1(N__31913),
            .in2(N__35429),
            .in3(N__37423),
            .lcout(n23_adj_1194),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i5_3_lut_LC_15_14_5.C_ON=1'b0;
    defparam mux_1502_i5_3_lut_LC_15_14_5.SEQ_MODE=4'b0000;
    defparam mux_1502_i5_3_lut_LC_15_14_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_1502_i5_3_lut_LC_15_14_5 (
            .in0(N__47811),
            .in1(N__34653),
            .in2(_gnd_net_),
            .in3(N__31889),
            .lcout(n4217),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i6_LC_15_14_6.C_ON=1'b0;
    defparam buf_device_acadc_i6_LC_15_14_6.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i6_LC_15_14_6.LUT_INIT=16'b0100111101000000;
    LogicCell40 buf_device_acadc_i6_LC_15_14_6 (
            .in0(N__51852),
            .in1(N__33789),
            .in2(N__31870),
            .in3(N__31798),
            .lcout(buf_device_acadc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51238),
            .ce(),
            .sr(_gnd_net_));
    defparam i13004_2_lut_LC_15_14_7.C_ON=1'b0;
    defparam i13004_2_lut_LC_15_14_7.SEQ_MODE=4'b0000;
    defparam i13004_2_lut_LC_15_14_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i13004_2_lut_LC_15_14_7 (
            .in0(N__31783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47804),
            .lcout(n15834),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i8_LC_15_15_1.C_ON=1'b0;
    defparam acadc_skipCount_i8_LC_15_15_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i8_LC_15_15_1.LUT_INIT=16'b0111010100100000;
    LogicCell40 acadc_skipCount_i8_LC_15_15_1 (
            .in0(N__41789),
            .in1(N__51880),
            .in2(N__34141),
            .in3(N__32271),
            .lcout(acadc_skipCount_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51253),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i2_LC_15_15_2.C_ON=1'b0;
    defparam acadc_skipCount_i2_LC_15_15_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i2_LC_15_15_2.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i2_LC_15_15_2 (
            .in0(N__51879),
            .in1(N__41790),
            .in2(N__31945),
            .in3(N__39996),
            .lcout(acadc_skipCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51253),
            .ce(),
            .sr(_gnd_net_));
    defparam i3173_3_lut_LC_15_15_3.C_ON=1'b0;
    defparam i3173_3_lut_LC_15_15_3.SEQ_MODE=4'b0000;
    defparam i3173_3_lut_LC_15_15_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i3173_3_lut_LC_15_15_3 (
            .in0(N__32057),
            .in1(N__37870),
            .in2(_gnd_net_),
            .in3(N__40534),
            .lcout(n8_adj_1225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_103_LC_15_15_4.C_ON=1'b0;
    defparam i4_4_lut_adj_103_LC_15_15_4.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_103_LC_15_15_4.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_adj_103_LC_15_15_4 (
            .in0(N__38166),
            .in1(N__38332),
            .in2(N__37771),
            .in3(N__42015),
            .lcout(),
            .ltout(n20_adj_1253_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_15_15_5.C_ON=1'b0;
    defparam i13_4_lut_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_15_15_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_LC_15_15_5 (
            .in0(N__34634),
            .in1(N__31760),
            .in2(N__31745),
            .in3(N__34298),
            .lcout(n29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12715_2_lut_LC_15_15_6.C_ON=1'b0;
    defparam i12715_2_lut_LC_15_15_6.SEQ_MODE=4'b0000;
    defparam i12715_2_lut_LC_15_15_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12715_2_lut_LC_15_15_6 (
            .in0(_gnd_net_),
            .in1(N__34134),
            .in2(_gnd_net_),
            .in3(N__32125),
            .lcout(n15546),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i23_LC_15_15_7 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i23_LC_15_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i23_LC_15_15_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i23_LC_15_15_7  (
            .in0(N__53605),
            .in1(N__46082),
            .in2(N__34470),
            .in3(N__53481),
            .lcout(cmd_rdadctmp_23_adj_1053),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51253),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i5_LC_15_16_1.C_ON=1'b0;
    defparam data_index_i5_LC_15_16_1.SEQ_MODE=4'b1000;
    defparam data_index_i5_LC_15_16_1.LUT_INIT=16'b0011000010101010;
    LogicCell40 data_index_i5_LC_15_16_1 (
            .in0(N__51508),
            .in1(N__51869),
            .in2(N__52489),
            .in3(N__52184),
            .lcout(data_index_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51270),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i6_LC_15_16_2.C_ON=1'b0;
    defparam acadc_skipCount_i6_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i6_LC_15_16_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i6_LC_15_16_2 (
            .in0(N__41820),
            .in1(N__33961),
            .in2(N__51917),
            .in3(N__34759),
            .lcout(acadc_skipCount_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51270),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i12_LC_15_16_3.C_ON=1'b0;
    defparam buf_dds_i12_LC_15_16_3.SEQ_MODE=4'b1000;
    defparam buf_dds_i12_LC_15_16_3.LUT_INIT=16'b1000100011110000;
    LogicCell40 buf_dds_i12_LC_15_16_3 (
            .in0(N__36995),
            .in1(N__41510),
            .in2(N__32031),
            .in3(N__41374),
            .lcout(buf_dds_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51270),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_15_16_4.C_ON=1'b0;
    defparam i6_4_lut_LC_15_16_4.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_15_16_4.LUT_INIT=16'b0111110110111110;
    LogicCell40 i6_4_lut_LC_15_16_4 (
            .in0(N__32009),
            .in1(N__31987),
            .in2(N__31967),
            .in3(N__31935),
            .lcout(n22_adj_1170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i3_LC_15_16_5.C_ON=1'b0;
    defparam req_data_cnt_i3_LC_15_16_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i3_LC_15_16_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 req_data_cnt_i3_LC_15_16_5 (
            .in0(N__51867),
            .in1(N__40470),
            .in2(N__44775),
            .in3(N__38170),
            .lcout(req_data_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51270),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i10_LC_15_16_6.C_ON=1'b0;
    defparam acadc_skipCount_i10_LC_15_16_6.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i10_LC_15_16_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i10_LC_15_16_6 (
            .in0(N__41819),
            .in1(N__34424),
            .in2(N__51916),
            .in3(N__34210),
            .lcout(acadc_skipCount_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51270),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i13_LC_15_16_7.C_ON=1'b0;
    defparam acadc_skipCount_i13_LC_15_16_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i13_LC_15_16_7.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i13_LC_15_16_7 (
            .in0(N__51866),
            .in1(N__41821),
            .in2(N__32215),
            .in3(N__33793),
            .lcout(acadc_skipCount_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51270),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_3_i15_4_lut_LC_15_17_0.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_3_i15_4_lut_LC_15_17_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_3_i15_4_lut_LC_15_17_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_394_Mux_3_i15_4_lut_LC_15_17_0 (
            .in0(N__52466),
            .in1(N__32500),
            .in2(N__51913),
            .in3(N__32488),
            .lcout(data_index_9_N_258_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13054_3_lut_4_lut_LC_15_17_2.C_ON=1'b0;
    defparam i13054_3_lut_4_lut_LC_15_17_2.SEQ_MODE=4'b0000;
    defparam i13054_3_lut_4_lut_LC_15_17_2.LUT_INIT=16'b0000000000000111;
    LogicCell40 i13054_3_lut_4_lut_LC_15_17_2 (
            .in0(N__32833),
            .in1(N__32926),
            .in2(N__32767),
            .in3(N__38127),
            .lcout(n8456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i3_LC_15_17_3.C_ON=1'b0;
    defparam acadc_skipCount_i3_LC_15_17_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i3_LC_15_17_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i3_LC_15_17_3 (
            .in0(N__51868),
            .in1(N__41822),
            .in2(N__44777),
            .in3(N__38146),
            .lcout(acadc_skipCount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51282),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i5_LC_15_17_4.C_ON=1'b0;
    defparam acadc_skipCount_i5_LC_15_17_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i5_LC_15_17_4.LUT_INIT=16'b0000110010101010;
    LogicCell40 acadc_skipCount_i5_LC_15_17_4 (
            .in0(N__37741),
            .in1(N__37882),
            .in2(N__51914),
            .in3(N__41823),
            .lcout(acadc_skipCount_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51282),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_15_17_5.C_ON=1'b0;
    defparam i4_4_lut_LC_15_17_5.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_15_17_5.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_LC_15_17_5 (
            .in0(N__32323),
            .in1(N__37740),
            .in2(N__32309),
            .in3(N__38145),
            .lcout(),
            .ltout(n20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_15_17_6.C_ON=1'b0;
    defparam i10_4_lut_LC_15_17_6.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_15_17_6.LUT_INIT=16'b1111111111110110;
    LogicCell40 i10_4_lut_LC_15_17_6 (
            .in0(N__32291),
            .in1(N__32272),
            .in2(N__32249),
            .in3(N__32189),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_46_i14_2_lut_LC_15_17_7.C_ON=1'b0;
    defparam equal_46_i14_2_lut_LC_15_17_7.SEQ_MODE=4'b0000;
    defparam equal_46_i14_2_lut_LC_15_17_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 equal_46_i14_2_lut_LC_15_17_7 (
            .in0(_gnd_net_),
            .in1(N__32234),
            .in2(_gnd_net_),
            .in3(N__32205),
            .lcout(n14_adj_1160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i8_LC_15_18_4 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i8_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i8_LC_15_18_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i8_LC_15_18_4  (
            .in0(N__53101),
            .in1(N__32140),
            .in2(N__32183),
            .in3(N__52897),
            .lcout(buf_adcdata1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51293),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_LC_15_18_7.C_ON=1'b0;
    defparam i2_4_lut_4_lut_LC_15_18_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_LC_15_18_7.LUT_INIT=16'b0000001000000011;
    LogicCell40 i2_4_lut_4_lut_LC_15_18_7 (
            .in0(N__32930),
            .in1(N__32834),
            .in2(N__32763),
            .in3(N__38132),
            .lcout(n9790),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i8_LC_15_19_0.C_ON=1'b0;
    defparam data_index_i8_LC_15_19_0.SEQ_MODE=4'b1000;
    defparam data_index_i8_LC_15_19_0.LUT_INIT=16'b0100111001000100;
    LogicCell40 data_index_i8_LC_15_19_0 (
            .in0(N__52469),
            .in1(N__42580),
            .in2(N__51931),
            .in3(N__42601),
            .lcout(data_index_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51302),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.dds_state_i2_LC_16_4_6 .C_ON=1'b0;
    defparam \CLOCK_DDS.dds_state_i2_LC_16_4_6 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.dds_state_i2_LC_16_4_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \CLOCK_DDS.dds_state_i2_LC_16_4_6  (
            .in0(_gnd_net_),
            .in1(N__35669),
            .in2(_gnd_net_),
            .in3(N__48420),
            .lcout(dds_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51117),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1481_i4_4_lut_LC_16_5_0.C_ON=1'b0;
    defparam mux_1481_i4_4_lut_LC_16_5_0.SEQ_MODE=4'b0000;
    defparam mux_1481_i4_4_lut_LC_16_5_0.LUT_INIT=16'b1010001110100000;
    LogicCell40 mux_1481_i4_4_lut_LC_16_5_0 (
            .in0(N__32633),
            .in1(N__48048),
            .in2(N__47309),
            .in3(N__32623),
            .lcout(n4149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_16_5_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_16_5_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_102_2_lut_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(N__32564),
            .in2(_gnd_net_),
            .in3(N__46561),
            .lcout(\comm_spi.data_tx_7__N_819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i1_LC_16_6_0.C_ON=1'b0;
    defparam comm_index_i1_LC_16_6_0.SEQ_MODE=4'b1000;
    defparam comm_index_i1_LC_16_6_0.LUT_INIT=16'b1101111100100000;
    LogicCell40 comm_index_i1_LC_16_6_0 (
            .in0(N__43298),
            .in1(N__43441),
            .in2(N__38693),
            .in3(N__33020),
            .lcout(comm_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51132),
            .ce(N__32522),
            .sr(N__33693));
    defparam comm_index_i0_LC_16_6_1.C_ON=1'b0;
    defparam comm_index_i0_LC_16_6_1.SEQ_MODE=4'b1000;
    defparam comm_index_i0_LC_16_6_1.LUT_INIT=16'b1001100111001100;
    LogicCell40 comm_index_i0_LC_16_6_1 (
            .in0(N__43440),
            .in1(N__38642),
            .in2(_gnd_net_),
            .in3(N__43297),
            .lcout(comm_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51132),
            .ce(N__32522),
            .sr(N__33693));
    defparam i12636_3_lut_4_lut_LC_16_7_0.C_ON=1'b0;
    defparam i12636_3_lut_4_lut_LC_16_7_0.SEQ_MODE=4'b0000;
    defparam i12636_3_lut_4_lut_LC_16_7_0.LUT_INIT=16'b1100100011000000;
    LogicCell40 i12636_3_lut_4_lut_LC_16_7_0 (
            .in0(N__40237),
            .in1(N__45302),
            .in2(N__33559),
            .in3(N__47236),
            .lcout(n15463),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12637_3_lut_4_lut_LC_16_7_1.C_ON=1'b0;
    defparam i12637_3_lut_4_lut_LC_16_7_1.SEQ_MODE=4'b0000;
    defparam i12637_3_lut_4_lut_LC_16_7_1.LUT_INIT=16'b1110000011000000;
    LogicCell40 i12637_3_lut_4_lut_LC_16_7_1 (
            .in0(N__47237),
            .in1(N__33371),
            .in2(N__45313),
            .in3(N__40238),
            .lcout(),
            .ltout(n15460_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i39_4_lut_adj_64_LC_16_7_2.C_ON=1'b0;
    defparam i39_4_lut_adj_64_LC_16_7_2.SEQ_MODE=4'b0000;
    defparam i39_4_lut_adj_64_LC_16_7_2.LUT_INIT=16'b1111000001000100;
    LogicCell40 i39_4_lut_adj_64_LC_16_7_2 (
            .in0(N__33649),
            .in1(N__33372),
            .in2(N__33596),
            .in3(N__45604),
            .lcout(),
            .ltout(n19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i3_LC_16_7_3.C_ON=1'b0;
    defparam comm_length_i3_LC_16_7_3.SEQ_MODE=4'b1000;
    defparam comm_length_i3_LC_16_7_3.LUT_INIT=16'b1011101000110000;
    LogicCell40 comm_length_i3_LC_16_7_3 (
            .in0(N__33373),
            .in1(N__47852),
            .in2(N__33593),
            .in3(N__36586),
            .lcout(comm_length_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51144),
            .ce(N__50660),
            .sr(N__33700));
    defparam i39_4_lut_LC_16_7_4.C_ON=1'b0;
    defparam i39_4_lut_LC_16_7_4.SEQ_MODE=4'b0000;
    defparam i39_4_lut_LC_16_7_4.LUT_INIT=16'b1100110000001010;
    LogicCell40 i39_4_lut_LC_16_7_4 (
            .in0(N__33555),
            .in1(N__33590),
            .in2(N__33650),
            .in3(N__45603),
            .lcout(),
            .ltout(n19_adj_1151_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i2_LC_16_7_5.C_ON=1'b0;
    defparam comm_length_i2_LC_16_7_5.SEQ_MODE=4'b1000;
    defparam comm_length_i2_LC_16_7_5.LUT_INIT=16'b1011101111111011;
    LogicCell40 comm_length_i2_LC_16_7_5 (
            .in0(N__33584),
            .in1(N__38996),
            .in2(N__33569),
            .in3(N__47853),
            .lcout(comm_length_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51144),
            .ce(N__50660),
            .sr(N__33700));
    defparam i2_4_lut_adj_281_LC_16_7_6.C_ON=1'b0;
    defparam i2_4_lut_adj_281_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_281_LC_16_7_6.LUT_INIT=16'b0110111111110110;
    LogicCell40 i2_4_lut_adj_281_LC_16_7_6 (
            .in0(N__33551),
            .in1(N__33486),
            .in2(N__33374),
            .in3(N__33320),
            .lcout(),
            .ltout(n6_adj_1281_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_283_LC_16_7_7.C_ON=1'b0;
    defparam i3_4_lut_adj_283_LC_16_7_7.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_283_LC_16_7_7.LUT_INIT=16'b1111110111111110;
    LogicCell40 i3_4_lut_adj_283_LC_16_7_7 (
            .in0(N__33715),
            .in1(N__32948),
            .in2(N__33215),
            .in3(N__38630),
            .lcout(n7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_200_i2_2_lut_LC_16_8_0.C_ON=1'b0;
    defparam equal_200_i2_2_lut_LC_16_8_0.SEQ_MODE=4'b0000;
    defparam equal_200_i2_2_lut_LC_16_8_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 equal_200_i2_2_lut_LC_16_8_0 (
            .in0(_gnd_net_),
            .in1(N__32938),
            .in2(_gnd_net_),
            .in3(N__33085),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_55_LC_16_8_1.C_ON=1'b0;
    defparam i1_4_lut_adj_55_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_55_LC_16_8_1.LUT_INIT=16'b1111010111000100;
    LogicCell40 i1_4_lut_adj_55_LC_16_8_1 (
            .in0(N__32939),
            .in1(N__40910),
            .in2(N__39475),
            .in3(N__41221),
            .lcout(),
            .ltout(n15119_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i1_LC_16_8_2.C_ON=1'b0;
    defparam comm_length_i1_LC_16_8_2.SEQ_MODE=4'b1000;
    defparam comm_length_i1_LC_16_8_2.LUT_INIT=16'b0111111111111111;
    LogicCell40 comm_length_i1_LC_16_8_2 (
            .in0(N__36605),
            .in1(N__40925),
            .in2(N__32942),
            .in3(N__33728),
            .lcout(comm_length_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51156),
            .ce(N__50656),
            .sr(N__33692));
    defparam i1_2_lut_3_lut_4_lut_LC_16_8_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_16_8_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_16_8_3.LUT_INIT=16'b1110111111101010;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_16_8_3 (
            .in0(N__40880),
            .in1(N__44969),
            .in2(N__47232),
            .in3(N__43198),
            .lcout(n5_adj_1282),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_209_i13_2_lut_3_lut_LC_16_8_4.C_ON=1'b0;
    defparam equal_209_i13_2_lut_3_lut_LC_16_8_4.SEQ_MODE=4'b0000;
    defparam equal_209_i13_2_lut_3_lut_LC_16_8_4.LUT_INIT=16'b1111111110111011;
    LogicCell40 equal_209_i13_2_lut_3_lut_LC_16_8_4 (
            .in0(N__43197),
            .in1(N__47095),
            .in2(_gnd_net_),
            .in3(N__40879),
            .lcout(n13),
            .ltout(n13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_54_LC_16_8_5.C_ON=1'b0;
    defparam i1_2_lut_adj_54_LC_16_8_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_54_LC_16_8_5.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_54_LC_16_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33731),
            .in3(N__38995),
            .lcout(n6_adj_1273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i0_LC_16_8_6.C_ON=1'b0;
    defparam comm_length_i0_LC_16_8_6.SEQ_MODE=4'b1000;
    defparam comm_length_i0_LC_16_8_6.LUT_INIT=16'b0101110111111111;
    LogicCell40 comm_length_i0_LC_16_8_6 (
            .in0(N__33722),
            .in1(N__33716),
            .in2(N__39476),
            .in3(N__41166),
            .lcout(comm_length_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51156),
            .ce(N__50656),
            .sr(N__33692));
    defparam i1_4_lut_adj_209_LC_16_8_7.C_ON=1'b0;
    defparam i1_4_lut_adj_209_LC_16_8_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_209_LC_16_8_7.LUT_INIT=16'b1111000000010000;
    LogicCell40 i1_4_lut_adj_209_LC_16_8_7 (
            .in0(N__50536),
            .in1(N__33656),
            .in2(N__52447),
            .in3(N__51841),
            .lcout(n8253),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9554_2_lut_LC_16_9_0.C_ON=1'b0;
    defparam i9554_2_lut_LC_16_9_0.SEQ_MODE=4'b0000;
    defparam i9554_2_lut_LC_16_9_0.LUT_INIT=16'b1110111011101110;
    LogicCell40 i9554_2_lut_LC_16_9_0 (
            .in0(N__47047),
            .in1(N__45229),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n12649),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_250_LC_16_9_1.C_ON=1'b0;
    defparam i1_4_lut_adj_250_LC_16_9_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_250_LC_16_9_1.LUT_INIT=16'b1010101100000000;
    LogicCell40 i1_4_lut_adj_250_LC_16_9_1 (
            .in0(N__52217),
            .in1(N__49531),
            .in2(N__42755),
            .in3(N__36595),
            .lcout(n8525),
            .ltout(n8525_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i5_LC_16_9_2.C_ON=1'b0;
    defparam buf_dds_i5_LC_16_9_2.SEQ_MODE=4'b1000;
    defparam buf_dds_i5_LC_16_9_2.LUT_INIT=16'b1010110011111100;
    LogicCell40 buf_dds_i5_LC_16_9_2 (
            .in0(N__37369),
            .in1(N__34234),
            .in2(N__33635),
            .in3(N__52218),
            .lcout(buf_dds_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51169),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_230_LC_16_9_3.C_ON=1'b0;
    defparam i1_4_lut_adj_230_LC_16_9_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_230_LC_16_9_3.LUT_INIT=16'b1010000010001000;
    LogicCell40 i1_4_lut_adj_230_LC_16_9_3 (
            .in0(N__40212),
            .in1(N__39590),
            .in2(N__36566),
            .in3(N__47046),
            .lcout(n4075),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds_333_LC_16_9_4.C_ON=1'b0;
    defparam trig_dds_333_LC_16_9_4.SEQ_MODE=4'b1000;
    defparam trig_dds_333_LC_16_9_4.LUT_INIT=16'b1111100001110000;
    LogicCell40 trig_dds_333_LC_16_9_4 (
            .in0(N__36596),
            .in1(N__33914),
            .in2(N__33907),
            .in3(N__41498),
            .lcout(trig_dds),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51169),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i0_LC_16_9_5.C_ON=1'b0;
    defparam buf_dds_i0_LC_16_9_5.SEQ_MODE=4'b1000;
    defparam buf_dds_i0_LC_16_9_5.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i0_LC_16_9_5 (
            .in0(N__36716),
            .in1(N__33870),
            .in2(N__41520),
            .in3(N__41313),
            .lcout(buf_dds_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51169),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i8_LC_16_9_6.C_ON=1'b0;
    defparam buf_dds_i8_LC_16_9_6.SEQ_MODE=4'b1000;
    defparam buf_dds_i8_LC_16_9_6.LUT_INIT=16'b1101100001010000;
    LogicCell40 buf_dds_i8_LC_16_9_6 (
            .in0(N__41312),
            .in1(N__34133),
            .in2(N__33850),
            .in3(N__41497),
            .lcout(buf_dds_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51169),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1494_i8_3_lut_LC_16_10_1.C_ON=1'b0;
    defparam mux_1494_i8_3_lut_LC_16_10_1.SEQ_MODE=4'b0000;
    defparam mux_1494_i8_3_lut_LC_16_10_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_1494_i8_3_lut_LC_16_10_1 (
            .in0(N__37298),
            .in1(N__47700),
            .in2(_gnd_net_),
            .in3(N__34921),
            .lcout(),
            .ltout(n4190_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i8_4_lut_LC_16_10_2.C_ON=1'b0;
    defparam mux_1507_i8_4_lut_LC_16_10_2.SEQ_MODE=4'b0000;
    defparam mux_1507_i8_4_lut_LC_16_10_2.LUT_INIT=16'b1110111011110000;
    LogicCell40 mux_1507_i8_4_lut_LC_16_10_2 (
            .in0(N__47701),
            .in1(N__33821),
            .in2(N__33809),
            .in3(N__45240),
            .lcout(n4227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i2_LC_16_10_3.C_ON=1'b0;
    defparam comm_buf_1__i2_LC_16_10_3.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i2_LC_16_10_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i2_LC_16_10_3 (
            .in0(N__40116),
            .in1(N__50123),
            .in2(_gnd_net_),
            .in3(N__33800),
            .lcout(comm_buf_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51187),
            .ce(N__44711),
            .sr(N__44653));
    defparam i9634_2_lut_3_lut_LC_16_10_5.C_ON=1'b0;
    defparam i9634_2_lut_3_lut_LC_16_10_5.SEQ_MODE=4'b0000;
    defparam i9634_2_lut_3_lut_LC_16_10_5.LUT_INIT=16'b0000000001000100;
    LogicCell40 i9634_2_lut_3_lut_LC_16_10_5 (
            .in0(N__49546),
            .in1(N__39970),
            .in2(_gnd_net_),
            .in3(N__50120),
            .lcout(n14_adj_1197),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9627_2_lut_3_lut_LC_16_10_6.C_ON=1'b0;
    defparam i9627_2_lut_3_lut_LC_16_10_6.SEQ_MODE=4'b0000;
    defparam i9627_2_lut_3_lut_LC_16_10_6.LUT_INIT=16'b0000000001000100;
    LogicCell40 i9627_2_lut_3_lut_LC_16_10_6 (
            .in0(N__50121),
            .in1(N__34592),
            .in2(_gnd_net_),
            .in3(N__49547),
            .lcout(n14_adj_1210),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9628_2_lut_3_lut_LC_16_10_7.C_ON=1'b0;
    defparam i9628_2_lut_3_lut_LC_16_10_7.SEQ_MODE=4'b0000;
    defparam i9628_2_lut_3_lut_LC_16_10_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i9628_2_lut_3_lut_LC_16_10_7 (
            .in0(N__49548),
            .in1(N__34409),
            .in2(_gnd_net_),
            .in3(N__50122),
            .lcout(n14_adj_1209),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9638_2_lut_3_lut_LC_16_11_1.C_ON=1'b0;
    defparam i9638_2_lut_3_lut_LC_16_11_1.SEQ_MODE=4'b0000;
    defparam i9638_2_lut_3_lut_LC_16_11_1.LUT_INIT=16'b0000000001000100;
    LogicCell40 i9638_2_lut_3_lut_LC_16_11_1 (
            .in0(N__49819),
            .in1(N__33775),
            .in2(_gnd_net_),
            .in3(N__49549),
            .lcout(n14_adj_1202),
            .ltout(n14_adj_1202_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i13_LC_16_11_2.C_ON=1'b0;
    defparam buf_dds_i13_LC_16_11_2.SEQ_MODE=4'b1000;
    defparam buf_dds_i13_LC_16_11_2.LUT_INIT=16'b1111010111001100;
    LogicCell40 buf_dds_i13_LC_16_11_2 (
            .in0(N__52300),
            .in1(N__34060),
            .in2(N__34070),
            .in3(N__41346),
            .lcout(buf_dds_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51205),
            .ce(),
            .sr(_gnd_net_));
    defparam i12856_2_lut_LC_16_11_3.C_ON=1'b0;
    defparam i12856_2_lut_LC_16_11_3.SEQ_MODE=4'b0000;
    defparam i12856_2_lut_LC_16_11_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12856_2_lut_LC_16_11_3 (
            .in0(N__34059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47824),
            .lcout(n15690),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i12_LC_16_11_4.C_ON=1'b0;
    defparam req_data_cnt_i12_LC_16_11_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i12_LC_16_11_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i12_LC_16_11_4 (
            .in0(N__40433),
            .in1(N__37718),
            .in2(_gnd_net_),
            .in3(N__34029),
            .lcout(req_data_cnt_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51205),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_206_i13_2_lut_3_lut_LC_16_11_5.C_ON=1'b0;
    defparam equal_206_i13_2_lut_3_lut_LC_16_11_5.SEQ_MODE=4'b0000;
    defparam equal_206_i13_2_lut_3_lut_LC_16_11_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 equal_206_i13_2_lut_3_lut_LC_16_11_5 (
            .in0(N__43199),
            .in1(N__47027),
            .in2(_gnd_net_),
            .in3(N__40875),
            .lcout(n13_adj_1026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_71_LC_16_11_6.C_ON=1'b0;
    defparam i1_4_lut_adj_71_LC_16_11_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_71_LC_16_11_6.LUT_INIT=16'b1110101011000000;
    LogicCell40 i1_4_lut_adj_71_LC_16_11_6 (
            .in0(N__34507),
            .in1(N__45597),
            .in2(N__37214),
            .in3(N__45264),
            .lcout(),
            .ltout(n78_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_77_LC_16_11_7.C_ON=1'b0;
    defparam i1_4_lut_adj_77_LC_16_11_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_77_LC_16_11_7.LUT_INIT=16'b1110111011000000;
    LogicCell40 i1_4_lut_adj_77_LC_16_11_7 (
            .in0(N__34001),
            .in1(N__47823),
            .in2(N__33992),
            .in3(N__41931),
            .lcout(n99_adj_1024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i7_LC_16_12_0.C_ON=1'b0;
    defparam comm_buf_1__i7_LC_16_12_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i7_LC_16_12_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i7_LC_16_12_0 (
            .in0(N__39361),
            .in1(N__50152),
            .in2(_gnd_net_),
            .in3(N__33977),
            .lcout(comm_buf_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51222),
            .ce(N__44712),
            .sr(N__44641));
    defparam comm_buf_1__i0_LC_16_12_1.C_ON=1'b0;
    defparam comm_buf_1__i0_LC_16_12_1.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i0_LC_16_12_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_1__i0_LC_16_12_1 (
            .in0(N__50149),
            .in1(N__39187),
            .in2(_gnd_net_),
            .in3(N__37088),
            .lcout(comm_buf_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51222),
            .ce(N__44712),
            .sr(N__44641));
    defparam comm_buf_1__i6_LC_16_12_2.C_ON=1'b0;
    defparam comm_buf_1__i6_LC_16_12_2.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i6_LC_16_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i6_LC_16_12_2 (
            .in0(N__40715),
            .in1(N__50151),
            .in2(_gnd_net_),
            .in3(N__34703),
            .lcout(comm_buf_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51222),
            .ce(N__44712),
            .sr(N__44641));
    defparam comm_buf_1__i1_LC_16_12_3.C_ON=1'b0;
    defparam comm_buf_1__i1_LC_16_12_3.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i1_LC_16_12_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_1__i1_LC_16_12_3 (
            .in0(N__50150),
            .in1(N__44158),
            .in2(_gnd_net_),
            .in3(N__42137),
            .lcout(comm_buf_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51222),
            .ce(N__44712),
            .sr(N__44641));
    defparam i105_4_lut_LC_16_13_0.C_ON=1'b0;
    defparam i105_4_lut_LC_16_13_0.SEQ_MODE=4'b0000;
    defparam i105_4_lut_LC_16_13_0.LUT_INIT=16'b0100010010100000;
    LogicCell40 i105_4_lut_LC_16_13_0 (
            .in0(N__45233),
            .in1(N__37649),
            .in2(N__34268),
            .in3(N__47744),
            .lcout(n66_adj_1158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i6_3_lut_LC_16_13_1.C_ON=1'b0;
    defparam mux_1498_i6_3_lut_LC_16_13_1.SEQ_MODE=4'b0000;
    defparam mux_1498_i6_3_lut_LC_16_13_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_1498_i6_3_lut_LC_16_13_1 (
            .in0(N__47745),
            .in1(_gnd_net_),
            .in2(N__34238),
            .in3(N__37512),
            .lcout(n4204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_228_LC_16_13_2.C_ON=1'b0;
    defparam i1_2_lut_adj_228_LC_16_13_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_228_LC_16_13_2.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_adj_228_LC_16_13_2 (
            .in0(N__45231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47742),
            .lcout(n93),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i130_3_lut_adj_85_LC_16_13_3.C_ON=1'b0;
    defparam i130_3_lut_adj_85_LC_16_13_3.SEQ_MODE=4'b0000;
    defparam i130_3_lut_adj_85_LC_16_13_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 i130_3_lut_adj_85_LC_16_13_3 (
            .in0(N__34186),
            .in1(N__45230),
            .in2(_gnd_net_),
            .in3(N__34214),
            .lcout(n90_adj_1167),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_215_LC_16_13_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_215_LC_16_13_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_215_LC_16_13_4.LUT_INIT=16'b0000000001000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_215_LC_16_13_4 (
            .in0(N__44963),
            .in1(N__47174),
            .in2(N__39664),
            .in3(N__40885),
            .lcout(n7485),
            .ltout(n7485_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam tacadc_rst_364_LC_16_13_5.C_ON=1'b0;
    defparam tacadc_rst_364_LC_16_13_5.SEQ_MODE=4'b1000;
    defparam tacadc_rst_364_LC_16_13_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 tacadc_rst_364_LC_16_13_5 (
            .in0(N__34187),
            .in1(_gnd_net_),
            .in2(N__34190),
            .in3(N__34419),
            .lcout(tacadc_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51239),
            .ce(),
            .sr(_gnd_net_));
    defparam i125_4_lut_LC_16_13_6.C_ON=1'b0;
    defparam i125_4_lut_LC_16_13_6.SEQ_MODE=4'b0000;
    defparam i125_4_lut_LC_16_13_6.LUT_INIT=16'b1111000010001000;
    LogicCell40 i125_4_lut_LC_16_13_6 (
            .in0(N__45232),
            .in1(N__34178),
            .in2(N__34163),
            .in3(N__47743),
            .lcout(n72_adj_1162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_start_366_LC_16_13_7.C_ON=1'b0;
    defparam eis_start_366_LC_16_13_7.SEQ_MODE=4'b1000;
    defparam eis_start_366_LC_16_13_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_start_366_LC_16_13_7 (
            .in0(N__34142),
            .in1(N__34519),
            .in2(_gnd_net_),
            .in3(N__41044),
            .lcout(eis_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51239),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_109_LC_16_14_0.C_ON=1'b0;
    defparam i2_4_lut_adj_109_LC_16_14_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_109_LC_16_14_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_109_LC_16_14_0 (
            .in0(N__42159),
            .in1(N__37811),
            .in2(N__34657),
            .in3(N__38228),
            .lcout(n18_adj_1217),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i7_3_lut_LC_16_14_1.C_ON=1'b0;
    defparam mux_1498_i7_3_lut_LC_16_14_1.SEQ_MODE=4'b0000;
    defparam mux_1498_i7_3_lut_LC_16_14_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_1498_i7_3_lut_LC_16_14_1 (
            .in0(N__47920),
            .in1(_gnd_net_),
            .in2(N__34624),
            .in3(N__41557),
            .lcout(n4203),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_stop_365_LC_16_14_2.C_ON=1'b0;
    defparam eis_stop_365_LC_16_14_2.SEQ_MODE=4'b1000;
    defparam eis_stop_365_LC_16_14_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_stop_365_LC_16_14_2 (
            .in0(N__34595),
            .in1(N__34523),
            .in2(_gnd_net_),
            .in3(N__34506),
            .lcout(eis_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51254),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i15_LC_16_14_4 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i15_LC_16_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i15_LC_16_14_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i15_LC_16_14_4  (
            .in0(N__53809),
            .in1(N__34441),
            .in2(N__34474),
            .in3(N__53433),
            .lcout(buf_adcdata2_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51254),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i10_LC_16_14_5.C_ON=1'b0;
    defparam buf_dds_i10_LC_16_14_5.SEQ_MODE=4'b1000;
    defparam buf_dds_i10_LC_16_14_5.LUT_INIT=16'b1000111110000000;
    LogicCell40 buf_dds_i10_LC_16_14_5 (
            .in0(N__34423),
            .in1(N__41525),
            .in2(N__41381),
            .in3(N__34341),
            .lcout(buf_dds_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51254),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i1_3_lut_LC_16_14_7.C_ON=1'b0;
    defparam mux_1502_i1_3_lut_LC_16_14_7.SEQ_MODE=4'b0000;
    defparam mux_1502_i1_3_lut_LC_16_14_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_1502_i1_3_lut_LC_16_14_7 (
            .in0(N__47919),
            .in1(N__34322),
            .in2(_gnd_net_),
            .in3(N__34285),
            .lcout(n4221),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_112_LC_16_15_0.C_ON=1'b0;
    defparam i1_4_lut_adj_112_LC_16_15_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_112_LC_16_15_0.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_112_LC_16_15_0 (
            .in0(N__34945),
            .in1(N__36648),
            .in2(N__37922),
            .in3(N__34284),
            .lcout(n17_adj_1214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i5_LC_16_15_1.C_ON=1'b0;
    defparam req_data_cnt_i5_LC_16_15_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i5_LC_16_15_1.LUT_INIT=16'b0101000011011000;
    LogicCell40 req_data_cnt_i5_LC_16_15_1 (
            .in0(N__40458),
            .in1(N__37874),
            .in2(N__37772),
            .in3(N__51895),
            .lcout(req_data_cnt_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51271),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i0_LC_16_15_2.C_ON=1'b0;
    defparam req_data_cnt_i0_LC_16_15_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i0_LC_16_15_2.LUT_INIT=16'b0111010000110000;
    LogicCell40 req_data_cnt_i0_LC_16_15_2 (
            .in0(N__51894),
            .in1(N__40459),
            .in2(N__34292),
            .in3(N__36713),
            .lcout(req_data_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51271),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i7_3_lut_LC_16_15_3.C_ON=1'b0;
    defparam mux_1502_i7_3_lut_LC_16_15_3.SEQ_MODE=4'b0000;
    defparam mux_1502_i7_3_lut_LC_16_15_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_1502_i7_3_lut_LC_16_15_3 (
            .in0(N__47922),
            .in1(N__34758),
            .in2(_gnd_net_),
            .in3(N__37921),
            .lcout(n4215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1494_i7_3_lut_LC_16_15_4.C_ON=1'b0;
    defparam mux_1494_i7_3_lut_LC_16_15_4.SEQ_MODE=4'b0000;
    defparam mux_1494_i7_3_lut_LC_16_15_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_1494_i7_3_lut_LC_16_15_4 (
            .in0(N__37346),
            .in1(N__47923),
            .in2(_gnd_net_),
            .in3(N__34944),
            .lcout(),
            .ltout(n4191_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i7_4_lut_LC_16_15_5.C_ON=1'b0;
    defparam mux_1507_i7_4_lut_LC_16_15_5.SEQ_MODE=4'b0000;
    defparam mux_1507_i7_4_lut_LC_16_15_5.LUT_INIT=16'b1110111011110000;
    LogicCell40 mux_1507_i7_4_lut_LC_16_15_5 (
            .in0(N__47924),
            .in1(N__34739),
            .in2(N__34724),
            .in3(N__45295),
            .lcout(),
            .ltout(n4228_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i7_3_lut_LC_16_15_6.C_ON=1'b0;
    defparam mux_1511_i7_3_lut_LC_16_15_6.SEQ_MODE=4'b0000;
    defparam mux_1511_i7_3_lut_LC_16_15_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_1511_i7_3_lut_LC_16_15_6 (
            .in0(_gnd_net_),
            .in1(N__34721),
            .in2(N__34715),
            .in3(N__45649),
            .lcout(),
            .ltout(n4248_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1513_i7_4_lut_LC_16_15_7.C_ON=1'b0;
    defparam mux_1513_i7_4_lut_LC_16_15_7.SEQ_MODE=4'b0000;
    defparam mux_1513_i7_4_lut_LC_16_15_7.LUT_INIT=16'b1100000011100010;
    LogicCell40 mux_1513_i7_4_lut_LC_16_15_7 (
            .in0(N__34712),
            .in1(N__47173),
            .in2(N__34706),
            .in3(N__45296),
            .lcout(n4258),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_cntvec_i0_i0_LC_16_16_0.C_ON=1'b1;
    defparam data_cntvec_i0_i0_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i0_LC_16_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i0_LC_16_16_0 (
            .in0(_gnd_net_),
            .in1(N__36649),
            .in2(_gnd_net_),
            .in3(N__34694),
            .lcout(data_cntvec_0),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(n13951),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i1_LC_16_16_1.C_ON=1'b1;
    defparam data_cntvec_i0_i1_LC_16_16_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i1_LC_16_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i1_LC_16_16_1 (
            .in0(_gnd_net_),
            .in1(N__38227),
            .in2(_gnd_net_),
            .in3(N__34691),
            .lcout(data_cntvec_1),
            .ltout(),
            .carryin(n13951),
            .carryout(n13952),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i2_LC_16_16_2.C_ON=1'b1;
    defparam data_cntvec_i0_i2_LC_16_16_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i2_LC_16_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i2_LC_16_16_2 (
            .in0(_gnd_net_),
            .in1(N__34683),
            .in2(_gnd_net_),
            .in3(N__34661),
            .lcout(data_cntvec_2),
            .ltout(),
            .carryin(n13952),
            .carryout(n13953),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i3_LC_16_16_3.C_ON=1'b1;
    defparam data_cntvec_i0_i3_LC_16_16_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i3_LC_16_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i3_LC_16_16_3 (
            .in0(_gnd_net_),
            .in1(N__42016),
            .in2(_gnd_net_),
            .in3(N__34955),
            .lcout(data_cntvec_3),
            .ltout(),
            .carryin(n13953),
            .carryout(n13954),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i4_LC_16_16_4.C_ON=1'b1;
    defparam data_cntvec_i0_i4_LC_16_16_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i4_LC_16_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i4_LC_16_16_4 (
            .in0(_gnd_net_),
            .in1(N__37810),
            .in2(_gnd_net_),
            .in3(N__34952),
            .lcout(data_cntvec_4),
            .ltout(),
            .carryin(n13954),
            .carryout(n13955),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i5_LC_16_16_5.C_ON=1'b1;
    defparam data_cntvec_i0_i5_LC_16_16_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i5_LC_16_16_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i5_LC_16_16_5 (
            .in0(_gnd_net_),
            .in1(N__38333),
            .in2(_gnd_net_),
            .in3(N__34949),
            .lcout(data_cntvec_5),
            .ltout(),
            .carryin(n13955),
            .carryout(n13956),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i6_LC_16_16_6.C_ON=1'b1;
    defparam data_cntvec_i0_i6_LC_16_16_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i6_LC_16_16_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i6_LC_16_16_6 (
            .in0(_gnd_net_),
            .in1(N__34946),
            .in2(_gnd_net_),
            .in3(N__34928),
            .lcout(data_cntvec_6),
            .ltout(),
            .carryin(n13956),
            .carryout(n13957),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i7_LC_16_16_7.C_ON=1'b1;
    defparam data_cntvec_i0_i7_LC_16_16_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i7_LC_16_16_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i7_LC_16_16_7 (
            .in0(_gnd_net_),
            .in1(N__34920),
            .in2(_gnd_net_),
            .in3(N__34892),
            .lcout(data_cntvec_7),
            .ltout(),
            .carryin(n13957),
            .carryout(n13958),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__38048),
            .sr(N__38006));
    defparam data_cntvec_i0_i8_LC_16_17_0.C_ON=1'b1;
    defparam data_cntvec_i0_i8_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i8_LC_16_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i8_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(N__34881),
            .in2(_gnd_net_),
            .in3(N__34859),
            .lcout(data_cntvec_8),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(n13959),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_cntvec_i0_i9_LC_16_17_1.C_ON=1'b1;
    defparam data_cntvec_i0_i9_LC_16_17_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i9_LC_16_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i9_LC_16_17_1 (
            .in0(_gnd_net_),
            .in1(N__34845),
            .in2(_gnd_net_),
            .in3(N__34823),
            .lcout(data_cntvec_9),
            .ltout(),
            .carryin(n13959),
            .carryout(n13960),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_cntvec_i0_i10_LC_16_17_2.C_ON=1'b1;
    defparam data_cntvec_i0_i10_LC_16_17_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i10_LC_16_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i10_LC_16_17_2 (
            .in0(_gnd_net_),
            .in1(N__34812),
            .in2(_gnd_net_),
            .in3(N__34790),
            .lcout(data_cntvec_10),
            .ltout(),
            .carryin(n13960),
            .carryout(n13961),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_cntvec_i0_i11_LC_16_17_3.C_ON=1'b1;
    defparam data_cntvec_i0_i11_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i11_LC_16_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i11_LC_16_17_3 (
            .in0(_gnd_net_),
            .in1(N__34782),
            .in2(_gnd_net_),
            .in3(N__34763),
            .lcout(data_cntvec_11),
            .ltout(),
            .carryin(n13961),
            .carryout(n13962),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_cntvec_i0_i12_LC_16_17_4.C_ON=1'b1;
    defparam data_cntvec_i0_i12_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i12_LC_16_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i12_LC_16_17_4 (
            .in0(_gnd_net_),
            .in1(N__35470),
            .in2(_gnd_net_),
            .in3(N__35456),
            .lcout(data_cntvec_12),
            .ltout(),
            .carryin(n13962),
            .carryout(n13963),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_cntvec_i0_i13_LC_16_17_5.C_ON=1'b1;
    defparam data_cntvec_i0_i13_LC_16_17_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i13_LC_16_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i13_LC_16_17_5 (
            .in0(_gnd_net_),
            .in1(N__35446),
            .in2(_gnd_net_),
            .in3(N__35432),
            .lcout(data_cntvec_13),
            .ltout(),
            .carryin(n13963),
            .carryout(n13964),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_cntvec_i0_i14_LC_16_17_6.C_ON=1'b1;
    defparam data_cntvec_i0_i14_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i14_LC_16_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i14_LC_16_17_6 (
            .in0(_gnd_net_),
            .in1(N__35422),
            .in2(_gnd_net_),
            .in3(N__35408),
            .lcout(data_cntvec_14),
            .ltout(),
            .carryin(n13964),
            .carryout(n13965),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_cntvec_i0_i15_LC_16_17_7.C_ON=1'b0;
    defparam data_cntvec_i0_i15_LC_16_17_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i15_LC_16_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i15_LC_16_17_7 (
            .in0(_gnd_net_),
            .in1(N__35395),
            .in2(_gnd_net_),
            .in3(N__35405),
            .lcout(data_cntvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__38042),
            .sr(N__38005));
    defparam data_count_i0_i0_LC_16_18_0.C_ON=1'b1;
    defparam data_count_i0_i0_LC_16_18_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i0_LC_16_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i0_LC_16_18_0 (
            .in0(_gnd_net_),
            .in1(N__35298),
            .in2(_gnd_net_),
            .in3(N__35276),
            .lcout(data_count_0),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(n13942),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i1_LC_16_18_1.C_ON=1'b1;
    defparam data_count_i0_i1_LC_16_18_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i1_LC_16_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i1_LC_16_18_1 (
            .in0(_gnd_net_),
            .in1(N__35193),
            .in2(_gnd_net_),
            .in3(N__35171),
            .lcout(data_count_1),
            .ltout(),
            .carryin(n13942),
            .carryout(n13943),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i2_LC_16_18_2.C_ON=1'b1;
    defparam data_count_i0_i2_LC_16_18_2.SEQ_MODE=4'b1000;
    defparam data_count_i0_i2_LC_16_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i2_LC_16_18_2 (
            .in0(_gnd_net_),
            .in1(N__35088),
            .in2(_gnd_net_),
            .in3(N__35066),
            .lcout(data_count_2),
            .ltout(),
            .carryin(n13943),
            .carryout(n13944),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i3_LC_16_18_3.C_ON=1'b1;
    defparam data_count_i0_i3_LC_16_18_3.SEQ_MODE=4'b1000;
    defparam data_count_i0_i3_LC_16_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i3_LC_16_18_3 (
            .in0(_gnd_net_),
            .in1(N__34980),
            .in2(_gnd_net_),
            .in3(N__34958),
            .lcout(data_count_3),
            .ltout(),
            .carryin(n13944),
            .carryout(n13945),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i4_LC_16_18_4.C_ON=1'b1;
    defparam data_count_i0_i4_LC_16_18_4.SEQ_MODE=4'b1000;
    defparam data_count_i0_i4_LC_16_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i4_LC_16_18_4 (
            .in0(_gnd_net_),
            .in1(N__36216),
            .in2(_gnd_net_),
            .in3(N__36194),
            .lcout(data_count_4),
            .ltout(),
            .carryin(n13945),
            .carryout(n13946),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i5_LC_16_18_5.C_ON=1'b1;
    defparam data_count_i0_i5_LC_16_18_5.SEQ_MODE=4'b1000;
    defparam data_count_i0_i5_LC_16_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i5_LC_16_18_5 (
            .in0(_gnd_net_),
            .in1(N__36108),
            .in2(_gnd_net_),
            .in3(N__36086),
            .lcout(data_count_5),
            .ltout(),
            .carryin(n13946),
            .carryout(n13947),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i6_LC_16_18_6.C_ON=1'b1;
    defparam data_count_i0_i6_LC_16_18_6.SEQ_MODE=4'b1000;
    defparam data_count_i0_i6_LC_16_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i6_LC_16_18_6 (
            .in0(_gnd_net_),
            .in1(N__36000),
            .in2(_gnd_net_),
            .in3(N__35978),
            .lcout(data_count_6),
            .ltout(),
            .carryin(n13947),
            .carryout(n13948),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i7_LC_16_18_7.C_ON=1'b1;
    defparam data_count_i0_i7_LC_16_18_7.SEQ_MODE=4'b1000;
    defparam data_count_i0_i7_LC_16_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i7_LC_16_18_7 (
            .in0(_gnd_net_),
            .in1(N__35895),
            .in2(_gnd_net_),
            .in3(N__35873),
            .lcout(data_count_7),
            .ltout(),
            .carryin(n13948),
            .carryout(n13949),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__38041),
            .sr(N__37995));
    defparam data_count_i0_i8_LC_16_19_0.C_ON=1'b0;
    defparam data_count_i0_i8_LC_16_19_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i8_LC_16_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i8_LC_16_19_0 (
            .in0(_gnd_net_),
            .in1(N__35787),
            .in2(_gnd_net_),
            .in3(N__35870),
            .lcout(data_count_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__38043),
            .sr(N__37994));
    defparam \CLOCK_DDS.dds_state_i1_LC_17_4_0 .C_ON=1'b0;
    defparam \CLOCK_DDS.dds_state_i1_LC_17_4_0 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.dds_state_i1_LC_17_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLOCK_DDS.dds_state_i1_LC_17_4_0  (
            .in0(_gnd_net_),
            .in1(N__35670),
            .in2(_gnd_net_),
            .in3(N__48380),
            .lcout(dds_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51124),
            .ce(N__48299),
            .sr(N__48538));
    defparam \comm_spi.data_rx_i0_7344_7345_set_LC_17_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_7344_7345_set_LC_17_5_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_rx_i0_7344_7345_set_LC_17_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_7344_7345_set_LC_17_5_0  (
            .in0(N__42236),
            .in1(N__45818),
            .in2(_gnd_net_),
            .in3(N__42260),
            .lcout(\comm_spi.n10455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42371),
            .ce(),
            .sr(N__42203));
    defparam \ADC_VAC2.i1_3_lut_LC_17_6_0 .C_ON=1'b0;
    defparam \ADC_VAC2.i1_3_lut_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i1_3_lut_LC_17_6_0 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \ADC_VAC2.i1_3_lut_LC_17_6_0  (
            .in0(N__53482),
            .in1(N__35539),
            .in2(_gnd_net_),
            .in3(N__35636),
            .lcout(\ADC_VAC2.n14926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.adc_state_i1_LC_17_6_1 .C_ON=1'b0;
    defparam \ADC_VAC2.adc_state_i1_LC_17_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.adc_state_i1_LC_17_6_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_VAC2.adc_state_i1_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__36485),
            .in2(_gnd_net_),
            .in3(N__53483),
            .lcout(adc_state_1_adj_1043),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51145),
            .ce(N__35510),
            .sr(N__36521));
    defparam \ADC_VAC2.i7600_2_lut_LC_17_6_3 .C_ON=1'b0;
    defparam \ADC_VAC2.i7600_2_lut_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC2.i7600_2_lut_LC_17_6_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ADC_VAC2.i7600_2_lut_LC_17_6_3  (
            .in0(N__36509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36484),
            .lcout(\ADC_VAC2.n10706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i7328_3_lut_LC_17_6_5 .C_ON=1'b0;
    defparam \comm_spi.i7328_3_lut_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i7328_3_lut_LC_17_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.i7328_3_lut_LC_17_6_5  (
            .in0(N__38465),
            .in1(N__37967),
            .in2(_gnd_net_),
            .in3(N__51335),
            .lcout(\comm_spi.iclk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i2_3_lut_LC_17_6_6 .C_ON=1'b0;
    defparam \comm_spi.i2_3_lut_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i2_3_lut_LC_17_6_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \comm_spi.i2_3_lut_LC_17_6_6  (
            .in0(N__36341),
            .in1(N__36357),
            .in2(_gnd_net_),
            .in3(N__36319),
            .lcout(\comm_spi.n12175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.bit_cnt_1603__i3_LC_17_7_0 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_1603__i3_LC_17_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_1603__i3_LC_17_7_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \comm_spi.bit_cnt_1603__i3_LC_17_7_0  (
            .in0(N__36359),
            .in1(N__38419),
            .in2(N__36326),
            .in3(N__36344),
            .lcout(\comm_spi.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_1603__i3C_net ),
            .ce(),
            .sr(N__46584));
    defparam \comm_spi.bit_cnt_1603__i2_LC_17_7_1 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_1603__i2_LC_17_7_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_1603__i2_LC_17_7_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \comm_spi.bit_cnt_1603__i2_LC_17_7_1  (
            .in0(N__36343),
            .in1(N__36322),
            .in2(_gnd_net_),
            .in3(N__36358),
            .lcout(\comm_spi.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_1603__i3C_net ),
            .ce(),
            .sr(N__46584));
    defparam \comm_spi.bit_cnt_1603__i1_LC_17_7_2 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_1603__i1_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_1603__i1_LC_17_7_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \comm_spi.bit_cnt_1603__i1_LC_17_7_2  (
            .in0(N__36321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36342),
            .lcout(\comm_spi.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_1603__i3C_net ),
            .ce(),
            .sr(N__46584));
    defparam \comm_spi.bit_cnt_1603__i0_LC_17_7_3 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_1603__i0_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_1603__i0_LC_17_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \comm_spi.bit_cnt_1603__i0_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36320),
            .lcout(\comm_spi.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_1603__i3C_net ),
            .ce(),
            .sr(N__46584));
    defparam i12087_2_lut_3_lut_LC_17_7_4.C_ON=1'b0;
    defparam i12087_2_lut_3_lut_LC_17_7_4.SEQ_MODE=4'b0000;
    defparam i12087_2_lut_3_lut_LC_17_7_4.LUT_INIT=16'b0100010000000000;
    LogicCell40 i12087_2_lut_3_lut_LC_17_7_4 (
            .in0(N__43445),
            .in1(N__50501),
            .in2(_gnd_net_),
            .in3(N__43267),
            .lcout(n15290),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_282_LC_17_7_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_282_LC_17_7_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_282_LC_17_7_5.LUT_INIT=16'b1101110111111111;
    LogicCell40 i1_2_lut_3_lut_adj_282_LC_17_7_5 (
            .in0(N__43268),
            .in1(N__43447),
            .in2(_gnd_net_),
            .in3(N__50499),
            .lcout(n4_adj_1179),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_175_LC_17_7_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_175_LC_17_7_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_175_LC_17_7_6.LUT_INIT=16'b0011001110111011;
    LogicCell40 i1_2_lut_3_lut_adj_175_LC_17_7_6 (
            .in0(N__43446),
            .in1(N__50500),
            .in2(_gnd_net_),
            .in3(N__43265),
            .lcout(n15198),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_3_lut_LC_17_7_7.C_ON=1'b0;
    defparam i3_2_lut_3_lut_LC_17_7_7.SEQ_MODE=4'b0000;
    defparam i3_2_lut_3_lut_LC_17_7_7.LUT_INIT=16'b1111111111101110;
    LogicCell40 i3_2_lut_3_lut_LC_17_7_7 (
            .in0(N__43266),
            .in1(N__43448),
            .in2(_gnd_net_),
            .in3(N__50498),
            .lcout(n8530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_378_Mux_1_i8_3_lut_4_lut_LC_17_8_0.C_ON=1'b0;
    defparam comm_state_3__I_0_378_Mux_1_i8_3_lut_4_lut_LC_17_8_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_378_Mux_1_i8_3_lut_4_lut_LC_17_8_0.LUT_INIT=16'b0000010110001101;
    LogicCell40 comm_state_3__I_0_378_Mux_1_i8_3_lut_4_lut_LC_17_8_0 (
            .in0(N__50510),
            .in1(N__49774),
            .in2(N__39443),
            .in3(N__36548),
            .lcout(n8_adj_1201),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12842_2_lut_LC_17_8_1.C_ON=1'b0;
    defparam i12842_2_lut_LC_17_8_1.SEQ_MODE=4'b0000;
    defparam i12842_2_lut_LC_17_8_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 i12842_2_lut_LC_17_8_1 (
            .in0(_gnd_net_),
            .in1(N__50509),
            .in2(_gnd_net_),
            .in3(N__42706),
            .lcout(),
            .ltout(n15668_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_1__bdd_4_lut_LC_17_8_2.C_ON=1'b0;
    defparam comm_state_1__bdd_4_lut_LC_17_8_2.SEQ_MODE=4'b0000;
    defparam comm_state_1__bdd_4_lut_LC_17_8_2.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_state_1__bdd_4_lut_LC_17_8_2 (
            .in0(N__39040),
            .in1(N__49773),
            .in2(N__36551),
            .in3(N__49480),
            .lcout(n16464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i244_2_lut_LC_17_8_3.C_ON=1'b0;
    defparam i244_2_lut_LC_17_8_3.SEQ_MODE=4'b0000;
    defparam i244_2_lut_LC_17_8_3.LUT_INIT=16'b0101000001010000;
    LogicCell40 i244_2_lut_LC_17_8_3 (
            .in0(N__43287),
            .in1(_gnd_net_),
            .in2(N__43438),
            .in3(_gnd_net_),
            .lcout(n1523),
            .ltout(n1523_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_378_Mux_1_i2_3_lut_4_lut_LC_17_8_4.C_ON=1'b0;
    defparam comm_state_3__I_0_378_Mux_1_i2_3_lut_4_lut_LC_17_8_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_378_Mux_1_i2_3_lut_4_lut_LC_17_8_4.LUT_INIT=16'b0100111001000100;
    LogicCell40 comm_state_3__I_0_378_Mux_1_i2_3_lut_4_lut_LC_17_8_4 (
            .in0(N__50511),
            .in1(N__43406),
            .in2(N__36542),
            .in3(N__49775),
            .lcout(),
            .ltout(n2_adj_1200_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n16464_bdd_4_lut_LC_17_8_5.C_ON=1'b0;
    defparam n16464_bdd_4_lut_LC_17_8_5.SEQ_MODE=4'b0000;
    defparam n16464_bdd_4_lut_LC_17_8_5.LUT_INIT=16'b1111101001000100;
    LogicCell40 n16464_bdd_4_lut_LC_17_8_5 (
            .in0(N__49481),
            .in1(N__50512),
            .in2(N__36539),
            .in3(N__36536),
            .lcout(),
            .ltout(n16467_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i1_LC_17_8_6.C_ON=1'b0;
    defparam comm_state_i1_LC_17_8_6.SEQ_MODE=4'b1000;
    defparam comm_state_i1_LC_17_8_6.LUT_INIT=16'b0111010000110000;
    LogicCell40 comm_state_i1_LC_17_8_6 (
            .in0(N__51927),
            .in1(N__52066),
            .in2(N__36530),
            .in3(N__36527),
            .lcout(comm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51170),
            .ce(N__36620),
            .sr(_gnd_net_));
    defparam i13037_4_lut_LC_17_8_7.C_ON=1'b0;
    defparam i13037_4_lut_LC_17_8_7.SEQ_MODE=4'b0000;
    defparam i13037_4_lut_LC_17_8_7.LUT_INIT=16'b1111010011110111;
    LogicCell40 i13037_4_lut_LC_17_8_7 (
            .in0(N__36629),
            .in1(N__50508),
            .in2(N__52165),
            .in3(N__36557),
            .lcout(n14_adj_1189),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_407_i13_2_lut_3_lut_4_lut_LC_17_9_0.C_ON=1'b0;
    defparam comm_cmd_6__I_0_407_i13_2_lut_3_lut_4_lut_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_407_i13_2_lut_3_lut_4_lut_LC_17_9_0.LUT_INIT=16'b1111111111111101;
    LogicCell40 comm_cmd_6__I_0_407_i13_2_lut_3_lut_4_lut_LC_17_9_0 (
            .in0(N__47509),
            .in1(N__45415),
            .in2(N__39013),
            .in3(N__45224),
            .lcout(n13_adj_1032),
            .ltout(n13_adj_1032_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_249_LC_17_9_1.C_ON=1'b0;
    defparam i1_3_lut_adj_249_LC_17_9_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_249_LC_17_9_1.LUT_INIT=16'b1100110011001111;
    LogicCell40 i1_3_lut_adj_249_LC_17_9_1 (
            .in0(_gnd_net_),
            .in1(N__43165),
            .in2(N__36599),
            .in3(N__50502),
            .lcout(n8519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_246_LC_17_9_2.C_ON=1'b0;
    defparam i1_2_lut_adj_246_LC_17_9_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_246_LC_17_9_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_246_LC_17_9_2 (
            .in0(_gnd_net_),
            .in1(N__47048),
            .in2(_gnd_net_),
            .in3(N__40862),
            .lcout(n12_adj_1027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_63_LC_17_9_3.C_ON=1'b0;
    defparam i1_4_lut_adj_63_LC_17_9_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_63_LC_17_9_3.LUT_INIT=16'b1010111010101010;
    LogicCell40 i1_4_lut_adj_63_LC_17_9_3 (
            .in0(N__40863),
            .in1(N__47508),
            .in2(N__47183),
            .in3(N__45454),
            .lcout(n22_adj_1115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i3_LC_17_9_4.C_ON=1'b0;
    defparam buf_dds_i3_LC_17_9_4.SEQ_MODE=4'b1000;
    defparam buf_dds_i3_LC_17_9_4.LUT_INIT=16'b1110001011101110;
    LogicCell40 buf_dds_i3_LC_17_9_4 (
            .in0(N__40965),
            .in1(N__41314),
            .in2(N__43916),
            .in3(N__52302),
            .lcout(buf_dds_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51188),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_296_LC_17_9_5.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_296_LC_17_9_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_296_LC_17_9_5.LUT_INIT=16'b1111111010101010;
    LogicCell40 i1_4_lut_4_lut_adj_296_LC_17_9_5 (
            .in0(N__40861),
            .in1(N__44967),
            .in2(N__47184),
            .in3(N__43188),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12836_2_lut_3_lut_LC_17_9_6.C_ON=1'b0;
    defparam i12836_2_lut_3_lut_LC_17_9_6.SEQ_MODE=4'b0000;
    defparam i12836_2_lut_3_lut_LC_17_9_6.LUT_INIT=16'b0100010000000000;
    LogicCell40 i12836_2_lut_3_lut_LC_17_9_6 (
            .in0(N__47507),
            .in1(N__45414),
            .in2(_gnd_net_),
            .in3(N__45223),
            .lcout(n15651),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12628_3_lut_LC_17_9_7.C_ON=1'b0;
    defparam i12628_3_lut_LC_17_9_7.SEQ_MODE=4'b0000;
    defparam i12628_3_lut_LC_17_9_7.LUT_INIT=16'b0001000100000000;
    LogicCell40 i12628_3_lut_LC_17_9_7 (
            .in0(N__43449),
            .in1(N__43289),
            .in2(_gnd_net_),
            .in3(N__49741),
            .lcout(n15526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12680_4_lut_4_lut_LC_17_10_0.C_ON=1'b0;
    defparam i12680_4_lut_4_lut_LC_17_10_0.SEQ_MODE=4'b0000;
    defparam i12680_4_lut_4_lut_LC_17_10_0.LUT_INIT=16'b1101100001010000;
    LogicCell40 i12680_4_lut_4_lut_LC_17_10_0 (
            .in0(N__46908),
            .in1(N__40196),
            .in2(N__36972),
            .in3(N__37687),
            .lcout(n15584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_115_LC_17_10_1.C_ON=1'b0;
    defparam i1_4_lut_adj_115_LC_17_10_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_115_LC_17_10_1.LUT_INIT=16'b1010100000000000;
    LogicCell40 i1_4_lut_adj_115_LC_17_10_1 (
            .in0(N__40195),
            .in1(N__47594),
            .in2(N__37016),
            .in3(N__46909),
            .lcout(),
            .ltout(n8058_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_271_LC_17_10_2.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_271_LC_17_10_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_271_LC_17_10_2.LUT_INIT=16'b1010001010100000;
    LogicCell40 i1_3_lut_4_lut_adj_271_LC_17_10_2 (
            .in0(N__45279),
            .in1(N__46911),
            .in2(N__36998),
            .in3(N__36973),
            .lcout(),
            .ltout(n83_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12771_4_lut_LC_17_10_3.C_ON=1'b0;
    defparam i12771_4_lut_LC_17_10_3.SEQ_MODE=4'b0000;
    defparam i12771_4_lut_LC_17_10_3.LUT_INIT=16'b1010100010100000;
    LogicCell40 i12771_4_lut_LC_17_10_3 (
            .in0(N__45537),
            .in1(N__36896),
            .in2(N__36890),
            .in3(N__47595),
            .lcout(n15581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i21_LC_17_10_4 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i21_LC_17_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i21_LC_17_10_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i21_LC_17_10_4  (
            .in0(N__44404),
            .in1(N__49268),
            .in2(N__36844),
            .in3(N__36877),
            .lcout(buf_adcdata3_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51206),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_301_LC_17_10_5.C_ON=1'b0;
    defparam i1_4_lut_adj_301_LC_17_10_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_301_LC_17_10_5.LUT_INIT=16'b1101000011000000;
    LogicCell40 i1_4_lut_adj_301_LC_17_10_5 (
            .in0(N__45536),
            .in1(N__39410),
            .in2(N__40224),
            .in3(N__40753),
            .lcout(comm_state_3_N_402_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i15_LC_17_10_6 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i15_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i15_LC_17_10_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i15_LC_17_10_6  (
            .in0(N__44403),
            .in1(N__49267),
            .in2(N__36806),
            .in3(N__36762),
            .lcout(buf_adcdata3_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51206),
            .ce(),
            .sr(_gnd_net_));
    defparam i129_4_lut_LC_17_10_7.C_ON=1'b0;
    defparam i129_4_lut_LC_17_10_7.SEQ_MODE=4'b0000;
    defparam i129_4_lut_LC_17_10_7.LUT_INIT=16'b0010001011000000;
    LogicCell40 i129_4_lut_LC_17_10_7 (
            .in0(N__36743),
            .in1(N__47593),
            .in2(N__37169),
            .in3(N__45278),
            .lcout(n75_adj_1164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_idxvec_i0_LC_17_11_0.C_ON=1'b0;
    defparam data_idxvec_i0_LC_17_11_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i0_LC_17_11_0.LUT_INIT=16'b0011000010101010;
    LogicCell40 data_idxvec_i0_LC_17_11_0 (
            .in0(N__37049),
            .in1(N__51893),
            .in2(N__36705),
            .in3(N__52301),
            .lcout(data_idxvec_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51223),
            .ce(N__37556),
            .sr(_gnd_net_));
    defparam mux_1494_i1_3_lut_LC_17_11_1.C_ON=1'b0;
    defparam mux_1494_i1_3_lut_LC_17_11_1.SEQ_MODE=4'b0000;
    defparam mux_1494_i1_3_lut_LC_17_11_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_1494_i1_3_lut_LC_17_11_1 (
            .in0(N__37060),
            .in1(N__47540),
            .in2(_gnd_net_),
            .in3(N__36653),
            .lcout(),
            .ltout(n4197_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i1_4_lut_LC_17_11_2.C_ON=1'b0;
    defparam mux_1507_i1_4_lut_LC_17_11_2.SEQ_MODE=4'b0000;
    defparam mux_1507_i1_4_lut_LC_17_11_2.LUT_INIT=16'b0100010011110000;
    LogicCell40 mux_1507_i1_4_lut_LC_17_11_2 (
            .in0(N__47541),
            .in1(N__37145),
            .in2(N__37127),
            .in3(N__45183),
            .lcout(),
            .ltout(n4234_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i1_3_lut_LC_17_11_3.C_ON=1'b0;
    defparam mux_1511_i1_3_lut_LC_17_11_3.SEQ_MODE=4'b0000;
    defparam mux_1511_i1_3_lut_LC_17_11_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_1511_i1_3_lut_LC_17_11_3 (
            .in0(_gnd_net_),
            .in1(N__37124),
            .in2(N__37112),
            .in3(N__45436),
            .lcout(),
            .ltout(n4254_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1513_i1_4_lut_LC_17_11_4.C_ON=1'b0;
    defparam mux_1513_i1_4_lut_LC_17_11_4.SEQ_MODE=4'b0000;
    defparam mux_1513_i1_4_lut_LC_17_11_4.LUT_INIT=16'b1111000000100010;
    LogicCell40 mux_1513_i1_4_lut_LC_17_11_4 (
            .in0(N__37109),
            .in1(N__45184),
            .in2(N__37091),
            .in3(N__46835),
            .lcout(n4264),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i37_4_lut_4_lut_LC_17_11_6.C_ON=1'b0;
    defparam i37_4_lut_4_lut_LC_17_11_6.SEQ_MODE=4'b0000;
    defparam i37_4_lut_4_lut_LC_17_11_6.LUT_INIT=16'b1001001001010010;
    LogicCell40 i37_4_lut_4_lut_LC_17_11_6 (
            .in0(N__45435),
            .in1(N__45182),
            .in2(N__47670),
            .in3(N__46833),
            .lcout(),
            .ltout(n32_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12654_4_lut_LC_17_11_7.C_ON=1'b0;
    defparam i12654_4_lut_LC_17_11_7.SEQ_MODE=4'b0000;
    defparam i12654_4_lut_LC_17_11_7.LUT_INIT=16'b1111100000000000;
    LogicCell40 i12654_4_lut_LC_17_11_7 (
            .in0(N__46834),
            .in1(N__40754),
            .in2(N__37082),
            .in3(N__40164),
            .lcout(n15557),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_1441_2_lut_LC_17_12_0.C_ON=1'b1;
    defparam add_1441_2_lut_LC_17_12_0.SEQ_MODE=4'b0000;
    defparam add_1441_2_lut_LC_17_12_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_1441_2_lut_LC_17_12_0 (
            .in0(_gnd_net_),
            .in1(N__43615),
            .in2(N__37064),
            .in3(_gnd_net_),
            .lcout(data_idxvec_15_N_673_0),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(n14040),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_idxvec_i1_LC_17_12_1.C_ON=1'b1;
    defparam data_idxvec_i1_LC_17_12_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i1_LC_17_12_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i1_LC_17_12_1 (
            .in0(N__37492),
            .in1(N__38242),
            .in2(N__52456),
            .in3(N__37043),
            .lcout(data_idxvec_1),
            .ltout(),
            .carryin(n14040),
            .carryout(n14041),
            .clk(N__51240),
            .ce(N__37552),
            .sr(_gnd_net_));
    defparam data_idxvec_i2_LC_17_12_2.C_ON=1'b1;
    defparam data_idxvec_i2_LC_17_12_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i2_LC_17_12_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i2_LC_17_12_2 (
            .in0(N__40345),
            .in1(N__52394),
            .in2(N__37040),
            .in3(N__37019),
            .lcout(data_idxvec_2),
            .ltout(),
            .carryin(n14041),
            .carryout(n14042),
            .clk(N__51240),
            .ce(N__37552),
            .sr(_gnd_net_));
    defparam data_idxvec_i3_LC_17_12_3.C_ON=1'b1;
    defparam data_idxvec_i3_LC_17_12_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i3_LC_17_12_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i3_LC_17_12_3 (
            .in0(N__43909),
            .in1(N__42031),
            .in2(N__52457),
            .in3(N__37403),
            .lcout(data_idxvec_3),
            .ltout(),
            .carryin(n14042),
            .carryout(n14043),
            .clk(N__51240),
            .ce(N__37552),
            .sr(_gnd_net_));
    defparam data_idxvec_i4_LC_17_12_4.C_ON=1'b1;
    defparam data_idxvec_i4_LC_17_12_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i4_LC_17_12_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i4_LC_17_12_4 (
            .in0(N__37399),
            .in1(N__52398),
            .in2(N__37829),
            .in3(N__37376),
            .lcout(data_idxvec_4),
            .ltout(),
            .carryin(n14043),
            .carryout(n14044),
            .clk(N__51240),
            .ce(N__37552),
            .sr(_gnd_net_));
    defparam data_idxvec_i5_LC_17_12_5.C_ON=1'b1;
    defparam data_idxvec_i5_LC_17_12_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i5_LC_17_12_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i5_LC_17_12_5 (
            .in0(N__37373),
            .in1(N__38347),
            .in2(N__52458),
            .in3(N__37349),
            .lcout(data_idxvec_5),
            .ltout(),
            .carryin(n14044),
            .carryout(n14045),
            .clk(N__51240),
            .ce(N__37552),
            .sr(_gnd_net_));
    defparam data_idxvec_i6_LC_17_12_6.C_ON=1'b1;
    defparam data_idxvec_i6_LC_17_12_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i6_LC_17_12_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i6_LC_17_12_6 (
            .in0(N__37945),
            .in1(N__52402),
            .in2(N__37345),
            .in3(N__37325),
            .lcout(data_idxvec_6),
            .ltout(),
            .carryin(n14045),
            .carryout(n14046),
            .clk(N__51240),
            .ce(N__37552),
            .sr(_gnd_net_));
    defparam data_idxvec_i7_LC_17_12_7.C_ON=1'b1;
    defparam data_idxvec_i7_LC_17_12_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i7_LC_17_12_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i7_LC_17_12_7 (
            .in0(N__37322),
            .in1(N__37294),
            .in2(N__52459),
            .in3(N__37280),
            .lcout(data_idxvec_7),
            .ltout(),
            .carryin(n14046),
            .carryout(n14047),
            .clk(N__51240),
            .ce(N__37552),
            .sr(_gnd_net_));
    defparam data_idxvec_i8_LC_17_13_0.C_ON=1'b1;
    defparam data_idxvec_i8_LC_17_13_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i8_LC_17_13_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i8_LC_17_13_0 (
            .in0(N__37277),
            .in1(N__52406),
            .in2(N__41003),
            .in3(N__37241),
            .lcout(data_idxvec_8),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(n14048),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam data_idxvec_i9_LC_17_13_1.C_ON=1'b1;
    defparam data_idxvec_i9_LC_17_13_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i9_LC_17_13_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i9_LC_17_13_1 (
            .in0(N__37237),
            .in1(N__37207),
            .in2(N__52460),
            .in3(N__37193),
            .lcout(data_idxvec_9),
            .ltout(),
            .carryin(n14048),
            .carryout(n14049),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam data_idxvec_i10_LC_17_13_2.C_ON=1'b1;
    defparam data_idxvec_i10_LC_17_13_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i10_LC_17_13_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i10_LC_17_13_2 (
            .in0(N__37189),
            .in1(N__52410),
            .in2(N__37168),
            .in3(N__37148),
            .lcout(data_idxvec_10),
            .ltout(),
            .carryin(n14049),
            .carryout(n14050),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam data_idxvec_i11_LC_17_13_3.C_ON=1'b1;
    defparam data_idxvec_i11_LC_17_13_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i11_LC_17_13_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i11_LC_17_13_3 (
            .in0(N__43492),
            .in1(N__40579),
            .in2(N__52461),
            .in3(N__37721),
            .lcout(data_idxvec_11),
            .ltout(),
            .carryin(n14050),
            .carryout(n14051),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam data_idxvec_i12_LC_17_13_4.C_ON=1'b1;
    defparam data_idxvec_i12_LC_17_13_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i12_LC_17_13_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i12_LC_17_13_4 (
            .in0(N__37711),
            .in1(N__52414),
            .in2(N__37688),
            .in3(N__37670),
            .lcout(data_idxvec_12),
            .ltout(),
            .carryin(n14051),
            .carryout(n14052),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam data_idxvec_i13_LC_17_13_5.C_ON=1'b1;
    defparam data_idxvec_i13_LC_17_13_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i13_LC_17_13_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i13_LC_17_13_5 (
            .in0(N__37667),
            .in1(N__37648),
            .in2(N__52462),
            .in3(N__37634),
            .lcout(data_idxvec_13),
            .ltout(),
            .carryin(n14052),
            .carryout(n14053),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam data_idxvec_i14_LC_17_13_6.C_ON=1'b1;
    defparam data_idxvec_i14_LC_17_13_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i14_LC_17_13_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i14_LC_17_13_6 (
            .in0(N__37631),
            .in1(N__52418),
            .in2(N__37606),
            .in3(N__37586),
            .lcout(data_idxvec_14),
            .ltout(),
            .carryin(n14053),
            .carryout(n14054),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam data_idxvec_i15_LC_17_13_7.C_ON=1'b0;
    defparam data_idxvec_i15_LC_17_13_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i15_LC_17_13_7.LUT_INIT=16'b1000110111011000;
    LogicCell40 data_idxvec_i15_LC_17_13_7 (
            .in0(N__52419),
            .in1(N__37582),
            .in2(N__41675),
            .in3(N__37559),
            .lcout(data_idxvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51255),
            .ce(N__37545),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i13_LC_17_14_1 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i13_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i13_LC_17_14_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i13_LC_17_14_1  (
            .in0(N__49077),
            .in1(N__44398),
            .in2(N__41957),
            .in3(N__37516),
            .lcout(buf_adcdata3_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51272),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i1_LC_17_14_2.C_ON=1'b0;
    defparam req_data_cnt_i1_LC_17_14_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i1_LC_17_14_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i1_LC_17_14_2 (
            .in0(N__37496),
            .in1(N__40462),
            .in2(_gnd_net_),
            .in3(N__42161),
            .lcout(req_data_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51272),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i14_LC_17_14_3 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i14_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i14_LC_17_14_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i14_LC_17_14_3  (
            .in0(N__53115),
            .in1(N__37441),
            .in2(N__37475),
            .in3(N__52794),
            .lcout(buf_adcdata1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51272),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i11_LC_17_14_4.C_ON=1'b0;
    defparam req_data_cnt_i11_LC_17_14_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i11_LC_17_14_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i11_LC_17_14_4 (
            .in0(N__43493),
            .in1(N__40461),
            .in2(_gnd_net_),
            .in3(N__37422),
            .lcout(req_data_cnt_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51272),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i22_LC_17_14_5 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i22_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i22_LC_17_14_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i22_LC_17_14_5  (
            .in0(N__49078),
            .in1(N__41574),
            .in2(N__41956),
            .in3(N__48810),
            .lcout(cmd_rdadctmp_22_adj_1090),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51272),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i6_LC_17_14_6.C_ON=1'b0;
    defparam req_data_cnt_i6_LC_17_14_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i6_LC_17_14_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i6_LC_17_14_6 (
            .in0(N__37949),
            .in1(N__40463),
            .in2(_gnd_net_),
            .in3(N__37917),
            .lcout(req_data_cnt_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51272),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i15_LC_17_14_7.C_ON=1'b0;
    defparam acadc_skipCount_i15_LC_17_14_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i15_LC_17_14_7.LUT_INIT=16'b0011000010111000;
    LogicCell40 acadc_skipCount_i15_LC_17_14_7 (
            .in0(N__38923),
            .in1(N__41757),
            .in2(N__41657),
            .in3(N__51896),
            .lcout(acadc_skipCount_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51272),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i6_3_lut_LC_17_15_0.C_ON=1'b0;
    defparam mux_1511_i6_3_lut_LC_17_15_0.SEQ_MODE=4'b0000;
    defparam mux_1511_i6_3_lut_LC_17_15_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_1511_i6_3_lut_LC_17_15_0 (
            .in0(N__37727),
            .in1(N__45602),
            .in2(_gnd_net_),
            .in3(N__38300),
            .lcout(),
            .ltout(n4249_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1513_i6_4_lut_LC_17_15_1.C_ON=1'b0;
    defparam mux_1513_i6_4_lut_LC_17_15_1.SEQ_MODE=4'b0000;
    defparam mux_1513_i6_4_lut_LC_17_15_1.LUT_INIT=16'b1111000001000100;
    LogicCell40 mux_1513_i6_4_lut_LC_17_15_1 (
            .in0(N__45263),
            .in1(N__37901),
            .in2(N__37889),
            .in3(N__47266),
            .lcout(),
            .ltout(n4259_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i5_LC_17_15_2.C_ON=1'b0;
    defparam comm_buf_1__i5_LC_17_15_2.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i5_LC_17_15_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i5_LC_17_15_2 (
            .in0(N__39765),
            .in1(_gnd_net_),
            .in2(N__37886),
            .in3(N__50289),
            .lcout(comm_buf_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51284),
            .ce(N__44717),
            .sr(N__44652));
    defparam mux_1494_i5_3_lut_LC_17_15_3.C_ON=1'b0;
    defparam mux_1494_i5_3_lut_LC_17_15_3.SEQ_MODE=4'b0000;
    defparam mux_1494_i5_3_lut_LC_17_15_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_1494_i5_3_lut_LC_17_15_3 (
            .in0(N__37828),
            .in1(N__47792),
            .in2(_gnd_net_),
            .in3(N__37806),
            .lcout(),
            .ltout(n4193_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i5_4_lut_LC_17_15_4.C_ON=1'b0;
    defparam mux_1507_i5_4_lut_LC_17_15_4.SEQ_MODE=4'b0000;
    defparam mux_1507_i5_4_lut_LC_17_15_4.LUT_INIT=16'b0010001011110000;
    LogicCell40 mux_1507_i5_4_lut_LC_17_15_4 (
            .in0(N__37790),
            .in1(N__47798),
            .in2(N__37775),
            .in3(N__45261),
            .lcout(n4230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i6_3_lut_LC_17_15_5.C_ON=1'b0;
    defparam mux_1502_i6_3_lut_LC_17_15_5.SEQ_MODE=4'b0000;
    defparam mux_1502_i6_3_lut_LC_17_15_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_1502_i6_3_lut_LC_17_15_5 (
            .in0(N__47799),
            .in1(N__37767),
            .in2(_gnd_net_),
            .in3(N__37748),
            .lcout(n4216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1494_i6_3_lut_LC_17_15_6.C_ON=1'b0;
    defparam mux_1494_i6_3_lut_LC_17_15_6.SEQ_MODE=4'b0000;
    defparam mux_1494_i6_3_lut_LC_17_15_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_1494_i6_3_lut_LC_17_15_6 (
            .in0(N__47793),
            .in1(N__38348),
            .in2(_gnd_net_),
            .in3(N__38331),
            .lcout(),
            .ltout(n4192_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i6_4_lut_LC_17_15_7.C_ON=1'b0;
    defparam mux_1507_i6_4_lut_LC_17_15_7.SEQ_MODE=4'b0000;
    defparam mux_1507_i6_4_lut_LC_17_15_7.LUT_INIT=16'b1111101011011000;
    LogicCell40 mux_1507_i6_4_lut_LC_17_15_7 (
            .in0(N__45262),
            .in1(N__38315),
            .in2(N__38303),
            .in3(N__47794),
            .lcout(n4229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i10_LC_17_16_0 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i10_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i10_LC_17_16_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i10_LC_17_16_0  (
            .in0(N__53752),
            .in1(N__38257),
            .in2(N__38294),
            .in3(N__53493),
            .lcout(buf_adcdata2_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51295),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1494_i2_3_lut_LC_17_16_2.C_ON=1'b0;
    defparam mux_1494_i2_3_lut_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam mux_1494_i2_3_lut_LC_17_16_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_1494_i2_3_lut_LC_17_16_2 (
            .in0(N__38243),
            .in1(N__38223),
            .in2(_gnd_net_),
            .in3(N__47791),
            .lcout(n4196),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i17_LC_17_16_4 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i17_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i17_LC_17_16_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i17_LC_17_16_4  (
            .in0(N__38200),
            .in1(N__49212),
            .in2(N__44535),
            .in3(N__48809),
            .lcout(cmd_rdadctmp_17_adj_1095),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51295),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i4_3_lut_LC_17_17_4.C_ON=1'b0;
    defparam mux_1502_i4_3_lut_LC_17_17_4.SEQ_MODE=4'b0000;
    defparam mux_1502_i4_3_lut_LC_17_17_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_1502_i4_3_lut_LC_17_17_4 (
            .in0(N__47928),
            .in1(N__38174),
            .in2(_gnd_net_),
            .in3(N__38150),
            .lcout(n4218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7374_2_lut_LC_17_19_5.C_ON=1'b0;
    defparam i7374_2_lut_LC_17_19_5.SEQ_MODE=4'b0000;
    defparam i7374_2_lut_LC_17_19_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i7374_2_lut_LC_17_19_5 (
            .in0(_gnd_net_),
            .in1(N__38131),
            .in2(_gnd_net_),
            .in3(N__38047),
            .lcout(n10483),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13067_4_lut_3_lut_LC_18_3_1 .C_ON=1'b0;
    defparam \comm_spi.i13067_4_lut_3_lut_LC_18_3_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13067_4_lut_3_lut_LC_18_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i13067_4_lut_3_lut_LC_18_3_1  (
            .in0(N__46560),
            .in1(N__51390),
            .in2(_gnd_net_),
            .in3(N__37960),
            .lcout(\comm_spi.n16887 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_7326_7327_reset_LC_18_4_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_7326_7327_reset_LC_18_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.iclk_40_7326_7327_reset_LC_18_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.iclk_40_7326_7327_reset_LC_18_4_0  (
            .in0(N__51397),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n10438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51133),
            .ce(),
            .sr(N__38453));
    defparam \comm_spi.i13087_4_lut_3_lut_LC_18_5_4 .C_ON=1'b0;
    defparam \comm_spi.i13087_4_lut_3_lut_LC_18_5_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13087_4_lut_3_lut_LC_18_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i13087_4_lut_3_lut_LC_18_5_4  (
            .in0(N__46503),
            .in1(N__42889),
            .in2(_gnd_net_),
            .in3(N__38438),
            .lcout(\comm_spi.n16890 ),
            .ltout(\comm_spi.n16890_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i7346_3_lut_LC_18_5_5 .C_ON=1'b0;
    defparam \comm_spi.i7346_3_lut_LC_18_5_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i7346_3_lut_LC_18_5_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.i7346_3_lut_LC_18_5_5  (
            .in0(_gnd_net_),
            .in1(N__38432),
            .in2(N__38426),
            .in3(N__42473),
            .lcout(comm_rx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i7_LC_18_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i7_LC_18_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i7_LC_18_6_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i7_LC_18_6_0  (
            .in0(N__38418),
            .in1(N__40628),
            .in2(_gnd_net_),
            .in3(N__38377),
            .lcout(comm_rx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42381),
            .ce(),
            .sr(N__46555));
    defparam \comm_spi.data_rx_i6_LC_18_6_1 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i6_LC_18_6_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i6_LC_18_6_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i6_LC_18_6_1  (
            .in0(N__38376),
            .in1(N__39688),
            .in2(_gnd_net_),
            .in3(N__38417),
            .lcout(comm_rx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42381),
            .ce(),
            .sr(N__46555));
    defparam \comm_spi.data_rx_i5_LC_18_6_2 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i5_LC_18_6_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i5_LC_18_6_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i5_LC_18_6_2  (
            .in0(N__38416),
            .in1(N__39832),
            .in2(_gnd_net_),
            .in3(N__38375),
            .lcout(comm_rx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42381),
            .ce(),
            .sr(N__46555));
    defparam \comm_spi.data_rx_i4_LC_18_6_3 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i4_LC_18_6_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i4_LC_18_6_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i4_LC_18_6_3  (
            .in0(N__38374),
            .in1(N__44807),
            .in2(_gnd_net_),
            .in3(N__38415),
            .lcout(comm_rx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42381),
            .ce(),
            .sr(N__46555));
    defparam \comm_spi.data_rx_i3_LC_18_6_4 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i3_LC_18_6_4 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i3_LC_18_6_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i3_LC_18_6_4  (
            .in0(N__38414),
            .in1(N__40021),
            .in2(_gnd_net_),
            .in3(N__38373),
            .lcout(comm_rx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42381),
            .ce(),
            .sr(N__46555));
    defparam \comm_spi.data_rx_i2_LC_18_6_5 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i2_LC_18_6_5 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i2_LC_18_6_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i2_LC_18_6_5  (
            .in0(N__38372),
            .in1(N__44074),
            .in2(_gnd_net_),
            .in3(N__38413),
            .lcout(comm_rx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42381),
            .ce(),
            .sr(N__46555));
    defparam \comm_spi.data_rx_i1_LC_18_6_6 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i1_LC_18_6_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i1_LC_18_6_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \comm_spi.data_rx_i1_LC_18_6_6  (
            .in0(N__38412),
            .in1(N__38371),
            .in2(_gnd_net_),
            .in3(N__39118),
            .lcout(comm_rx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42381),
            .ce(),
            .sr(N__46555));
    defparam i12171_3_lut_LC_18_6_7.C_ON=1'b0;
    defparam i12171_3_lut_LC_18_6_7.SEQ_MODE=4'b0000;
    defparam i12171_3_lut_LC_18_6_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i12171_3_lut_LC_18_6_7 (
            .in0(N__38978),
            .in1(N__38927),
            .in2(_gnd_net_),
            .in3(N__38689),
            .lcout(n15381),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_378_Mux_3_i7_4_lut_LC_18_7_0.C_ON=1'b0;
    defparam comm_state_3__I_0_378_Mux_3_i7_4_lut_LC_18_7_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_378_Mux_3_i7_4_lut_LC_18_7_0.LUT_INIT=16'b1101110111110000;
    LogicCell40 comm_state_3__I_0_378_Mux_3_i7_4_lut_LC_18_7_0 (
            .in0(N__49735),
            .in1(N__39023),
            .in2(N__42748),
            .in3(N__49550),
            .lcout(),
            .ltout(n12846_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i3_LC_18_7_1.C_ON=1'b0;
    defparam comm_state_i3_LC_18_7_1.SEQ_MODE=4'b1000;
    defparam comm_state_i3_LC_18_7_1.LUT_INIT=16'b0010011100000101;
    LogicCell40 comm_state_i3_LC_18_7_1 (
            .in0(N__52033),
            .in1(N__51923),
            .in2(N__38570),
            .in3(N__39425),
            .lcout(comm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51171),
            .ce(N__38477),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_65_LC_18_7_2.C_ON=1'b0;
    defparam i1_4_lut_adj_65_LC_18_7_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_65_LC_18_7_2.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_65_LC_18_7_2 (
            .in0(N__38567),
            .in1(N__39065),
            .in2(N__42815),
            .in3(N__38486),
            .lcout(n15130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_276_LC_18_7_3.C_ON=1'b0;
    defparam i1_4_lut_adj_276_LC_18_7_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_276_LC_18_7_3.LUT_INIT=16'b1110111011100000;
    LogicCell40 i1_4_lut_adj_276_LC_18_7_3 (
            .in0(N__38533),
            .in1(N__39082),
            .in2(N__43166),
            .in3(N__39073),
            .lcout(),
            .ltout(n4_adj_1184_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_277_LC_18_7_4.C_ON=1'b0;
    defparam i2_4_lut_adj_277_LC_18_7_4.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_277_LC_18_7_4.LUT_INIT=16'b1111000010110000;
    LogicCell40 i2_4_lut_adj_277_LC_18_7_4 (
            .in0(N__49734),
            .in1(N__43379),
            .in2(N__38501),
            .in3(N__50621),
            .lcout(n15108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_174_LC_18_7_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_174_LC_18_7_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_174_LC_18_7_5.LUT_INIT=16'b1110111011111111;
    LogicCell40 i1_2_lut_3_lut_adj_174_LC_18_7_5 (
            .in0(N__52032),
            .in1(N__49733),
            .in2(_gnd_net_),
            .in3(N__49402),
            .lcout(n15241),
            .ltout(n15241_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_285_LC_18_7_6.C_ON=1'b0;
    defparam i1_4_lut_adj_285_LC_18_7_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_285_LC_18_7_6.LUT_INIT=16'b1010001000000000;
    LogicCell40 i1_4_lut_adj_285_LC_18_7_6 (
            .in0(N__43205),
            .in1(N__38498),
            .in2(N__38489),
            .in3(N__38485),
            .lcout(n15128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_18_7_7.C_ON=1'b0;
    defparam i1_3_lut_LC_18_7_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_18_7_7.LUT_INIT=16'b1110111010101010;
    LogicCell40 i1_3_lut_LC_18_7_7 (
            .in0(N__43460),
            .in1(N__39083),
            .in2(_gnd_net_),
            .in3(N__39074),
            .lcout(n15266),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12200_4_lut_LC_18_8_0.C_ON=1'b0;
    defparam i12200_4_lut_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam i12200_4_lut_LC_18_8_0.LUT_INIT=16'b1110111011110000;
    LogicCell40 i12200_4_lut_LC_18_8_0 (
            .in0(N__39041),
            .in1(N__39029),
            .in2(N__39050),
            .in3(N__49438),
            .lcout(),
            .ltout(n15410_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i0_LC_18_8_1.C_ON=1'b0;
    defparam comm_state_i0_LC_18_8_1.SEQ_MODE=4'b1000;
    defparam comm_state_i0_LC_18_8_1.LUT_INIT=16'b0101010111110000;
    LogicCell40 comm_state_i0_LC_18_8_1 (
            .in0(N__51922),
            .in1(_gnd_net_),
            .in2(N__39059),
            .in3(N__52074),
            .lcout(comm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51189),
            .ce(N__39056),
            .sr(_gnd_net_));
    defparam i12198_3_lut_LC_18_8_3.C_ON=1'b0;
    defparam i12198_3_lut_LC_18_8_3.SEQ_MODE=4'b0000;
    defparam i12198_3_lut_LC_18_8_3.LUT_INIT=16'b1110111001010101;
    LogicCell40 i12198_3_lut_LC_18_8_3 (
            .in0(N__50507),
            .in1(N__43391),
            .in2(_gnd_net_),
            .in3(N__49939),
            .lcout(n15408),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7283_2_lut_LC_18_8_4.C_ON=1'b0;
    defparam i7283_2_lut_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam i7283_2_lut_LC_18_8_4.LUT_INIT=16'b1011101110111011;
    LogicCell40 i7283_2_lut_LC_18_8_4 (
            .in0(N__43394),
            .in1(N__50506),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n10394),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12980_3_lut_LC_18_8_5.C_ON=1'b0;
    defparam i12980_3_lut_LC_18_8_5.SEQ_MODE=4'b0000;
    defparam i12980_3_lut_LC_18_8_5.LUT_INIT=16'b1100110010001000;
    LogicCell40 i12980_3_lut_LC_18_8_5 (
            .in0(N__42727),
            .in1(N__49938),
            .in2(_gnd_net_),
            .in3(N__39254),
            .lcout(n16190),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12728_2_lut_3_lut_LC_18_8_6.C_ON=1'b0;
    defparam i12728_2_lut_3_lut_LC_18_8_6.SEQ_MODE=4'b0000;
    defparam i12728_2_lut_3_lut_LC_18_8_6.LUT_INIT=16'b1110111011111111;
    LogicCell40 i12728_2_lut_3_lut_LC_18_8_6 (
            .in0(N__43392),
            .in1(N__42726),
            .in2(_gnd_net_),
            .in3(N__50558),
            .lcout(n15635),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i22_3_lut_4_lut_LC_18_8_7.C_ON=1'b0;
    defparam i22_3_lut_4_lut_LC_18_8_7.SEQ_MODE=4'b0000;
    defparam i22_3_lut_4_lut_LC_18_8_7.LUT_INIT=16'b0001101000001010;
    LogicCell40 i22_3_lut_4_lut_LC_18_8_7 (
            .in0(N__50505),
            .in1(N__43393),
            .in2(N__50143),
            .in3(N__43288),
            .lcout(n7_adj_1190),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9584_3_lut_4_lut_LC_18_9_0.C_ON=1'b0;
    defparam i9584_3_lut_4_lut_LC_18_9_0.SEQ_MODE=4'b0000;
    defparam i9584_3_lut_4_lut_LC_18_9_0.LUT_INIT=16'b1111101011111000;
    LogicCell40 i9584_3_lut_4_lut_LC_18_9_0 (
            .in0(N__44968),
            .in1(N__47496),
            .in2(N__39017),
            .in3(N__40944),
            .lcout(n12622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i31_3_lut_4_lut_3_lut_LC_18_9_2.C_ON=1'b0;
    defparam i31_3_lut_4_lut_3_lut_LC_18_9_2.SEQ_MODE=4'b0000;
    defparam i31_3_lut_4_lut_3_lut_LC_18_9_2.LUT_INIT=16'b0100010000100010;
    LogicCell40 i31_3_lut_4_lut_3_lut_LC_18_9_2 (
            .in0(N__45410),
            .in1(N__47491),
            .in2(_gnd_net_),
            .in3(N__45221),
            .lcout(n14_adj_1152),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_53_LC_18_9_3.C_ON=1'b0;
    defparam i1_4_lut_adj_53_LC_18_9_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_53_LC_18_9_3.LUT_INIT=16'b1011000011100000;
    LogicCell40 i1_4_lut_adj_53_LC_18_9_3 (
            .in0(N__46963),
            .in1(N__39552),
            .in2(N__40225),
            .in3(N__45413),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12103_3_lut_4_lut_LC_18_9_4.C_ON=1'b0;
    defparam i12103_3_lut_4_lut_LC_18_9_4.SEQ_MODE=4'b0000;
    defparam i12103_3_lut_4_lut_LC_18_9_4.LUT_INIT=16'b1111111110111111;
    LogicCell40 i12103_3_lut_4_lut_LC_18_9_4 (
            .in0(N__45412),
            .in1(N__47495),
            .in2(N__47181),
            .in3(N__40860),
            .lcout(),
            .ltout(n15309_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_39_LC_18_9_5.C_ON=1'b0;
    defparam i1_4_lut_adj_39_LC_18_9_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_39_LC_18_9_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 i1_4_lut_adj_39_LC_18_9_5 (
            .in0(N__39452),
            .in1(N__39416),
            .in2(N__39446),
            .in3(N__40793),
            .lcout(comm_state_3_N_418_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12762_2_lut_LC_18_9_6.C_ON=1'b0;
    defparam i12762_2_lut_LC_18_9_6.SEQ_MODE=4'b0000;
    defparam i12762_2_lut_LC_18_9_6.LUT_INIT=16'b0011001100000000;
    LogicCell40 i12762_2_lut_LC_18_9_6 (
            .in0(_gnd_net_),
            .in1(N__50513),
            .in2(_gnd_net_),
            .in3(N__39436),
            .lcout(n15637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_119_i13_2_lut_3_lut_4_lut_LC_18_9_7.C_ON=1'b0;
    defparam equal_119_i13_2_lut_3_lut_4_lut_LC_18_9_7.SEQ_MODE=4'b0000;
    defparam equal_119_i13_2_lut_3_lut_4_lut_LC_18_9_7.LUT_INIT=16'b1111111111111011;
    LogicCell40 equal_119_i13_2_lut_3_lut_4_lut_LC_18_9_7 (
            .in0(N__45222),
            .in1(N__45411),
            .in2(N__47601),
            .in3(N__41211),
            .lcout(n13_adj_1040),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_18_10_0.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_18_10_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_18_10_0.LUT_INIT=16'b0111010100000000;
    LogicCell40 i1_3_lut_4_lut_LC_18_10_0 (
            .in0(N__45455),
            .in1(N__45041),
            .in2(N__47741),
            .in3(N__46898),
            .lcout(n22_adj_1078),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i7_LC_18_10_1.C_ON=1'b0;
    defparam comm_cmd_i7_LC_18_10_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i7_LC_18_10_1.LUT_INIT=16'b1101100001010000;
    LogicCell40 comm_cmd_i7_LC_18_10_1 (
            .in0(N__44035),
            .in1(N__43995),
            .in2(N__39255),
            .in3(N__39307),
            .lcout(comm_cmd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51224),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i0_LC_18_10_2.C_ON=1'b0;
    defparam comm_cmd_i0_LC_18_10_2.SEQ_MODE=4'b1000;
    defparam comm_cmd_i0_LC_18_10_2.LUT_INIT=16'b1110001000100010;
    LogicCell40 comm_cmd_i0_LC_18_10_2 (
            .in0(N__47599),
            .in1(N__44032),
            .in2(N__44002),
            .in3(N__39142),
            .lcout(comm_cmd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51224),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i2_LC_18_10_3.C_ON=1'b0;
    defparam comm_cmd_i2_LC_18_10_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i2_LC_18_10_3.LUT_INIT=16'b1101100001010000;
    LogicCell40 comm_cmd_i2_LC_18_10_3 (
            .in0(N__44033),
            .in1(N__43994),
            .in2(N__45465),
            .in3(N__40036),
            .lcout(comm_cmd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51224),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_114_i8_2_lut_LC_18_10_4.C_ON=1'b0;
    defparam equal_114_i8_2_lut_LC_18_10_4.SEQ_MODE=4'b0000;
    defparam equal_114_i8_2_lut_LC_18_10_4.LUT_INIT=16'b1111111100110011;
    LogicCell40 equal_114_i8_2_lut_LC_18_10_4 (
            .in0(_gnd_net_),
            .in1(N__45405),
            .in2(_gnd_net_),
            .in3(N__45040),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i2_LC_18_10_5.C_ON=1'b0;
    defparam buf_dds_i2_LC_18_10_5.SEQ_MODE=4'b1000;
    defparam buf_dds_i2_LC_18_10_5.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i2_LC_18_10_5 (
            .in0(N__39998),
            .in1(N__43681),
            .in2(N__41519),
            .in3(N__41378),
            .lcout(buf_dds_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51224),
            .ce(),
            .sr(_gnd_net_));
    defparam i7266_2_lut_LC_18_10_6.C_ON=1'b0;
    defparam i7266_2_lut_LC_18_10_6.SEQ_MODE=4'b0000;
    defparam i7266_2_lut_LC_18_10_6.LUT_INIT=16'b0011001100000000;
    LogicCell40 i7266_2_lut_LC_18_10_6 (
            .in0(_gnd_net_),
            .in1(N__52082),
            .in2(_gnd_net_),
            .in3(N__49965),
            .lcout(n10363),
            .ltout(n10363_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i4_LC_18_10_7.C_ON=1'b0;
    defparam comm_cmd_i4_LC_18_10_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i4_LC_18_10_7.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i4_LC_18_10_7 (
            .in0(N__44034),
            .in1(N__39878),
            .in2(N__39812),
            .in3(N__40288),
            .lcout(comm_cmd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51224),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i3_LC_18_11_0.C_ON=1'b0;
    defparam comm_cmd_i3_LC_18_11_0.SEQ_MODE=4'b1000;
    defparam comm_cmd_i3_LC_18_11_0.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i3_LC_18_11_0 (
            .in0(N__43996),
            .in1(N__44039),
            .in2(N__44883),
            .in3(N__46818),
            .lcout(comm_cmd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51241),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i5_LC_18_11_1.C_ON=1'b0;
    defparam comm_cmd_i5_LC_18_11_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i5_LC_18_11_1.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i5_LC_18_11_1 (
            .in0(N__40303),
            .in1(N__43997),
            .in2(N__39731),
            .in3(N__44041),
            .lcout(comm_cmd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51241),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_6__355_LC_18_11_2.C_ON=1'b0;
    defparam buf_control_6__355_LC_18_11_2.SEQ_MODE=4'b1000;
    defparam buf_control_6__355_LC_18_11_2.LUT_INIT=16'b1111000011011000;
    LogicCell40 buf_control_6__355_LC_18_11_2 (
            .in0(N__39665),
            .in1(N__41895),
            .in2(N__42986),
            .in3(N__41126),
            .lcout(buf_control_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51241),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_18_11_3.C_ON=1'b0;
    defparam i2_3_lut_LC_18_11_3.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_18_11_3.LUT_INIT=16'b1111111110111011;
    LogicCell40 i2_3_lut_LC_18_11_3 (
            .in0(N__40302),
            .in1(N__40284),
            .in2(_gnd_net_),
            .in3(N__40266),
            .lcout(n8085),
            .ltout(n8085_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_251_LC_18_11_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_251_LC_18_11_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_251_LC_18_11_4.LUT_INIT=16'b1111110011111111;
    LogicCell40 i1_2_lut_3_lut_adj_251_LC_18_11_4 (
            .in0(_gnd_net_),
            .in1(N__47488),
            .in2(N__39593),
            .in3(N__46817),
            .lcout(n8094),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_2_lut_LC_18_11_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_2_lut_LC_18_11_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_2_lut_LC_18_11_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 i1_2_lut_3_lut_2_lut_LC_18_11_5 (
            .in0(N__47489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45058),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i6_LC_18_11_6.C_ON=1'b0;
    defparam comm_cmd_i6_LC_18_11_6.SEQ_MODE=4'b1000;
    defparam comm_cmd_i6_LC_18_11_6.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i6_LC_18_11_6 (
            .in0(N__40267),
            .in1(N__40657),
            .in2(N__44003),
            .in3(N__44040),
            .lcout(comm_cmd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51241),
            .ce(),
            .sr(_gnd_net_));
    defparam i129_4_lut_adj_104_LC_18_11_7.C_ON=1'b0;
    defparam i129_4_lut_adj_104_LC_18_11_7.SEQ_MODE=4'b0000;
    defparam i129_4_lut_adj_104_LC_18_11_7.LUT_INIT=16'b0100010010100000;
    LogicCell40 i129_4_lut_adj_104_LC_18_11_7 (
            .in0(N__47490),
            .in1(N__40595),
            .in2(N__40583),
            .in3(N__45059),
            .lcout(n75),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_300_LC_18_12_1.C_ON=1'b0;
    defparam i1_2_lut_adj_300_LC_18_12_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_300_LC_18_12_1.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_300_LC_18_12_1 (
            .in0(_gnd_net_),
            .in1(N__46819),
            .in2(_gnd_net_),
            .in3(N__40830),
            .lcout(n12),
            .ltout(n12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2992_3_lut_4_lut_LC_18_12_2.C_ON=1'b0;
    defparam i2992_3_lut_4_lut_LC_18_12_2.SEQ_MODE=4'b0000;
    defparam i2992_3_lut_4_lut_LC_18_12_2.LUT_INIT=16'b1111111111111011;
    LogicCell40 i2992_3_lut_4_lut_LC_18_12_2 (
            .in0(N__50537),
            .in1(N__47602),
            .in2(N__40550),
            .in3(N__40946),
            .lcout(n6301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9546_2_lut_3_lut_3_lut_3_lut_LC_18_12_3.C_ON=1'b0;
    defparam i9546_2_lut_3_lut_3_lut_3_lut_LC_18_12_3.SEQ_MODE=4'b0000;
    defparam i9546_2_lut_3_lut_3_lut_3_lut_LC_18_12_3.LUT_INIT=16'b1111111110011001;
    LogicCell40 i9546_2_lut_3_lut_3_lut_3_lut_LC_18_12_3 (
            .in0(N__47603),
            .in1(N__45539),
            .in2(_gnd_net_),
            .in3(N__45105),
            .lcout(n12702),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i2_LC_18_12_4.C_ON=1'b0;
    defparam req_data_cnt_i2_LC_18_12_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i2_LC_18_12_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i2_LC_18_12_4 (
            .in0(N__40456),
            .in1(N__40349),
            .in2(_gnd_net_),
            .in3(N__40323),
            .lcout(req_data_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51256),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_297_LC_18_12_5.C_ON=1'b0;
    defparam i1_3_lut_adj_297_LC_18_12_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_297_LC_18_12_5.LUT_INIT=16'b0000000001000100;
    LogicCell40 i1_3_lut_adj_297_LC_18_12_5 (
            .in0(N__40304),
            .in1(N__40289),
            .in2(_gnd_net_),
            .in3(N__40268),
            .lcout(n8043),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_18_12_6.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_18_12_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_18_12_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_4_lut_LC_18_12_6 (
            .in0(N__45540),
            .in1(N__47604),
            .in2(N__45215),
            .in3(N__41210),
            .lcout(n7511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i1_LC_18_12_7.C_ON=1'b0;
    defparam buf_dds_i1_LC_18_12_7.SEQ_MODE=4'b1000;
    defparam buf_dds_i1_LC_18_12_7.LUT_INIT=16'b1101100001010000;
    LogicCell40 buf_dds_i1_LC_18_12_7 (
            .in0(N__41368),
            .in1(N__41524),
            .in2(N__42124),
            .in3(N__41097),
            .lcout(buf_dds_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51256),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_84_LC_18_13_0.C_ON=1'b0;
    defparam i1_4_lut_adj_84_LC_18_13_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_84_LC_18_13_0.LUT_INIT=16'b1010000010100010;
    LogicCell40 i1_4_lut_adj_84_LC_18_13_0 (
            .in0(N__52081),
            .in1(N__41180),
            .in2(N__51825),
            .in3(N__50594),
            .lcout(n8250),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_290_LC_18_13_2.C_ON=1'b0;
    defparam i1_4_lut_adj_290_LC_18_13_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_290_LC_18_13_2.LUT_INIT=16'b1110110010100000;
    LogicCell40 i1_4_lut_adj_290_LC_18_13_2 (
            .in0(N__45544),
            .in1(N__41040),
            .in2(N__41002),
            .in3(N__45153),
            .lcout(n78_adj_1022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i4_3_lut_LC_18_13_4.C_ON=1'b0;
    defparam mux_1498_i4_3_lut_LC_18_13_4.SEQ_MODE=4'b0000;
    defparam mux_1498_i4_3_lut_LC_18_13_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_1498_i4_3_lut_LC_18_13_4 (
            .in0(N__40970),
            .in1(N__47636),
            .in2(_gnd_net_),
            .in3(N__43774),
            .lcout(n4206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12098_3_lut_4_lut_LC_18_13_5.C_ON=1'b0;
    defparam i12098_3_lut_4_lut_LC_18_13_5.SEQ_MODE=4'b0000;
    defparam i12098_3_lut_4_lut_LC_18_13_5.LUT_INIT=16'b1111111100101111;
    LogicCell40 i12098_3_lut_4_lut_LC_18_13_5 (
            .in0(N__40945),
            .in1(N__41913),
            .in2(N__47790),
            .in3(N__41200),
            .lcout(n15188),
            .ltout(n15188_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_18_13_6.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_18_13_6.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_18_13_6.LUT_INIT=16'b1111000011100000;
    LogicCell40 i2_3_lut_4_lut_LC_18_13_6 (
            .in0(N__40906),
            .in1(N__46931),
            .in2(N__40889),
            .in3(N__40859),
            .lcout(),
            .ltout(n6_adj_1171_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_4_lut_LC_18_13_7.C_ON=1'b0;
    defparam i3_4_lut_4_lut_LC_18_13_7.SEQ_MODE=4'b0000;
    defparam i3_4_lut_4_lut_LC_18_13_7.LUT_INIT=16'b1101000011100000;
    LogicCell40 i3_4_lut_4_lut_LC_18_13_7 (
            .in0(N__45154),
            .in1(N__43636),
            .in2(N__40796),
            .in3(N__45545),
            .lcout(n15190),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i12_LC_18_14_0 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i12_LC_18_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i12_LC_18_14_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i12_LC_18_14_0  (
            .in0(N__49220),
            .in1(N__44382),
            .in2(N__40782),
            .in3(N__48598),
            .lcout(buf_adcdata3_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51285),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i21_LC_18_14_1 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i21_LC_18_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i21_LC_18_14_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i21_LC_18_14_1  (
            .in0(N__41949),
            .in1(N__49221),
            .in2(N__48599),
            .in3(N__48832),
            .lcout(cmd_rdadctmp_21_adj_1091),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51285),
            .ce(),
            .sr(_gnd_net_));
    defparam i9560_2_lut_LC_18_14_2.C_ON=1'b0;
    defparam i9560_2_lut_LC_18_14_2.SEQ_MODE=4'b0000;
    defparam i9560_2_lut_LC_18_14_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 i9560_2_lut_LC_18_14_2 (
            .in0(_gnd_net_),
            .in1(N__45541),
            .in2(_gnd_net_),
            .in3(N__45151),
            .lcout(n4_adj_1041),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i14_LC_18_14_4.C_ON=1'b0;
    defparam acadc_skipCount_i14_LC_18_14_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i14_LC_18_14_4.LUT_INIT=16'b0011101100001000;
    LogicCell40 acadc_skipCount_i14_LC_18_14_4 (
            .in0(N__41894),
            .in1(N__41756),
            .in2(N__51930),
            .in3(N__41697),
            .lcout(acadc_skipCount_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51285),
            .ce(),
            .sr(_gnd_net_));
    defparam i12647_4_lut_LC_18_14_5.C_ON=1'b0;
    defparam i12647_4_lut_LC_18_14_5.SEQ_MODE=4'b0000;
    defparam i12647_4_lut_LC_18_14_5.LUT_INIT=16'b1100010010000000;
    LogicCell40 i12647_4_lut_LC_18_14_5 (
            .in0(N__45542),
            .in1(N__46946),
            .in2(N__41674),
            .in3(N__41652),
            .lcout(n15468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i5_3_lut_LC_18_14_6.C_ON=1'b0;
    defparam mux_1511_i5_3_lut_LC_18_14_6.SEQ_MODE=4'b0000;
    defparam mux_1511_i5_3_lut_LC_18_14_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_1511_i5_3_lut_LC_18_14_6 (
            .in0(N__41615),
            .in1(N__45543),
            .in2(_gnd_net_),
            .in3(N__41606),
            .lcout(n4250),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i14_LC_18_15_0 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i14_LC_18_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i14_LC_18_15_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \ADC_VAC3.ADC_DATA_i14_LC_18_15_0  (
            .in0(N__41550),
            .in1(N__41578),
            .in2(N__49266),
            .in3(N__44399),
            .lcout(buf_adcdata3_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51296),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds_i11_LC_18_15_1.C_ON=1'b0;
    defparam buf_dds_i11_LC_18_15_1.SEQ_MODE=4'b1000;
    defparam buf_dds_i11_LC_18_15_1.LUT_INIT=16'b1010000011001100;
    LogicCell40 buf_dds_i11_LC_18_15_1 (
            .in0(N__43562),
            .in1(N__41241),
            .in2(N__41528),
            .in3(N__41379),
            .lcout(buf_dds_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51296),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_208_i13_2_lut_3_lut_4_lut_LC_18_15_3.C_ON=1'b0;
    defparam equal_208_i13_2_lut_3_lut_4_lut_LC_18_15_3.SEQ_MODE=4'b0000;
    defparam equal_208_i13_2_lut_3_lut_4_lut_LC_18_15_3.LUT_INIT=16'b1111111011111111;
    LogicCell40 equal_208_i13_2_lut_3_lut_4_lut_LC_18_15_3 (
            .in0(N__45234),
            .in1(N__45605),
            .in2(N__41222),
            .in3(N__47795),
            .lcout(n13_adj_1025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1502_i2_3_lut_LC_18_15_4.C_ON=1'b0;
    defparam mux_1502_i2_3_lut_LC_18_15_4.SEQ_MODE=4'b0000;
    defparam mux_1502_i2_3_lut_LC_18_15_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_1502_i2_3_lut_LC_18_15_4 (
            .in0(N__47797),
            .in1(N__42191),
            .in2(_gnd_net_),
            .in3(N__42160),
            .lcout(),
            .ltout(n4220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i2_3_lut_LC_18_15_5.C_ON=1'b0;
    defparam mux_1511_i2_3_lut_LC_18_15_5.SEQ_MODE=4'b0000;
    defparam mux_1511_i2_3_lut_LC_18_15_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_1511_i2_3_lut_LC_18_15_5 (
            .in0(_gnd_net_),
            .in1(N__42041),
            .in2(N__42143),
            .in3(N__45606),
            .lcout(),
            .ltout(n4253_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1513_i2_4_lut_LC_18_15_6.C_ON=1'b0;
    defparam mux_1513_i2_4_lut_LC_18_15_6.SEQ_MODE=4'b0000;
    defparam mux_1513_i2_4_lut_LC_18_15_6.LUT_INIT=16'b1111000000100010;
    LogicCell40 mux_1513_i2_4_lut_LC_18_15_6 (
            .in0(N__42068),
            .in1(N__45235),
            .in2(N__42140),
            .in3(N__46965),
            .lcout(n4263),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i2_3_lut_LC_18_15_7.C_ON=1'b0;
    defparam mux_1498_i2_3_lut_LC_18_15_7.SEQ_MODE=4'b0000;
    defparam mux_1498_i2_3_lut_LC_18_15_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_1498_i2_3_lut_LC_18_15_7 (
            .in0(N__42120),
            .in1(N__42088),
            .in2(_gnd_net_),
            .in3(N__47796),
            .lcout(n4208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i2_4_lut_LC_18_16_0.C_ON=1'b0;
    defparam mux_1507_i2_4_lut_LC_18_16_0.SEQ_MODE=4'b0000;
    defparam mux_1507_i2_4_lut_LC_18_16_0.LUT_INIT=16'b0111001101000000;
    LogicCell40 mux_1507_i2_4_lut_LC_18_16_0 (
            .in0(N__47800),
            .in1(N__45236),
            .in2(N__42062),
            .in3(N__42047),
            .lcout(n4233),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1494_i4_3_lut_LC_18_16_2.C_ON=1'b0;
    defparam mux_1494_i4_3_lut_LC_18_16_2.SEQ_MODE=4'b0000;
    defparam mux_1494_i4_3_lut_LC_18_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_1494_i4_3_lut_LC_18_16_2 (
            .in0(N__42035),
            .in1(N__47802),
            .in2(_gnd_net_),
            .in3(N__42017),
            .lcout(),
            .ltout(n4194_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1507_i4_4_lut_LC_18_16_3.C_ON=1'b0;
    defparam mux_1507_i4_4_lut_LC_18_16_3.SEQ_MODE=4'b0000;
    defparam mux_1507_i4_4_lut_LC_18_16_3.LUT_INIT=16'b1111101011011000;
    LogicCell40 mux_1507_i4_4_lut_LC_18_16_3 (
            .in0(N__45237),
            .in1(N__41996),
            .in2(N__41981),
            .in3(N__47801),
            .lcout(),
            .ltout(n4231_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1511_i4_3_lut_LC_18_16_4.C_ON=1'b0;
    defparam mux_1511_i4_3_lut_LC_18_16_4.SEQ_MODE=4'b0000;
    defparam mux_1511_i4_3_lut_LC_18_16_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_1511_i4_3_lut_LC_18_16_4 (
            .in0(_gnd_net_),
            .in1(N__41978),
            .in2(N__41972),
            .in3(N__45607),
            .lcout(),
            .ltout(n4251_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1513_i4_4_lut_LC_18_16_5.C_ON=1'b0;
    defparam mux_1513_i4_4_lut_LC_18_16_5.SEQ_MODE=4'b0000;
    defparam mux_1513_i4_4_lut_LC_18_16_5.LUT_INIT=16'b1111000001000100;
    LogicCell40 mux_1513_i4_4_lut_LC_18_16_5 (
            .in0(N__45238),
            .in1(N__41969),
            .in2(N__41960),
            .in3(N__46966),
            .lcout(n4261),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1457_i2_4_lut_LC_18_17_4.C_ON=1'b0;
    defparam mux_1457_i2_4_lut_LC_18_17_4.SEQ_MODE=4'b0000;
    defparam mux_1457_i2_4_lut_LC_18_17_4.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1457_i2_4_lut_LC_18_17_4 (
            .in0(N__42686),
            .in1(N__47803),
            .in2(N__42674),
            .in3(N__46964),
            .lcout(n4063),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i11_LC_18_18_3 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i11_LC_18_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i11_LC_18_18_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i11_LC_18_18_3  (
            .in0(N__53810),
            .in1(N__53492),
            .in2(N__46181),
            .in3(N__42616),
            .lcout(buf_adcdata2_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51312),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_8_i15_4_lut_LC_18_19_2.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_8_i15_4_lut_LC_18_19_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_8_i15_4_lut_LC_18_19_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_394_Mux_8_i15_4_lut_LC_18_19_2 (
            .in0(N__52183),
            .in1(N__42602),
            .in2(N__51929),
            .in3(N__42581),
            .lcout(data_index_9_N_258_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_7330_7331_set_LC_19_4_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_7330_7331_set_LC_19_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imosi_44_7330_7331_set_LC_19_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_7330_7331_set_LC_19_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45795),
            .lcout(\comm_spi.n10441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51146),
            .ce(),
            .sr(N__42953));
    defparam \comm_spi.data_rx_i0_7344_7345_reset_LC_19_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_7344_7345_reset_LC_19_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i0_7344_7345_reset_LC_19_5_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_rx_i0_7344_7345_reset_LC_19_5_0  (
            .in0(N__42228),
            .in1(N__42253),
            .in2(_gnd_net_),
            .in3(N__45814),
            .lcout(\comm_spi.n10456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42375),
            .ce(),
            .sr(N__42878));
    defparam \comm_spi.i13072_4_lut_3_lut_LC_19_6_1 .C_ON=1'b0;
    defparam \comm_spi.i13072_4_lut_3_lut_LC_19_6_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13072_4_lut_3_lut_LC_19_6_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.i13072_4_lut_3_lut_LC_19_6_1  (
            .in0(N__45797),
            .in1(N__46462),
            .in2(_gnd_net_),
            .in3(N__42252),
            .lcout(\comm_spi.n16893 ),
            .ltout(\comm_spi.n16893_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i7332_3_lut_LC_19_6_2 .C_ON=1'b0;
    defparam \comm_spi.i7332_3_lut_LC_19_6_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i7332_3_lut_LC_19_6_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.i7332_3_lut_LC_19_6_2  (
            .in0(_gnd_net_),
            .in1(N__42232),
            .in2(N__42209),
            .in3(N__45813),
            .lcout(\comm_spi.imosi ),
            .ltout(\comm_spi.imosi_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_19_6_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_19_6_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_19_6_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \comm_spi.RESET_I_0_86_2_lut_LC_19_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42206),
            .in3(N__46464),
            .lcout(\comm_spi.DOUT_7__N_785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_19_6_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_19_6_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_19_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_88_2_lut_LC_19_6_4  (
            .in0(N__46463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45796),
            .lcout(\comm_spi.imosi_N_791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i1_LC_19_6_5 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i1_LC_19_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i1_LC_19_6_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i1_LC_19_6_5  (
            .in0(N__53751),
            .in1(N__42904),
            .in2(N__42944),
            .in3(N__53533),
            .lcout(buf_adcdata2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51172),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_19_6_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_19_6_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_19_6_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.RESET_I_0_87_2_lut_LC_19_6_7  (
            .in0(_gnd_net_),
            .in1(N__46465),
            .in2(_gnd_net_),
            .in3(N__42890),
            .lcout(\comm_spi.DOUT_7__N_786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_274_LC_19_7_0.C_ON=1'b0;
    defparam i1_4_lut_adj_274_LC_19_7_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_274_LC_19_7_0.LUT_INIT=16'b1000101010001000;
    LogicCell40 i1_4_lut_adj_274_LC_19_7_0 (
            .in0(N__42849),
            .in1(N__42811),
            .in2(N__50550),
            .in3(N__43614),
            .lcout(n15191),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2727_2_lut_LC_19_7_2.C_ON=1'b0;
    defparam i2727_2_lut_LC_19_7_2.SEQ_MODE=4'b0000;
    defparam i2727_2_lut_LC_19_7_2.LUT_INIT=16'b1111111110101010;
    LogicCell40 i2727_2_lut_LC_19_7_2 (
            .in0(N__50476),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50282),
            .lcout(n10148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_clear_330_LC_19_7_3.C_ON=1'b0;
    defparam comm_clear_330_LC_19_7_3.SEQ_MODE=4'b1000;
    defparam comm_clear_330_LC_19_7_3.LUT_INIT=16'b0101010111011101;
    LogicCell40 comm_clear_330_LC_19_7_3 (
            .in0(N__50283),
            .in1(N__50477),
            .in2(_gnd_net_),
            .in3(N__52073),
            .lcout(comm_clear),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51190),
            .ce(N__50633),
            .sr(_gnd_net_));
    defparam i22_4_lut_LC_19_8_1.C_ON=1'b0;
    defparam i22_4_lut_LC_19_8_1.SEQ_MODE=4'b0000;
    defparam i22_4_lut_LC_19_8_1.LUT_INIT=16'b1011001110100010;
    LogicCell40 i22_4_lut_LC_19_8_1 (
            .in0(N__49434),
            .in1(N__50559),
            .in2(N__42731),
            .in3(N__43301),
            .lcout(n8_adj_1193),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12879_4_lut_LC_19_8_2.C_ON=1'b0;
    defparam i12879_4_lut_LC_19_8_2.SEQ_MODE=4'b0000;
    defparam i12879_4_lut_LC_19_8_2.LUT_INIT=16'b0000100001001100;
    LogicCell40 i12879_4_lut_LC_19_8_2 (
            .in0(N__50560),
            .in1(N__49435),
            .in2(N__43436),
            .in3(N__42707),
            .lcout(),
            .ltout(n15711_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i2_LC_19_8_3.C_ON=1'b0;
    defparam comm_state_i2_LC_19_8_3.SEQ_MODE=4'b1000;
    defparam comm_state_i2_LC_19_8_3.LUT_INIT=16'b0111001001010000;
    LogicCell40 comm_state_i2_LC_19_8_3 (
            .in0(N__50286),
            .in1(N__43398),
            .in2(N__42695),
            .in3(N__42692),
            .lcout(comm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51207),
            .ce(N__43469),
            .sr(N__52424));
    defparam i1_4_lut_adj_41_LC_19_8_4.C_ON=1'b0;
    defparam i1_4_lut_adj_41_LC_19_8_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_41_LC_19_8_4.LUT_INIT=16'b0000001010111100;
    LogicCell40 i1_4_lut_adj_41_LC_19_8_4 (
            .in0(N__43300),
            .in1(N__50285),
            .in2(N__43437),
            .in3(N__49433),
            .lcout(),
            .ltout(n26_adj_1192_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13040_2_lut_3_lut_LC_19_8_5.C_ON=1'b0;
    defparam i13040_2_lut_3_lut_LC_19_8_5.SEQ_MODE=4'b0000;
    defparam i13040_2_lut_3_lut_LC_19_8_5.LUT_INIT=16'b1101111111011111;
    LogicCell40 i13040_2_lut_3_lut_LC_19_8_5 (
            .in0(N__50504),
            .in1(N__52062),
            .in2(N__43472),
            .in3(_gnd_net_),
            .lcout(n18_adj_1191),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_229_LC_19_8_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_229_LC_19_8_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_229_LC_19_8_6.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_229_LC_19_8_6 (
            .in0(N__52061),
            .in1(N__50284),
            .in2(_gnd_net_),
            .in3(N__49432),
            .lcout(n15245),
            .ltout(n15245_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_LC_19_8_7.C_ON=1'b0;
    defparam i1_4_lut_4_lut_LC_19_8_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_LC_19_8_7.LUT_INIT=16'b1111010111111100;
    LogicCell40 i1_4_lut_4_lut_LC_19_8_7 (
            .in0(N__50503),
            .in1(N__43402),
            .in2(N__43304),
            .in3(N__43299),
            .lcout(n8544),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_206_i9_2_lut_3_lut_LC_19_9_0.C_ON=1'b0;
    defparam equal_206_i9_2_lut_3_lut_LC_19_9_0.SEQ_MODE=4'b0000;
    defparam equal_206_i9_2_lut_3_lut_LC_19_9_0.LUT_INIT=16'b1110111011111111;
    LogicCell40 equal_206_i9_2_lut_3_lut_LC_19_9_0 (
            .in0(N__47542),
            .in1(N__45437),
            .in2(_gnd_net_),
            .in3(N__45225),
            .lcout(n9_adj_1028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_177_LC_19_9_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_177_LC_19_9_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_177_LC_19_9_3.LUT_INIT=16'b1111111111011101;
    LogicCell40 i1_2_lut_3_lut_adj_177_LC_19_9_3 (
            .in0(N__52185),
            .in1(N__50093),
            .in2(_gnd_net_),
            .in3(N__49403),
            .lcout(n9011),
            .ltout(n9011_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_287_LC_19_9_4.C_ON=1'b0;
    defparam i1_4_lut_adj_287_LC_19_9_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_287_LC_19_9_4.LUT_INIT=16'b1110000011000000;
    LogicCell40 i1_4_lut_adj_287_LC_19_9_4 (
            .in0(N__49404),
            .in1(N__52186),
            .in2(N__43142),
            .in3(N__45689),
            .lcout(n9215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1469_i4_4_lut_LC_19_9_5.C_ON=1'b0;
    defparam mux_1469_i4_4_lut_LC_19_9_5.SEQ_MODE=4'b0000;
    defparam mux_1469_i4_4_lut_LC_19_9_5.LUT_INIT=16'b1010001110100000;
    LogicCell40 mux_1469_i4_4_lut_LC_19_9_5 (
            .in0(N__43040),
            .in1(N__47543),
            .in2(N__47182),
            .in3(N__43024),
            .lcout(comm_buf_3_7_N_501_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i111_4_lut_adj_133_LC_19_10_0.C_ON=1'b0;
    defparam i111_4_lut_adj_133_LC_19_10_0.SEQ_MODE=4'b0000;
    defparam i111_4_lut_adj_133_LC_19_10_0.LUT_INIT=16'b0011000010001000;
    LogicCell40 i111_4_lut_adj_133_LC_19_10_0 (
            .in0(N__43707),
            .in1(N__45464),
            .in2(N__42985),
            .in3(N__46910),
            .lcout(n60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i0_LC_19_10_1 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i0_LC_19_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i0_LC_19_10_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC3.ADC_DATA_i0_LC_19_10_1  (
            .in0(N__44400),
            .in1(N__43800),
            .in2(N__43853),
            .in3(N__49265),
            .lcout(buf_adcdata3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51242),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i11_LC_19_10_2 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i11_LC_19_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i11_LC_19_10_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i11_LC_19_10_2  (
            .in0(N__49262),
            .in1(N__44401),
            .in2(N__49286),
            .in3(N__43767),
            .lcout(buf_adcdata3_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51242),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i22_LC_19_10_3 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i22_LC_19_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i22_LC_19_10_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i22_LC_19_10_3  (
            .in0(N__44402),
            .in1(N__49263),
            .in2(N__43748),
            .in3(N__43708),
            .lcout(buf_adcdata3_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51242),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_4_lut_adj_272_LC_19_10_4.C_ON=1'b0;
    defparam i1_4_lut_4_lut_4_lut_adj_272_LC_19_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_4_lut_adj_272_LC_19_10_4.LUT_INIT=16'b1110001111100000;
    LogicCell40 i1_4_lut_4_lut_4_lut_adj_272_LC_19_10_4 (
            .in0(N__50108),
            .in1(N__49469),
            .in2(N__52423),
            .in3(N__43694),
            .lcout(n8618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1498_i3_3_lut_LC_19_10_5.C_ON=1'b0;
    defparam mux_1498_i3_3_lut_LC_19_10_5.SEQ_MODE=4'b0000;
    defparam mux_1498_i3_3_lut_LC_19_10_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_1498_i3_3_lut_LC_19_10_5 (
            .in0(N__43677),
            .in1(N__44199),
            .in2(_gnd_net_),
            .in3(N__47600),
            .lcout(n4207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i19_LC_19_10_7 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i19_LC_19_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i19_LC_19_10_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i19_LC_19_10_7  (
            .in0(N__44509),
            .in1(N__49281),
            .in2(N__48845),
            .in3(N__49264),
            .lcout(cmd_rdadctmp_19_adj_1093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51242),
            .ce(),
            .sr(_gnd_net_));
    defparam i13023_2_lut_3_lut_LC_19_11_0.C_ON=1'b0;
    defparam i13023_2_lut_3_lut_LC_19_11_0.SEQ_MODE=4'b0000;
    defparam i13023_2_lut_3_lut_LC_19_11_0.LUT_INIT=16'b0100010000000000;
    LogicCell40 i13023_2_lut_3_lut_LC_19_11_0 (
            .in0(N__43635),
            .in1(N__45409),
            .in2(_gnd_net_),
            .in3(N__45042),
            .lcout(n729),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i19_LC_19_11_1 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i19_LC_19_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i19_LC_19_11_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i19_LC_19_11_1  (
            .in0(N__53774),
            .in1(N__43576),
            .in2(N__43877),
            .in3(N__53569),
            .lcout(buf_adcdata2_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51257),
            .ce(),
            .sr(_gnd_net_));
    defparam i9629_2_lut_3_lut_LC_19_11_2.C_ON=1'b0;
    defparam i9629_2_lut_3_lut_LC_19_11_2.SEQ_MODE=4'b0000;
    defparam i9629_2_lut_3_lut_LC_19_11_2.LUT_INIT=16'b0000000001000100;
    LogicCell40 i9629_2_lut_3_lut_LC_19_11_2 (
            .in0(N__50106),
            .in1(N__43559),
            .in2(_gnd_net_),
            .in3(N__49445),
            .lcout(n14_adj_1208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i2_LC_19_11_3 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i2_LC_19_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i2_LC_19_11_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i2_LC_19_11_3  (
            .in0(N__53116),
            .in1(N__44419),
            .in2(N__44471),
            .in3(N__52892),
            .lcout(buf_adcdata1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51257),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.ADC_DATA_i10_LC_19_11_6 .C_ON=1'b0;
    defparam \ADC_VAC3.ADC_DATA_i10_LC_19_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.ADC_DATA_i10_LC_19_11_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC3.ADC_DATA_i10_LC_19_11_6  (
            .in0(N__44405),
            .in1(N__49243),
            .in2(N__44206),
            .in3(N__44510),
            .lcout(buf_adcdata3_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51257),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i1_LC_19_11_7.C_ON=1'b0;
    defparam comm_cmd_i1_LC_19_11_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i1_LC_19_11_7.LUT_INIT=16'b1100101000001010;
    LogicCell40 comm_cmd_i1_LC_19_11_7 (
            .in0(N__45043),
            .in1(N__44139),
            .in2(N__44042),
            .in3(N__44001),
            .lcout(comm_cmd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51257),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i26_LC_19_12_0 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i26_LC_19_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i26_LC_19_12_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i26_LC_19_12_0  (
            .in0(N__53534),
            .in1(N__43967),
            .in2(N__43892),
            .in3(N__46115),
            .lcout(cmd_rdadctmp_26_adj_1050),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51273),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i18_LC_19_12_1 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i18_LC_19_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i18_LC_19_12_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i18_LC_19_12_1  (
            .in0(N__53813),
            .in1(N__53536),
            .in2(N__43936),
            .in3(N__43891),
            .lcout(buf_adcdata2_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51273),
            .ce(),
            .sr(_gnd_net_));
    defparam i9641_2_lut_3_lut_LC_19_12_2.C_ON=1'b0;
    defparam i9641_2_lut_3_lut_LC_19_12_2.SEQ_MODE=4'b0000;
    defparam i9641_2_lut_3_lut_LC_19_12_2.LUT_INIT=16'b0000000000100010;
    LogicCell40 i9641_2_lut_3_lut_LC_19_12_2 (
            .in0(N__44764),
            .in1(N__50107),
            .in2(_gnd_net_),
            .in3(N__49446),
            .lcout(n14_adj_1215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i27_LC_19_12_3 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i27_LC_19_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i27_LC_19_12_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i27_LC_19_12_3  (
            .in0(N__46116),
            .in1(N__53537),
            .in2(N__43873),
            .in3(N__43890),
            .lcout(cmd_rdadctmp_27_adj_1049),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51273),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i28_LC_19_12_4 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i28_LC_19_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i28_LC_19_12_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i28_LC_19_12_4  (
            .in0(N__53535),
            .in1(N__43869),
            .in2(N__45730),
            .in3(N__46117),
            .lcout(cmd_rdadctmp_28_adj_1048),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51273),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i29_LC_19_12_5 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i29_LC_19_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i29_LC_19_12_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i29_LC_19_12_5  (
            .in0(N__46118),
            .in1(N__45726),
            .in2(N__46357),
            .in3(N__53538),
            .lcout(cmd_rdadctmp_29_adj_1047),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51273),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i30_LC_19_12_7 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i30_LC_19_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i30_LC_19_12_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i30_LC_19_12_7  (
            .in0(N__46119),
            .in1(N__53539),
            .in2(N__48202),
            .in3(N__46353),
            .lcout(cmd_rdadctmp_30_adj_1046),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51273),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_286_LC_19_13_0.C_ON=1'b0;
    defparam i1_2_lut_adj_286_LC_19_13_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_286_LC_19_13_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_286_LC_19_13_0 (
            .in0(_gnd_net_),
            .in1(N__50092),
            .in2(_gnd_net_),
            .in3(N__50593),
            .lcout(n4_adj_1250),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i12_LC_19_13_6 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i12_LC_19_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i12_LC_19_13_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i12_LC_19_13_6  (
            .in0(N__53811),
            .in1(N__45676),
            .in2(N__46145),
            .in3(N__53525),
            .lcout(buf_adcdata2_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51286),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_i9_2_lut_3_lut_LC_19_13_7.C_ON=1'b0;
    defparam comm_cmd_6__I_0_i9_2_lut_3_lut_LC_19_13_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_i9_2_lut_3_lut_LC_19_13_7.LUT_INIT=16'b1101110111111111;
    LogicCell40 comm_cmd_6__I_0_i9_2_lut_3_lut_LC_19_13_7 (
            .in0(N__47605),
            .in1(N__45500),
            .in2(_gnd_net_),
            .in3(N__45152),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i3_LC_19_14_7.C_ON=1'b0;
    defparam comm_buf_1__i3_LC_19_14_7.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i3_LC_19_14_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i3_LC_19_14_7 (
            .in0(N__44884),
            .in1(N__50109),
            .in2(_gnd_net_),
            .in3(N__44786),
            .lcout(comm_buf_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51297),
            .ce(N__44716),
            .sr(N__44657));
    defparam \ADC_VAC1.ADC_DATA_i13_LC_19_15_0 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i13_LC_19_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i13_LC_19_15_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC1.ADC_DATA_i13_LC_19_15_0  (
            .in0(N__52894),
            .in1(N__53129),
            .in2(N__44567),
            .in3(N__44603),
            .lcout(buf_adcdata1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51304),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i18_LC_19_15_4 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i18_LC_19_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i18_LC_19_15_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i18_LC_19_15_4  (
            .in0(N__49213),
            .in1(N__44542),
            .in2(N__44508),
            .in3(N__48830),
            .lcout(cmd_rdadctmp_18_adj_1094),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51304),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i13_LC_19_15_6 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i13_LC_19_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i13_LC_19_15_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i13_LC_19_15_6  (
            .in0(N__53799),
            .in1(N__44485),
            .in2(N__45908),
            .in3(N__53527),
            .lcout(buf_adcdata2_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51304),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i12_LC_19_15_7 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i12_LC_19_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i12_LC_19_15_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i12_LC_19_15_7  (
            .in0(N__53128),
            .in1(N__46252),
            .in2(N__46292),
            .in3(N__52895),
            .lcout(buf_adcdata1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51304),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i9_LC_19_16_0 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i9_LC_19_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i9_LC_19_16_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i9_LC_19_16_0  (
            .in0(N__53798),
            .in1(N__46195),
            .in2(N__46238),
            .in3(N__53572),
            .lcout(buf_adcdata2_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51310),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i20_LC_19_16_4 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i20_LC_19_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i20_LC_19_16_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i20_LC_19_16_4  (
            .in0(N__46177),
            .in1(N__46108),
            .in2(N__46141),
            .in3(N__53573),
            .lcout(cmd_rdadctmp_20_adj_1056),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51310),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i21_LC_19_16_5 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i21_LC_19_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i21_LC_19_16_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i21_LC_19_16_5  (
            .in0(N__53570),
            .in1(N__46137),
            .in2(N__46120),
            .in3(N__45903),
            .lcout(cmd_rdadctmp_21_adj_1055),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51310),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.cmd_rdadctmp_i22_LC_19_16_7 .C_ON=1'b0;
    defparam \ADC_VAC2.cmd_rdadctmp_i22_LC_19_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.cmd_rdadctmp_i22_LC_19_16_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_VAC2.cmd_rdadctmp_i22_LC_19_16_7  (
            .in0(N__53571),
            .in1(N__53592),
            .in2(N__46121),
            .in3(N__45904),
            .lcout(cmd_rdadctmp_22_adj_1054),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51310),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1469_i8_4_lut_LC_20_3_4.C_ON=1'b0;
    defparam mux_1469_i8_4_lut_LC_20_3_4.SEQ_MODE=4'b0000;
    defparam mux_1469_i8_4_lut_LC_20_3_4.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1469_i8_4_lut_LC_20_3_4 (
            .in0(N__45890),
            .in1(N__47929),
            .in2(N__45877),
            .in3(N__47267),
            .lcout(n4101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_7330_7331_reset_LC_20_5_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_7330_7331_reset_LC_20_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imosi_44_7330_7331_reset_LC_20_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_7330_7331_reset_LC_20_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45777),
            .lcout(\comm_spi.n10442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51173),
            .ce(),
            .sr(N__45740));
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_20_6_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_20_6_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_20_6_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_89_2_lut_LC_20_6_4  (
            .in0(N__45794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46470),
            .lcout(\comm_spi.imosi_N_792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i20_LC_20_6_6 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i20_LC_20_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i20_LC_20_6_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i20_LC_20_6_6  (
            .in0(N__53733),
            .in1(N__45703),
            .in2(N__45734),
            .in3(N__53532),
            .lcout(buf_adcdata2_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51191),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i23_LC_20_6_7 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i23_LC_20_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i23_LC_20_6_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i23_LC_20_6_7  (
            .in0(N__53531),
            .in1(N__53734),
            .in2(N__48158),
            .in3(N__48118),
            .lcout(buf_adcdata2_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51191),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_1469_i1_4_lut_LC_20_7_0.C_ON=1'b0;
    defparam mux_1469_i1_4_lut_LC_20_7_0.SEQ_MODE=4'b0000;
    defparam mux_1469_i1_4_lut_LC_20_7_0.LUT_INIT=16'b1010101000110000;
    LogicCell40 mux_1469_i1_4_lut_LC_20_7_0 (
            .in0(N__48104),
            .in1(N__47854),
            .in2(N__47378),
            .in3(N__47094),
            .lcout(n4108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i2_LC_20_7_3 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i2_LC_20_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i2_LC_20_7_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i2_LC_20_7_3  (
            .in0(N__53754),
            .in1(N__46667),
            .in2(N__46706),
            .in3(N__53575),
            .lcout(buf_adcdata2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51208),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_20_7_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_20_7_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_20_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_95_2_lut_LC_20_7_4  (
            .in0(N__46638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46501),
            .lcout(\comm_spi.data_tx_7__N_808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_20_7_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_20_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_90_2_lut_LC_20_7_5  (
            .in0(N__51374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46469),
            .lcout(\comm_spi.iclk_N_801 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i13102_4_lut_3_lut_LC_20_7_6 .C_ON=1'b0;
    defparam \comm_spi.i13102_4_lut_3_lut_LC_20_7_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i13102_4_lut_3_lut_LC_20_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.i13102_4_lut_3_lut_LC_20_7_6  (
            .in0(N__46639),
            .in1(N__46502),
            .in2(_gnd_net_),
            .in3(N__46377),
            .lcout(\comm_spi.n16899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i21_LC_20_7_7 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i21_LC_20_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i21_LC_20_7_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i21_LC_20_7_7  (
            .in0(N__53753),
            .in1(N__46327),
            .in2(N__46361),
            .in3(N__53574),
            .lcout(buf_adcdata2_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51208),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_response_331_LC_20_8_0.C_ON=1'b0;
    defparam comm_response_331_LC_20_8_0.SEQ_MODE=4'b1000;
    defparam comm_response_331_LC_20_8_0.LUT_INIT=16'b0001000000011010;
    LogicCell40 comm_response_331_LC_20_8_0 (
            .in0(N__50141),
            .in1(N__49406),
            .in2(N__52356),
            .in3(N__50554),
            .lcout(ICE_GPMI_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51225),
            .ce(N__49298),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_4_lut_LC_20_8_3.C_ON=1'b0;
    defparam i1_4_lut_4_lut_4_lut_LC_20_8_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_4_lut_LC_20_8_3.LUT_INIT=16'b1100110111000010;
    LogicCell40 i1_4_lut_4_lut_4_lut_LC_20_8_3 (
            .in0(N__50552),
            .in1(N__52220),
            .in2(N__50292),
            .in3(N__49436),
            .lcout(n8576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_20_8_5.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_20_8_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_20_8_5.LUT_INIT=16'b1111101111111011;
    LogicCell40 i2_2_lut_3_lut_LC_20_8_5 (
            .in0(N__50553),
            .in1(N__52221),
            .in2(N__50293),
            .in3(_gnd_net_),
            .lcout(n8117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_adj_226_LC_20_8_6.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_226_LC_20_8_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_226_LC_20_8_6.LUT_INIT=16'b1110111011111111;
    LogicCell40 i2_2_lut_3_lut_adj_226_LC_20_8_6 (
            .in0(N__52219),
            .in1(N__49405),
            .in2(_gnd_net_),
            .in3(N__50551),
            .lcout(n6_adj_1175),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_4_lut_LC_20_9_1.C_ON=1'b0;
    defparam i1_3_lut_4_lut_4_lut_LC_20_9_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_4_lut_LC_20_9_1.LUT_INIT=16'b1111000011101111;
    LogicCell40 i1_3_lut_4_lut_4_lut_LC_20_9_1 (
            .in0(N__50595),
            .in1(N__50142),
            .in2(N__52390),
            .in3(N__49437),
            .lcout(n8129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC3.cmd_rdadctmp_i20_LC_20_9_5 .C_ON=1'b0;
    defparam \ADC_VAC3.cmd_rdadctmp_i20_LC_20_9_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC3.cmd_rdadctmp_i20_LC_20_9_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC3.cmd_rdadctmp_i20_LC_20_9_5  (
            .in0(N__49285),
            .in1(N__49242),
            .in2(N__48589),
            .in3(N__48841),
            .lcout(cmd_rdadctmp_20_adj_1092),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51243),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLOCK_DDS.dds_state_i0_LC_20_10_0 .C_ON=1'b0;
    defparam \CLOCK_DDS.dds_state_i0_LC_20_10_0 .SEQ_MODE=4'b1000;
    defparam \CLOCK_DDS.dds_state_i0_LC_20_10_0 .LUT_INIT=16'b1010000000110011;
    LogicCell40 \CLOCK_DDS.dds_state_i0_LC_20_10_0  (
            .in0(N__48572),
            .in1(N__48334),
            .in2(N__48563),
            .in3(N__48542),
            .lcout(dds_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51258),
            .ce(N__48298),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i16_LC_20_11_5 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i16_LC_20_11_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i16_LC_20_11_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i16_LC_20_11_5  (
            .in0(N__53117),
            .in1(N__48226),
            .in2(N__48272),
            .in3(N__52893),
            .lcout(buf_adcdata1_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51274),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i22_LC_20_11_6 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i22_LC_20_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i22_LC_20_11_6 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \ADC_VAC2.ADC_DATA_i22_LC_20_11_6  (
            .in0(N__48201),
            .in1(N__53775),
            .in2(N__53576),
            .in3(N__48172),
            .lcout(buf_adcdata2_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51274),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC2.ADC_DATA_i14_LC_20_13_5 .C_ON=1'b0;
    defparam \ADC_VAC2.ADC_DATA_i14_LC_20_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC2.ADC_DATA_i14_LC_20_13_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC2.ADC_DATA_i14_LC_20_13_5  (
            .in0(N__53812),
            .in1(N__53143),
            .in2(N__53609),
            .in3(N__53526),
            .lcout(buf_adcdata2_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51298),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC1.ADC_DATA_i10_LC_20_17_3 .C_ON=1'b0;
    defparam \ADC_VAC1.ADC_DATA_i10_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC1.ADC_DATA_i10_LC_20_17_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_VAC1.ADC_DATA_i10_LC_20_17_3  (
            .in0(N__53114),
            .in1(N__52504),
            .in2(N__52934),
            .in3(N__52896),
            .lcout(buf_adcdata1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51316),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_394_Mux_5_i15_4_lut_LC_20_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_394_Mux_5_i15_4_lut_LC_20_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_394_Mux_5_i15_4_lut_LC_20_19_4.LUT_INIT=16'b0011101100001000;
    LogicCell40 comm_state_3__I_0_394_Mux_5_i15_4_lut_LC_20_19_4 (
            .in0(N__52490),
            .in1(N__52455),
            .in2(N__51932),
            .in3(N__51515),
            .lcout(data_index_9_N_258_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_7326_7327_set_LC_23_7_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_7326_7327_set_LC_23_7_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.iclk_40_7326_7327_set_LC_23_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_7326_7327_set_LC_23_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51375),
            .lcout(\comm_spi.n10437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51261),
            .ce(),
            .sr(N__50672));
endmodule // zimaux
