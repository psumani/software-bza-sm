-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 3 2023 14:37:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "zim" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of zim
entity zim is
port (
    VAC_DRDY : in std_logic;
    IAC_FLT1 : out std_logic;
    DDS_SCK : out std_logic;
    ICE_IOR_166 : in std_logic;
    ICE_IOR_119 : in std_logic;
    DDS_MOSI : out std_logic;
    VAC_MISO : in std_logic;
    DDS_MOSI1 : out std_logic;
    ICE_IOR_146 : in std_logic;
    VDC_CLK : out std_logic;
    ICE_IOT_222 : in std_logic;
    IAC_CS : out std_logic;
    ICE_IOL_18B : in std_logic;
    ICE_IOL_13A : in std_logic;
    ICE_IOB_81 : in std_logic;
    VAC_OSR1 : out std_logic;
    IAC_MOSI : out std_logic;
    DDS_CS1 : out std_logic;
    ICE_IOL_4B : in std_logic;
    ICE_IOB_94 : in std_logic;
    VAC_CS : out std_logic;
    VAC_CLK : out std_logic;
    ICE_SPI_CE0 : in std_logic;
    ICE_IOR_167 : in std_logic;
    ICE_IOR_118 : in std_logic;
    RTD_SDO : in std_logic;
    IAC_OSR0 : out std_logic;
    VDC_SCLK : out std_logic;
    VAC_FLT1 : out std_logic;
    ICE_SPI_MOSI : in std_logic;
    ICE_IOR_165 : in std_logic;
    ICE_IOR_147 : in std_logic;
    ICE_IOL_14A : in std_logic;
    ICE_IOL_13B : in std_logic;
    ICE_IOB_91 : in std_logic;
    ICE_GPMO_0 : in std_logic;
    DDS_RNG_0 : out std_logic;
    VDC_RNG0 : out std_logic;
    ICE_SPI_SCLK : in std_logic;
    ICE_IOR_152 : in std_logic;
    ICE_IOL_12A : in std_logic;
    RTD_DRDY : in std_logic;
    ICE_SPI_MISO : out std_logic;
    ICE_IOT_177 : in std_logic;
    ICE_IOR_141 : in std_logic;
    ICE_IOB_80 : in std_logic;
    ICE_IOB_102 : in std_logic;
    ICE_GPMO_2 : in std_logic;
    ICE_GPMI_0 : out std_logic;
    IAC_MISO : in std_logic;
    VAC_OSR0 : out std_logic;
    VAC_MOSI : out std_logic;
    TEST_LED : out std_logic;
    ICE_IOR_148 : in std_logic;
    STAT_COMM : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_IOR_161 : in std_logic;
    ICE_IOB_95 : in std_logic;
    ICE_IOB_82 : in std_logic;
    ICE_IOB_104 : in std_logic;
    IAC_CLK : out std_logic;
    DDS_CS : out std_logic;
    SELIRNG0 : out std_logic;
    RTD_SDI : out std_logic;
    ICE_IOT_221 : in std_logic;
    ICE_IOT_197 : in std_logic;
    DDS_MCLK : out std_logic;
    RTD_SCLK : out std_logic;
    RTD_CS : out std_logic;
    ICE_IOR_137 : in std_logic;
    IAC_OSR1 : out std_logic;
    VAC_FLT0 : out std_logic;
    ICE_IOR_144 : in std_logic;
    ICE_IOR_128 : in std_logic;
    ICE_GPMO_1 : in std_logic;
    IAC_SCLK : out std_logic;
    EIS_SYNCCLK : in std_logic;
    ICE_IOR_139 : in std_logic;
    ICE_IOL_4A : in std_logic;
    VAC_SCLK : out std_logic;
    THERMOSTAT : in std_logic;
    ICE_IOR_164 : in std_logic;
    ICE_IOB_103 : in std_logic;
    AMPV_POW : out std_logic;
    VDC_SDO : in std_logic;
    ICE_IOT_174 : in std_logic;
    ICE_IOR_140 : in std_logic;
    ICE_IOB_96 : in std_logic;
    CONT_SD : out std_logic;
    AC_ADC_SYNC : out std_logic;
    SELIRNG1 : out std_logic;
    ICE_IOL_12B : in std_logic;
    ICE_IOR_160 : in std_logic;
    ICE_IOR_136 : in std_logic;
    DDS_MCLK1 : out std_logic;
    ICE_IOT_198 : in std_logic;
    ICE_IOT_173 : in std_logic;
    IAC_DRDY : in std_logic;
    ICE_IOT_178 : in std_logic;
    ICE_IOR_138 : in std_logic;
    ICE_IOR_120 : in std_logic;
    IAC_FLT0 : out std_logic;
    DDS_SCK1 : out std_logic);
end zim;

-- Architecture of zim
-- View name is \INTERFACE\
architecture \INTERFACE\ of zim is

signal \N__59563\ : std_logic;
signal \N__59562\ : std_logic;
signal \N__59561\ : std_logic;
signal \N__59554\ : std_logic;
signal \N__59553\ : std_logic;
signal \N__59552\ : std_logic;
signal \N__59545\ : std_logic;
signal \N__59544\ : std_logic;
signal \N__59543\ : std_logic;
signal \N__59536\ : std_logic;
signal \N__59535\ : std_logic;
signal \N__59534\ : std_logic;
signal \N__59527\ : std_logic;
signal \N__59526\ : std_logic;
signal \N__59525\ : std_logic;
signal \N__59518\ : std_logic;
signal \N__59517\ : std_logic;
signal \N__59516\ : std_logic;
signal \N__59509\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59507\ : std_logic;
signal \N__59500\ : std_logic;
signal \N__59499\ : std_logic;
signal \N__59498\ : std_logic;
signal \N__59491\ : std_logic;
signal \N__59490\ : std_logic;
signal \N__59489\ : std_logic;
signal \N__59482\ : std_logic;
signal \N__59481\ : std_logic;
signal \N__59480\ : std_logic;
signal \N__59473\ : std_logic;
signal \N__59472\ : std_logic;
signal \N__59471\ : std_logic;
signal \N__59464\ : std_logic;
signal \N__59463\ : std_logic;
signal \N__59462\ : std_logic;
signal \N__59455\ : std_logic;
signal \N__59454\ : std_logic;
signal \N__59453\ : std_logic;
signal \N__59446\ : std_logic;
signal \N__59445\ : std_logic;
signal \N__59444\ : std_logic;
signal \N__59437\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59435\ : std_logic;
signal \N__59428\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59426\ : std_logic;
signal \N__59419\ : std_logic;
signal \N__59418\ : std_logic;
signal \N__59417\ : std_logic;
signal \N__59410\ : std_logic;
signal \N__59409\ : std_logic;
signal \N__59408\ : std_logic;
signal \N__59401\ : std_logic;
signal \N__59400\ : std_logic;
signal \N__59399\ : std_logic;
signal \N__59392\ : std_logic;
signal \N__59391\ : std_logic;
signal \N__59390\ : std_logic;
signal \N__59383\ : std_logic;
signal \N__59382\ : std_logic;
signal \N__59381\ : std_logic;
signal \N__59374\ : std_logic;
signal \N__59373\ : std_logic;
signal \N__59372\ : std_logic;
signal \N__59365\ : std_logic;
signal \N__59364\ : std_logic;
signal \N__59363\ : std_logic;
signal \N__59356\ : std_logic;
signal \N__59355\ : std_logic;
signal \N__59354\ : std_logic;
signal \N__59347\ : std_logic;
signal \N__59346\ : std_logic;
signal \N__59345\ : std_logic;
signal \N__59338\ : std_logic;
signal \N__59337\ : std_logic;
signal \N__59336\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59328\ : std_logic;
signal \N__59327\ : std_logic;
signal \N__59320\ : std_logic;
signal \N__59319\ : std_logic;
signal \N__59318\ : std_logic;
signal \N__59311\ : std_logic;
signal \N__59310\ : std_logic;
signal \N__59309\ : std_logic;
signal \N__59302\ : std_logic;
signal \N__59301\ : std_logic;
signal \N__59300\ : std_logic;
signal \N__59293\ : std_logic;
signal \N__59292\ : std_logic;
signal \N__59291\ : std_logic;
signal \N__59284\ : std_logic;
signal \N__59283\ : std_logic;
signal \N__59282\ : std_logic;
signal \N__59275\ : std_logic;
signal \N__59274\ : std_logic;
signal \N__59273\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59265\ : std_logic;
signal \N__59264\ : std_logic;
signal \N__59257\ : std_logic;
signal \N__59256\ : std_logic;
signal \N__59255\ : std_logic;
signal \N__59248\ : std_logic;
signal \N__59247\ : std_logic;
signal \N__59246\ : std_logic;
signal \N__59239\ : std_logic;
signal \N__59238\ : std_logic;
signal \N__59237\ : std_logic;
signal \N__59230\ : std_logic;
signal \N__59229\ : std_logic;
signal \N__59228\ : std_logic;
signal \N__59221\ : std_logic;
signal \N__59220\ : std_logic;
signal \N__59219\ : std_logic;
signal \N__59212\ : std_logic;
signal \N__59211\ : std_logic;
signal \N__59210\ : std_logic;
signal \N__59203\ : std_logic;
signal \N__59202\ : std_logic;
signal \N__59201\ : std_logic;
signal \N__59194\ : std_logic;
signal \N__59193\ : std_logic;
signal \N__59192\ : std_logic;
signal \N__59185\ : std_logic;
signal \N__59184\ : std_logic;
signal \N__59183\ : std_logic;
signal \N__59176\ : std_logic;
signal \N__59175\ : std_logic;
signal \N__59174\ : std_logic;
signal \N__59167\ : std_logic;
signal \N__59166\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59158\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59156\ : std_logic;
signal \N__59149\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59147\ : std_logic;
signal \N__59140\ : std_logic;
signal \N__59139\ : std_logic;
signal \N__59138\ : std_logic;
signal \N__59131\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59129\ : std_logic;
signal \N__59122\ : std_logic;
signal \N__59121\ : std_logic;
signal \N__59120\ : std_logic;
signal \N__59113\ : std_logic;
signal \N__59112\ : std_logic;
signal \N__59111\ : std_logic;
signal \N__59104\ : std_logic;
signal \N__59103\ : std_logic;
signal \N__59102\ : std_logic;
signal \N__59095\ : std_logic;
signal \N__59094\ : std_logic;
signal \N__59093\ : std_logic;
signal \N__59086\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59084\ : std_logic;
signal \N__59077\ : std_logic;
signal \N__59076\ : std_logic;
signal \N__59075\ : std_logic;
signal \N__59068\ : std_logic;
signal \N__59067\ : std_logic;
signal \N__59066\ : std_logic;
signal \N__59059\ : std_logic;
signal \N__59058\ : std_logic;
signal \N__59057\ : std_logic;
signal \N__59050\ : std_logic;
signal \N__59049\ : std_logic;
signal \N__59048\ : std_logic;
signal \N__59041\ : std_logic;
signal \N__59040\ : std_logic;
signal \N__59039\ : std_logic;
signal \N__59032\ : std_logic;
signal \N__59031\ : std_logic;
signal \N__59030\ : std_logic;
signal \N__59023\ : std_logic;
signal \N__59022\ : std_logic;
signal \N__59021\ : std_logic;
signal \N__59014\ : std_logic;
signal \N__59013\ : std_logic;
signal \N__59012\ : std_logic;
signal \N__59005\ : std_logic;
signal \N__59004\ : std_logic;
signal \N__59003\ : std_logic;
signal \N__58996\ : std_logic;
signal \N__58995\ : std_logic;
signal \N__58994\ : std_logic;
signal \N__58987\ : std_logic;
signal \N__58986\ : std_logic;
signal \N__58985\ : std_logic;
signal \N__58978\ : std_logic;
signal \N__58977\ : std_logic;
signal \N__58976\ : std_logic;
signal \N__58969\ : std_logic;
signal \N__58968\ : std_logic;
signal \N__58967\ : std_logic;
signal \N__58960\ : std_logic;
signal \N__58959\ : std_logic;
signal \N__58958\ : std_logic;
signal \N__58951\ : std_logic;
signal \N__58950\ : std_logic;
signal \N__58949\ : std_logic;
signal \N__58942\ : std_logic;
signal \N__58941\ : std_logic;
signal \N__58940\ : std_logic;
signal \N__58933\ : std_logic;
signal \N__58932\ : std_logic;
signal \N__58931\ : std_logic;
signal \N__58924\ : std_logic;
signal \N__58923\ : std_logic;
signal \N__58922\ : std_logic;
signal \N__58915\ : std_logic;
signal \N__58914\ : std_logic;
signal \N__58913\ : std_logic;
signal \N__58906\ : std_logic;
signal \N__58905\ : std_logic;
signal \N__58904\ : std_logic;
signal \N__58897\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58895\ : std_logic;
signal \N__58888\ : std_logic;
signal \N__58887\ : std_logic;
signal \N__58886\ : std_logic;
signal \N__58879\ : std_logic;
signal \N__58878\ : std_logic;
signal \N__58877\ : std_logic;
signal \N__58870\ : std_logic;
signal \N__58869\ : std_logic;
signal \N__58868\ : std_logic;
signal \N__58861\ : std_logic;
signal \N__58860\ : std_logic;
signal \N__58859\ : std_logic;
signal \N__58852\ : std_logic;
signal \N__58851\ : std_logic;
signal \N__58850\ : std_logic;
signal \N__58843\ : std_logic;
signal \N__58842\ : std_logic;
signal \N__58841\ : std_logic;
signal \N__58834\ : std_logic;
signal \N__58833\ : std_logic;
signal \N__58832\ : std_logic;
signal \N__58825\ : std_logic;
signal \N__58824\ : std_logic;
signal \N__58823\ : std_logic;
signal \N__58816\ : std_logic;
signal \N__58815\ : std_logic;
signal \N__58814\ : std_logic;
signal \N__58807\ : std_logic;
signal \N__58806\ : std_logic;
signal \N__58805\ : std_logic;
signal \N__58798\ : std_logic;
signal \N__58797\ : std_logic;
signal \N__58796\ : std_logic;
signal \N__58789\ : std_logic;
signal \N__58788\ : std_logic;
signal \N__58787\ : std_logic;
signal \N__58780\ : std_logic;
signal \N__58779\ : std_logic;
signal \N__58778\ : std_logic;
signal \N__58771\ : std_logic;
signal \N__58770\ : std_logic;
signal \N__58769\ : std_logic;
signal \N__58762\ : std_logic;
signal \N__58761\ : std_logic;
signal \N__58760\ : std_logic;
signal \N__58753\ : std_logic;
signal \N__58752\ : std_logic;
signal \N__58751\ : std_logic;
signal \N__58744\ : std_logic;
signal \N__58743\ : std_logic;
signal \N__58742\ : std_logic;
signal \N__58735\ : std_logic;
signal \N__58734\ : std_logic;
signal \N__58733\ : std_logic;
signal \N__58726\ : std_logic;
signal \N__58725\ : std_logic;
signal \N__58724\ : std_logic;
signal \N__58717\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58715\ : std_logic;
signal \N__58708\ : std_logic;
signal \N__58707\ : std_logic;
signal \N__58706\ : std_logic;
signal \N__58699\ : std_logic;
signal \N__58698\ : std_logic;
signal \N__58697\ : std_logic;
signal \N__58690\ : std_logic;
signal \N__58689\ : std_logic;
signal \N__58688\ : std_logic;
signal \N__58681\ : std_logic;
signal \N__58680\ : std_logic;
signal \N__58679\ : std_logic;
signal \N__58672\ : std_logic;
signal \N__58671\ : std_logic;
signal \N__58670\ : std_logic;
signal \N__58663\ : std_logic;
signal \N__58662\ : std_logic;
signal \N__58661\ : std_logic;
signal \N__58654\ : std_logic;
signal \N__58653\ : std_logic;
signal \N__58652\ : std_logic;
signal \N__58645\ : std_logic;
signal \N__58644\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58626\ : std_logic;
signal \N__58623\ : std_logic;
signal \N__58622\ : std_logic;
signal \N__58621\ : std_logic;
signal \N__58620\ : std_logic;
signal \N__58617\ : std_logic;
signal \N__58616\ : std_logic;
signal \N__58613\ : std_logic;
signal \N__58612\ : std_logic;
signal \N__58609\ : std_logic;
signal \N__58608\ : std_logic;
signal \N__58607\ : std_logic;
signal \N__58592\ : std_logic;
signal \N__58589\ : std_logic;
signal \N__58586\ : std_logic;
signal \N__58585\ : std_logic;
signal \N__58584\ : std_logic;
signal \N__58581\ : std_logic;
signal \N__58580\ : std_logic;
signal \N__58579\ : std_logic;
signal \N__58578\ : std_logic;
signal \N__58577\ : std_logic;
signal \N__58576\ : std_logic;
signal \N__58575\ : std_logic;
signal \N__58574\ : std_logic;
signal \N__58573\ : std_logic;
signal \N__58570\ : std_logic;
signal \N__58567\ : std_logic;
signal \N__58566\ : std_logic;
signal \N__58565\ : std_logic;
signal \N__58564\ : std_logic;
signal \N__58561\ : std_logic;
signal \N__58560\ : std_logic;
signal \N__58557\ : std_logic;
signal \N__58554\ : std_logic;
signal \N__58553\ : std_logic;
signal \N__58550\ : std_logic;
signal \N__58549\ : std_logic;
signal \N__58546\ : std_logic;
signal \N__58545\ : std_logic;
signal \N__58542\ : std_logic;
signal \N__58541\ : std_logic;
signal \N__58538\ : std_logic;
signal \N__58537\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58533\ : std_logic;
signal \N__58530\ : std_logic;
signal \N__58529\ : std_logic;
signal \N__58526\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58524\ : std_logic;
signal \N__58523\ : std_logic;
signal \N__58522\ : std_logic;
signal \N__58519\ : std_logic;
signal \N__58516\ : std_logic;
signal \N__58513\ : std_logic;
signal \N__58510\ : std_logic;
signal \N__58509\ : std_logic;
signal \N__58508\ : std_logic;
signal \N__58507\ : std_logic;
signal \N__58504\ : std_logic;
signal \N__58503\ : std_logic;
signal \N__58502\ : std_logic;
signal \N__58501\ : std_logic;
signal \N__58500\ : std_logic;
signal \N__58497\ : std_logic;
signal \N__58494\ : std_logic;
signal \N__58491\ : std_logic;
signal \N__58476\ : std_logic;
signal \N__58459\ : std_logic;
signal \N__58456\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58451\ : std_logic;
signal \N__58448\ : std_logic;
signal \N__58447\ : std_logic;
signal \N__58444\ : std_logic;
signal \N__58435\ : std_logic;
signal \N__58432\ : std_logic;
signal \N__58429\ : std_logic;
signal \N__58428\ : std_logic;
signal \N__58425\ : std_logic;
signal \N__58424\ : std_logic;
signal \N__58421\ : std_logic;
signal \N__58420\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58416\ : std_logic;
signal \N__58413\ : std_logic;
signal \N__58412\ : std_logic;
signal \N__58409\ : std_logic;
signal \N__58408\ : std_logic;
signal \N__58405\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58397\ : std_logic;
signal \N__58394\ : std_logic;
signal \N__58391\ : std_logic;
signal \N__58376\ : std_logic;
signal \N__58369\ : std_logic;
signal \N__58366\ : std_logic;
signal \N__58363\ : std_logic;
signal \N__58360\ : std_logic;
signal \N__58359\ : std_logic;
signal \N__58356\ : std_logic;
signal \N__58339\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58335\ : std_logic;
signal \N__58326\ : std_logic;
signal \N__58317\ : std_logic;
signal \N__58314\ : std_logic;
signal \N__58311\ : std_logic;
signal \N__58308\ : std_logic;
signal \N__58305\ : std_logic;
signal \N__58302\ : std_logic;
signal \N__58299\ : std_logic;
signal \N__58294\ : std_logic;
signal \N__58293\ : std_logic;
signal \N__58288\ : std_logic;
signal \N__58283\ : std_logic;
signal \N__58278\ : std_logic;
signal \N__58275\ : std_logic;
signal \N__58266\ : std_logic;
signal \N__58263\ : std_logic;
signal \N__58260\ : std_logic;
signal \N__58259\ : std_logic;
signal \N__58258\ : std_logic;
signal \N__58255\ : std_logic;
signal \N__58252\ : std_logic;
signal \N__58249\ : std_logic;
signal \N__58244\ : std_logic;
signal \N__58243\ : std_logic;
signal \N__58240\ : std_logic;
signal \N__58237\ : std_logic;
signal \N__58234\ : std_logic;
signal \N__58231\ : std_logic;
signal \N__58226\ : std_logic;
signal \N__58221\ : std_logic;
signal \N__58218\ : std_logic;
signal \N__58217\ : std_logic;
signal \N__58214\ : std_logic;
signal \N__58211\ : std_logic;
signal \N__58206\ : std_logic;
signal \N__58205\ : std_logic;
signal \N__58202\ : std_logic;
signal \N__58199\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58193\ : std_logic;
signal \N__58190\ : std_logic;
signal \N__58187\ : std_logic;
signal \N__58184\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58176\ : std_logic;
signal \N__58175\ : std_logic;
signal \N__58172\ : std_logic;
signal \N__58169\ : std_logic;
signal \N__58164\ : std_logic;
signal \N__58161\ : std_logic;
signal \N__58160\ : std_logic;
signal \N__58157\ : std_logic;
signal \N__58154\ : std_logic;
signal \N__58151\ : std_logic;
signal \N__58148\ : std_logic;
signal \N__58145\ : std_logic;
signal \N__58142\ : std_logic;
signal \N__58139\ : std_logic;
signal \N__58136\ : std_logic;
signal \N__58131\ : std_logic;
signal \N__58130\ : std_logic;
signal \N__58127\ : std_logic;
signal \N__58124\ : std_logic;
signal \N__58119\ : std_logic;
signal \N__58116\ : std_logic;
signal \N__58115\ : std_logic;
signal \N__58112\ : std_logic;
signal \N__58109\ : std_logic;
signal \N__58104\ : std_logic;
signal \N__58103\ : std_logic;
signal \N__58100\ : std_logic;
signal \N__58097\ : std_logic;
signal \N__58094\ : std_logic;
signal \N__58089\ : std_logic;
signal \N__58088\ : std_logic;
signal \N__58085\ : std_logic;
signal \N__58082\ : std_logic;
signal \N__58077\ : std_logic;
signal \N__58074\ : std_logic;
signal \N__58071\ : std_logic;
signal \N__58070\ : std_logic;
signal \N__58067\ : std_logic;
signal \N__58064\ : std_logic;
signal \N__58059\ : std_logic;
signal \N__58056\ : std_logic;
signal \N__58055\ : std_logic;
signal \N__58052\ : std_logic;
signal \N__58049\ : std_logic;
signal \N__58044\ : std_logic;
signal \N__58043\ : std_logic;
signal \N__58040\ : std_logic;
signal \N__58037\ : std_logic;
signal \N__58034\ : std_logic;
signal \N__58029\ : std_logic;
signal \N__58028\ : std_logic;
signal \N__58025\ : std_logic;
signal \N__58022\ : std_logic;
signal \N__58017\ : std_logic;
signal \N__58014\ : std_logic;
signal \N__58011\ : std_logic;
signal \N__58010\ : std_logic;
signal \N__58007\ : std_logic;
signal \N__58006\ : std_logic;
signal \N__58005\ : std_logic;
signal \N__58004\ : std_logic;
signal \N__58003\ : std_logic;
signal \N__58002\ : std_logic;
signal \N__57999\ : std_logic;
signal \N__57996\ : std_logic;
signal \N__57993\ : std_logic;
signal \N__57986\ : std_logic;
signal \N__57983\ : std_logic;
signal \N__57978\ : std_logic;
signal \N__57975\ : std_logic;
signal \N__57972\ : std_logic;
signal \N__57963\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57959\ : std_logic;
signal \N__57956\ : std_logic;
signal \N__57953\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57947\ : std_logic;
signal \N__57944\ : std_logic;
signal \N__57941\ : std_logic;
signal \N__57936\ : std_logic;
signal \N__57935\ : std_logic;
signal \N__57932\ : std_logic;
signal \N__57929\ : std_logic;
signal \N__57924\ : std_logic;
signal \N__57921\ : std_logic;
signal \N__57920\ : std_logic;
signal \N__57917\ : std_logic;
signal \N__57914\ : std_logic;
signal \N__57909\ : std_logic;
signal \N__57908\ : std_logic;
signal \N__57905\ : std_logic;
signal \N__57902\ : std_logic;
signal \N__57899\ : std_logic;
signal \N__57894\ : std_logic;
signal \N__57891\ : std_logic;
signal \N__57890\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57884\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57876\ : std_logic;
signal \N__57873\ : std_logic;
signal \N__57870\ : std_logic;
signal \N__57867\ : std_logic;
signal \N__57864\ : std_logic;
signal \N__57861\ : std_logic;
signal \N__57858\ : std_logic;
signal \N__57855\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57843\ : std_logic;
signal \N__57840\ : std_logic;
signal \N__57837\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57831\ : std_logic;
signal \N__57828\ : std_logic;
signal \N__57825\ : std_logic;
signal \N__57824\ : std_logic;
signal \N__57823\ : std_logic;
signal \N__57822\ : std_logic;
signal \N__57821\ : std_logic;
signal \N__57820\ : std_logic;
signal \N__57819\ : std_logic;
signal \N__57818\ : std_logic;
signal \N__57817\ : std_logic;
signal \N__57816\ : std_logic;
signal \N__57815\ : std_logic;
signal \N__57814\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57812\ : std_logic;
signal \N__57809\ : std_logic;
signal \N__57808\ : std_logic;
signal \N__57807\ : std_logic;
signal \N__57806\ : std_logic;
signal \N__57805\ : std_logic;
signal \N__57804\ : std_logic;
signal \N__57803\ : std_logic;
signal \N__57802\ : std_logic;
signal \N__57801\ : std_logic;
signal \N__57800\ : std_logic;
signal \N__57797\ : std_logic;
signal \N__57796\ : std_logic;
signal \N__57795\ : std_logic;
signal \N__57794\ : std_logic;
signal \N__57793\ : std_logic;
signal \N__57792\ : std_logic;
signal \N__57789\ : std_logic;
signal \N__57788\ : std_logic;
signal \N__57787\ : std_logic;
signal \N__57786\ : std_logic;
signal \N__57785\ : std_logic;
signal \N__57784\ : std_logic;
signal \N__57783\ : std_logic;
signal \N__57782\ : std_logic;
signal \N__57781\ : std_logic;
signal \N__57780\ : std_logic;
signal \N__57779\ : std_logic;
signal \N__57778\ : std_logic;
signal \N__57777\ : std_logic;
signal \N__57776\ : std_logic;
signal \N__57773\ : std_logic;
signal \N__57770\ : std_logic;
signal \N__57767\ : std_logic;
signal \N__57764\ : std_logic;
signal \N__57763\ : std_logic;
signal \N__57760\ : std_logic;
signal \N__57759\ : std_logic;
signal \N__57758\ : std_logic;
signal \N__57757\ : std_logic;
signal \N__57756\ : std_logic;
signal \N__57755\ : std_logic;
signal \N__57754\ : std_logic;
signal \N__57751\ : std_logic;
signal \N__57750\ : std_logic;
signal \N__57749\ : std_logic;
signal \N__57748\ : std_logic;
signal \N__57747\ : std_logic;
signal \N__57744\ : std_logic;
signal \N__57741\ : std_logic;
signal \N__57740\ : std_logic;
signal \N__57739\ : std_logic;
signal \N__57738\ : std_logic;
signal \N__57737\ : std_logic;
signal \N__57736\ : std_logic;
signal \N__57729\ : std_logic;
signal \N__57724\ : std_logic;
signal \N__57717\ : std_logic;
signal \N__57714\ : std_logic;
signal \N__57705\ : std_logic;
signal \N__57702\ : std_logic;
signal \N__57701\ : std_logic;
signal \N__57700\ : std_logic;
signal \N__57699\ : std_logic;
signal \N__57698\ : std_logic;
signal \N__57695\ : std_logic;
signal \N__57690\ : std_logic;
signal \N__57685\ : std_logic;
signal \N__57682\ : std_logic;
signal \N__57675\ : std_logic;
signal \N__57672\ : std_logic;
signal \N__57669\ : std_logic;
signal \N__57668\ : std_logic;
signal \N__57667\ : std_logic;
signal \N__57666\ : std_logic;
signal \N__57665\ : std_logic;
signal \N__57662\ : std_logic;
signal \N__57661\ : std_logic;
signal \N__57658\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57654\ : std_logic;
signal \N__57653\ : std_logic;
signal \N__57652\ : std_logic;
signal \N__57651\ : std_logic;
signal \N__57648\ : std_logic;
signal \N__57643\ : std_logic;
signal \N__57642\ : std_logic;
signal \N__57641\ : std_logic;
signal \N__57638\ : std_logic;
signal \N__57635\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57627\ : std_logic;
signal \N__57626\ : std_logic;
signal \N__57625\ : std_logic;
signal \N__57624\ : std_logic;
signal \N__57619\ : std_logic;
signal \N__57618\ : std_logic;
signal \N__57617\ : std_logic;
signal \N__57616\ : std_logic;
signal \N__57615\ : std_logic;
signal \N__57614\ : std_logic;
signal \N__57611\ : std_logic;
signal \N__57608\ : std_logic;
signal \N__57605\ : std_logic;
signal \N__57604\ : std_logic;
signal \N__57603\ : std_logic;
signal \N__57600\ : std_logic;
signal \N__57597\ : std_logic;
signal \N__57594\ : std_logic;
signal \N__57593\ : std_logic;
signal \N__57592\ : std_logic;
signal \N__57591\ : std_logic;
signal \N__57590\ : std_logic;
signal \N__57589\ : std_logic;
signal \N__57588\ : std_logic;
signal \N__57585\ : std_logic;
signal \N__57582\ : std_logic;
signal \N__57579\ : std_logic;
signal \N__57576\ : std_logic;
signal \N__57573\ : std_logic;
signal \N__57572\ : std_logic;
signal \N__57569\ : std_logic;
signal \N__57564\ : std_logic;
signal \N__57561\ : std_logic;
signal \N__57558\ : std_logic;
signal \N__57555\ : std_logic;
signal \N__57554\ : std_logic;
signal \N__57553\ : std_logic;
signal \N__57550\ : std_logic;
signal \N__57547\ : std_logic;
signal \N__57544\ : std_logic;
signal \N__57539\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57527\ : std_logic;
signal \N__57524\ : std_logic;
signal \N__57521\ : std_logic;
signal \N__57508\ : std_logic;
signal \N__57505\ : std_logic;
signal \N__57500\ : std_logic;
signal \N__57499\ : std_logic;
signal \N__57498\ : std_logic;
signal \N__57493\ : std_logic;
signal \N__57490\ : std_logic;
signal \N__57487\ : std_logic;
signal \N__57484\ : std_logic;
signal \N__57481\ : std_logic;
signal \N__57478\ : std_logic;
signal \N__57477\ : std_logic;
signal \N__57476\ : std_logic;
signal \N__57475\ : std_logic;
signal \N__57474\ : std_logic;
signal \N__57467\ : std_logic;
signal \N__57462\ : std_logic;
signal \N__57459\ : std_logic;
signal \N__57456\ : std_logic;
signal \N__57451\ : std_logic;
signal \N__57446\ : std_logic;
signal \N__57443\ : std_logic;
signal \N__57440\ : std_logic;
signal \N__57437\ : std_logic;
signal \N__57434\ : std_logic;
signal \N__57423\ : std_logic;
signal \N__57416\ : std_logic;
signal \N__57411\ : std_logic;
signal \N__57404\ : std_logic;
signal \N__57399\ : std_logic;
signal \N__57394\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57388\ : std_logic;
signal \N__57387\ : std_logic;
signal \N__57386\ : std_logic;
signal \N__57385\ : std_logic;
signal \N__57384\ : std_logic;
signal \N__57383\ : std_logic;
signal \N__57382\ : std_logic;
signal \N__57381\ : std_logic;
signal \N__57370\ : std_logic;
signal \N__57367\ : std_logic;
signal \N__57362\ : std_logic;
signal \N__57355\ : std_logic;
signal \N__57352\ : std_logic;
signal \N__57349\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57335\ : std_logic;
signal \N__57330\ : std_logic;
signal \N__57323\ : std_logic;
signal \N__57320\ : std_logic;
signal \N__57317\ : std_logic;
signal \N__57312\ : std_logic;
signal \N__57303\ : std_logic;
signal \N__57300\ : std_logic;
signal \N__57293\ : std_logic;
signal \N__57288\ : std_logic;
signal \N__57281\ : std_logic;
signal \N__57278\ : std_logic;
signal \N__57263\ : std_logic;
signal \N__57262\ : std_logic;
signal \N__57261\ : std_logic;
signal \N__57258\ : std_logic;
signal \N__57251\ : std_logic;
signal \N__57246\ : std_logic;
signal \N__57241\ : std_logic;
signal \N__57232\ : std_logic;
signal \N__57225\ : std_logic;
signal \N__57222\ : std_logic;
signal \N__57215\ : std_logic;
signal \N__57208\ : std_logic;
signal \N__57199\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57181\ : std_logic;
signal \N__57156\ : std_logic;
signal \N__57153\ : std_logic;
signal \N__57150\ : std_logic;
signal \N__57147\ : std_logic;
signal \N__57144\ : std_logic;
signal \N__57143\ : std_logic;
signal \N__57140\ : std_logic;
signal \N__57139\ : std_logic;
signal \N__57138\ : std_logic;
signal \N__57135\ : std_logic;
signal \N__57134\ : std_logic;
signal \N__57133\ : std_logic;
signal \N__57132\ : std_logic;
signal \N__57127\ : std_logic;
signal \N__57126\ : std_logic;
signal \N__57125\ : std_logic;
signal \N__57124\ : std_logic;
signal \N__57123\ : std_logic;
signal \N__57122\ : std_logic;
signal \N__57119\ : std_logic;
signal \N__57118\ : std_logic;
signal \N__57115\ : std_logic;
signal \N__57110\ : std_logic;
signal \N__57109\ : std_logic;
signal \N__57108\ : std_logic;
signal \N__57105\ : std_logic;
signal \N__57102\ : std_logic;
signal \N__57099\ : std_logic;
signal \N__57098\ : std_logic;
signal \N__57097\ : std_logic;
signal \N__57096\ : std_logic;
signal \N__57095\ : std_logic;
signal \N__57094\ : std_logic;
signal \N__57093\ : std_logic;
signal \N__57092\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57090\ : std_logic;
signal \N__57089\ : std_logic;
signal \N__57088\ : std_logic;
signal \N__57087\ : std_logic;
signal \N__57082\ : std_logic;
signal \N__57079\ : std_logic;
signal \N__57076\ : std_logic;
signal \N__57073\ : std_logic;
signal \N__57070\ : std_logic;
signal \N__57069\ : std_logic;
signal \N__57068\ : std_logic;
signal \N__57067\ : std_logic;
signal \N__57066\ : std_logic;
signal \N__57065\ : std_logic;
signal \N__57064\ : std_logic;
signal \N__57063\ : std_logic;
signal \N__57062\ : std_logic;
signal \N__57061\ : std_logic;
signal \N__57060\ : std_logic;
signal \N__57059\ : std_logic;
signal \N__57056\ : std_logic;
signal \N__57053\ : std_logic;
signal \N__57050\ : std_logic;
signal \N__57049\ : std_logic;
signal \N__57046\ : std_logic;
signal \N__57043\ : std_logic;
signal \N__57038\ : std_logic;
signal \N__57035\ : std_logic;
signal \N__57032\ : std_logic;
signal \N__57029\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57025\ : std_logic;
signal \N__57024\ : std_logic;
signal \N__57023\ : std_logic;
signal \N__57022\ : std_logic;
signal \N__57021\ : std_logic;
signal \N__57016\ : std_logic;
signal \N__57015\ : std_logic;
signal \N__57014\ : std_logic;
signal \N__57013\ : std_logic;
signal \N__57008\ : std_logic;
signal \N__57005\ : std_logic;
signal \N__57004\ : std_logic;
signal \N__57001\ : std_logic;
signal \N__57000\ : std_logic;
signal \N__56999\ : std_logic;
signal \N__56996\ : std_logic;
signal \N__56993\ : std_logic;
signal \N__56992\ : std_logic;
signal \N__56983\ : std_logic;
signal \N__56980\ : std_logic;
signal \N__56973\ : std_logic;
signal \N__56968\ : std_logic;
signal \N__56959\ : std_logic;
signal \N__56958\ : std_logic;
signal \N__56957\ : std_logic;
signal \N__56956\ : std_logic;
signal \N__56955\ : std_logic;
signal \N__56954\ : std_logic;
signal \N__56953\ : std_logic;
signal \N__56948\ : std_logic;
signal \N__56947\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56945\ : std_logic;
signal \N__56940\ : std_logic;
signal \N__56937\ : std_logic;
signal \N__56936\ : std_logic;
signal \N__56935\ : std_logic;
signal \N__56934\ : std_logic;
signal \N__56933\ : std_logic;
signal \N__56932\ : std_logic;
signal \N__56931\ : std_logic;
signal \N__56930\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56928\ : std_logic;
signal \N__56927\ : std_logic;
signal \N__56926\ : std_logic;
signal \N__56925\ : std_logic;
signal \N__56924\ : std_logic;
signal \N__56923\ : std_logic;
signal \N__56920\ : std_logic;
signal \N__56917\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56902\ : std_logic;
signal \N__56901\ : std_logic;
signal \N__56900\ : std_logic;
signal \N__56899\ : std_logic;
signal \N__56888\ : std_logic;
signal \N__56885\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56872\ : std_logic;
signal \N__56869\ : std_logic;
signal \N__56868\ : std_logic;
signal \N__56867\ : std_logic;
signal \N__56866\ : std_logic;
signal \N__56865\ : std_logic;
signal \N__56864\ : std_logic;
signal \N__56863\ : std_logic;
signal \N__56860\ : std_logic;
signal \N__56857\ : std_logic;
signal \N__56854\ : std_logic;
signal \N__56853\ : std_logic;
signal \N__56852\ : std_logic;
signal \N__56845\ : std_logic;
signal \N__56842\ : std_logic;
signal \N__56835\ : std_logic;
signal \N__56832\ : std_logic;
signal \N__56831\ : std_logic;
signal \N__56830\ : std_logic;
signal \N__56827\ : std_logic;
signal \N__56826\ : std_logic;
signal \N__56825\ : std_logic;
signal \N__56824\ : std_logic;
signal \N__56823\ : std_logic;
signal \N__56822\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56808\ : std_logic;
signal \N__56801\ : std_logic;
signal \N__56796\ : std_logic;
signal \N__56787\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56773\ : std_logic;
signal \N__56768\ : std_logic;
signal \N__56763\ : std_logic;
signal \N__56760\ : std_logic;
signal \N__56757\ : std_logic;
signal \N__56752\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56732\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56724\ : std_logic;
signal \N__56715\ : std_logic;
signal \N__56708\ : std_logic;
signal \N__56703\ : std_logic;
signal \N__56694\ : std_logic;
signal \N__56693\ : std_logic;
signal \N__56692\ : std_logic;
signal \N__56689\ : std_logic;
signal \N__56686\ : std_logic;
signal \N__56683\ : std_logic;
signal \N__56676\ : std_logic;
signal \N__56671\ : std_logic;
signal \N__56668\ : std_logic;
signal \N__56651\ : std_logic;
signal \N__56640\ : std_logic;
signal \N__56629\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56621\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56595\ : std_logic;
signal \N__56594\ : std_logic;
signal \N__56591\ : std_logic;
signal \N__56588\ : std_logic;
signal \N__56585\ : std_logic;
signal \N__56582\ : std_logic;
signal \N__56579\ : std_logic;
signal \N__56576\ : std_logic;
signal \N__56571\ : std_logic;
signal \N__56568\ : std_logic;
signal \N__56567\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56563\ : std_logic;
signal \N__56562\ : std_logic;
signal \N__56561\ : std_logic;
signal \N__56560\ : std_logic;
signal \N__56559\ : std_logic;
signal \N__56558\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56556\ : std_logic;
signal \N__56555\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56553\ : std_logic;
signal \N__56552\ : std_logic;
signal \N__56551\ : std_logic;
signal \N__56550\ : std_logic;
signal \N__56549\ : std_logic;
signal \N__56548\ : std_logic;
signal \N__56547\ : std_logic;
signal \N__56546\ : std_logic;
signal \N__56545\ : std_logic;
signal \N__56544\ : std_logic;
signal \N__56541\ : std_logic;
signal \N__56540\ : std_logic;
signal \N__56539\ : std_logic;
signal \N__56532\ : std_logic;
signal \N__56527\ : std_logic;
signal \N__56520\ : std_logic;
signal \N__56519\ : std_logic;
signal \N__56518\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56516\ : std_logic;
signal \N__56513\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56506\ : std_logic;
signal \N__56505\ : std_logic;
signal \N__56504\ : std_logic;
signal \N__56501\ : std_logic;
signal \N__56500\ : std_logic;
signal \N__56499\ : std_logic;
signal \N__56498\ : std_logic;
signal \N__56497\ : std_logic;
signal \N__56494\ : std_logic;
signal \N__56489\ : std_logic;
signal \N__56488\ : std_logic;
signal \N__56485\ : std_logic;
signal \N__56484\ : std_logic;
signal \N__56483\ : std_logic;
signal \N__56482\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56480\ : std_logic;
signal \N__56479\ : std_logic;
signal \N__56478\ : std_logic;
signal \N__56477\ : std_logic;
signal \N__56476\ : std_logic;
signal \N__56475\ : std_logic;
signal \N__56474\ : std_logic;
signal \N__56473\ : std_logic;
signal \N__56472\ : std_logic;
signal \N__56471\ : std_logic;
signal \N__56468\ : std_logic;
signal \N__56467\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56459\ : std_logic;
signal \N__56456\ : std_logic;
signal \N__56453\ : std_logic;
signal \N__56452\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56450\ : std_logic;
signal \N__56447\ : std_logic;
signal \N__56446\ : std_logic;
signal \N__56445\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56433\ : std_logic;
signal \N__56430\ : std_logic;
signal \N__56427\ : std_logic;
signal \N__56424\ : std_logic;
signal \N__56421\ : std_logic;
signal \N__56420\ : std_logic;
signal \N__56419\ : std_logic;
signal \N__56414\ : std_logic;
signal \N__56409\ : std_logic;
signal \N__56406\ : std_logic;
signal \N__56401\ : std_logic;
signal \N__56400\ : std_logic;
signal \N__56395\ : std_logic;
signal \N__56390\ : std_logic;
signal \N__56387\ : std_logic;
signal \N__56384\ : std_logic;
signal \N__56379\ : std_logic;
signal \N__56364\ : std_logic;
signal \N__56361\ : std_logic;
signal \N__56358\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56356\ : std_logic;
signal \N__56351\ : std_logic;
signal \N__56348\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56344\ : std_logic;
signal \N__56343\ : std_logic;
signal \N__56334\ : std_logic;
signal \N__56331\ : std_logic;
signal \N__56328\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56321\ : std_logic;
signal \N__56320\ : std_logic;
signal \N__56317\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56315\ : std_logic;
signal \N__56312\ : std_logic;
signal \N__56305\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56293\ : std_logic;
signal \N__56292\ : std_logic;
signal \N__56291\ : std_logic;
signal \N__56288\ : std_logic;
signal \N__56281\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56275\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56267\ : std_logic;
signal \N__56264\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56240\ : std_logic;
signal \N__56237\ : std_logic;
signal \N__56232\ : std_logic;
signal \N__56229\ : std_logic;
signal \N__56228\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56223\ : std_logic;
signal \N__56222\ : std_logic;
signal \N__56221\ : std_logic;
signal \N__56220\ : std_logic;
signal \N__56215\ : std_logic;
signal \N__56212\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56203\ : std_logic;
signal \N__56202\ : std_logic;
signal \N__56199\ : std_logic;
signal \N__56196\ : std_logic;
signal \N__56191\ : std_logic;
signal \N__56188\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56180\ : std_logic;
signal \N__56179\ : std_logic;
signal \N__56176\ : std_logic;
signal \N__56175\ : std_logic;
signal \N__56174\ : std_logic;
signal \N__56171\ : std_logic;
signal \N__56170\ : std_logic;
signal \N__56169\ : std_logic;
signal \N__56168\ : std_logic;
signal \N__56165\ : std_logic;
signal \N__56160\ : std_logic;
signal \N__56157\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56143\ : std_logic;
signal \N__56136\ : std_logic;
signal \N__56129\ : std_logic;
signal \N__56124\ : std_logic;
signal \N__56121\ : std_logic;
signal \N__56116\ : std_logic;
signal \N__56109\ : std_logic;
signal \N__56100\ : std_logic;
signal \N__56091\ : std_logic;
signal \N__56084\ : std_logic;
signal \N__56075\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56054\ : std_logic;
signal \N__56031\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56027\ : std_logic;
signal \N__56024\ : std_logic;
signal \N__56021\ : std_logic;
signal \N__56018\ : std_logic;
signal \N__56015\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56004\ : std_logic;
signal \N__56001\ : std_logic;
signal \N__55998\ : std_logic;
signal \N__55995\ : std_logic;
signal \N__55992\ : std_logic;
signal \N__55989\ : std_logic;
signal \N__55986\ : std_logic;
signal \N__55983\ : std_logic;
signal \N__55980\ : std_logic;
signal \N__55977\ : std_logic;
signal \N__55974\ : std_logic;
signal \N__55971\ : std_logic;
signal \N__55968\ : std_logic;
signal \N__55967\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55958\ : std_logic;
signal \N__55955\ : std_logic;
signal \N__55952\ : std_logic;
signal \N__55949\ : std_logic;
signal \N__55946\ : std_logic;
signal \N__55943\ : std_logic;
signal \N__55940\ : std_logic;
signal \N__55937\ : std_logic;
signal \N__55934\ : std_logic;
signal \N__55931\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55925\ : std_logic;
signal \N__55922\ : std_logic;
signal \N__55917\ : std_logic;
signal \N__55914\ : std_logic;
signal \N__55911\ : std_logic;
signal \N__55908\ : std_logic;
signal \N__55905\ : std_logic;
signal \N__55902\ : std_logic;
signal \N__55901\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55897\ : std_logic;
signal \N__55894\ : std_logic;
signal \N__55891\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55874\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55871\ : std_logic;
signal \N__55870\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55868\ : std_logic;
signal \N__55867\ : std_logic;
signal \N__55866\ : std_logic;
signal \N__55865\ : std_logic;
signal \N__55862\ : std_logic;
signal \N__55859\ : std_logic;
signal \N__55858\ : std_logic;
signal \N__55857\ : std_logic;
signal \N__55854\ : std_logic;
signal \N__55851\ : std_logic;
signal \N__55850\ : std_logic;
signal \N__55849\ : std_logic;
signal \N__55848\ : std_logic;
signal \N__55847\ : std_logic;
signal \N__55844\ : std_logic;
signal \N__55843\ : std_logic;
signal \N__55840\ : std_logic;
signal \N__55837\ : std_logic;
signal \N__55834\ : std_logic;
signal \N__55833\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55831\ : std_logic;
signal \N__55828\ : std_logic;
signal \N__55827\ : std_logic;
signal \N__55824\ : std_logic;
signal \N__55821\ : std_logic;
signal \N__55820\ : std_logic;
signal \N__55819\ : std_logic;
signal \N__55818\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55816\ : std_logic;
signal \N__55811\ : std_logic;
signal \N__55810\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55792\ : std_logic;
signal \N__55787\ : std_logic;
signal \N__55782\ : std_logic;
signal \N__55779\ : std_logic;
signal \N__55778\ : std_logic;
signal \N__55777\ : std_logic;
signal \N__55772\ : std_logic;
signal \N__55769\ : std_logic;
signal \N__55766\ : std_logic;
signal \N__55765\ : std_logic;
signal \N__55764\ : std_logic;
signal \N__55763\ : std_logic;
signal \N__55760\ : std_logic;
signal \N__55759\ : std_logic;
signal \N__55758\ : std_logic;
signal \N__55757\ : std_logic;
signal \N__55752\ : std_logic;
signal \N__55749\ : std_logic;
signal \N__55742\ : std_logic;
signal \N__55739\ : std_logic;
signal \N__55736\ : std_logic;
signal \N__55733\ : std_logic;
signal \N__55730\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55720\ : std_logic;
signal \N__55717\ : std_logic;
signal \N__55714\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55699\ : std_logic;
signal \N__55696\ : std_logic;
signal \N__55689\ : std_logic;
signal \N__55680\ : std_logic;
signal \N__55677\ : std_logic;
signal \N__55674\ : std_logic;
signal \N__55667\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55649\ : std_logic;
signal \N__55638\ : std_logic;
signal \N__55637\ : std_logic;
signal \N__55636\ : std_logic;
signal \N__55633\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55627\ : std_logic;
signal \N__55624\ : std_logic;
signal \N__55621\ : std_logic;
signal \N__55618\ : std_logic;
signal \N__55615\ : std_logic;
signal \N__55614\ : std_logic;
signal \N__55611\ : std_logic;
signal \N__55608\ : std_logic;
signal \N__55605\ : std_logic;
signal \N__55602\ : std_logic;
signal \N__55601\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55595\ : std_logic;
signal \N__55590\ : std_logic;
signal \N__55587\ : std_logic;
signal \N__55578\ : std_logic;
signal \N__55575\ : std_logic;
signal \N__55572\ : std_logic;
signal \N__55569\ : std_logic;
signal \N__55566\ : std_logic;
signal \N__55563\ : std_logic;
signal \N__55560\ : std_logic;
signal \N__55557\ : std_logic;
signal \N__55556\ : std_logic;
signal \N__55553\ : std_logic;
signal \N__55552\ : std_logic;
signal \N__55551\ : std_logic;
signal \N__55550\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55547\ : std_logic;
signal \N__55546\ : std_logic;
signal \N__55545\ : std_logic;
signal \N__55544\ : std_logic;
signal \N__55543\ : std_logic;
signal \N__55542\ : std_logic;
signal \N__55541\ : std_logic;
signal \N__55538\ : std_logic;
signal \N__55535\ : std_logic;
signal \N__55526\ : std_logic;
signal \N__55525\ : std_logic;
signal \N__55524\ : std_logic;
signal \N__55523\ : std_logic;
signal \N__55522\ : std_logic;
signal \N__55519\ : std_logic;
signal \N__55518\ : std_logic;
signal \N__55517\ : std_logic;
signal \N__55516\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55514\ : std_logic;
signal \N__55513\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55511\ : std_logic;
signal \N__55510\ : std_logic;
signal \N__55507\ : std_logic;
signal \N__55504\ : std_logic;
signal \N__55501\ : std_logic;
signal \N__55500\ : std_logic;
signal \N__55499\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55486\ : std_logic;
signal \N__55481\ : std_logic;
signal \N__55480\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55467\ : std_logic;
signal \N__55464\ : std_logic;
signal \N__55459\ : std_logic;
signal \N__55452\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55434\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55429\ : std_logic;
signal \N__55426\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55422\ : std_logic;
signal \N__55421\ : std_logic;
signal \N__55418\ : std_logic;
signal \N__55415\ : std_logic;
signal \N__55412\ : std_logic;
signal \N__55409\ : std_logic;
signal \N__55408\ : std_logic;
signal \N__55407\ : std_logic;
signal \N__55406\ : std_logic;
signal \N__55405\ : std_logic;
signal \N__55404\ : std_logic;
signal \N__55397\ : std_logic;
signal \N__55394\ : std_logic;
signal \N__55391\ : std_logic;
signal \N__55388\ : std_logic;
signal \N__55385\ : std_logic;
signal \N__55380\ : std_logic;
signal \N__55375\ : std_logic;
signal \N__55370\ : std_logic;
signal \N__55365\ : std_logic;
signal \N__55360\ : std_logic;
signal \N__55357\ : std_logic;
signal \N__55354\ : std_logic;
signal \N__55353\ : std_logic;
signal \N__55352\ : std_logic;
signal \N__55351\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55349\ : std_logic;
signal \N__55348\ : std_logic;
signal \N__55339\ : std_logic;
signal \N__55336\ : std_logic;
signal \N__55331\ : std_logic;
signal \N__55326\ : std_logic;
signal \N__55317\ : std_logic;
signal \N__55314\ : std_logic;
signal \N__55309\ : std_logic;
signal \N__55302\ : std_logic;
signal \N__55299\ : std_logic;
signal \N__55296\ : std_logic;
signal \N__55287\ : std_logic;
signal \N__55282\ : std_logic;
signal \N__55277\ : std_logic;
signal \N__55270\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55248\ : std_logic;
signal \N__55245\ : std_logic;
signal \N__55242\ : std_logic;
signal \N__55239\ : std_logic;
signal \N__55236\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55233\ : std_logic;
signal \N__55232\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55225\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55219\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55216\ : std_logic;
signal \N__55215\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55213\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55211\ : std_logic;
signal \N__55210\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55208\ : std_logic;
signal \N__55205\ : std_logic;
signal \N__55200\ : std_logic;
signal \N__55195\ : std_logic;
signal \N__55190\ : std_logic;
signal \N__55189\ : std_logic;
signal \N__55188\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55184\ : std_logic;
signal \N__55177\ : std_logic;
signal \N__55176\ : std_logic;
signal \N__55175\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55173\ : std_logic;
signal \N__55172\ : std_logic;
signal \N__55171\ : std_logic;
signal \N__55170\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55161\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55159\ : std_logic;
signal \N__55158\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55155\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55153\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55150\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55148\ : std_logic;
signal \N__55147\ : std_logic;
signal \N__55146\ : std_logic;
signal \N__55145\ : std_logic;
signal \N__55142\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55140\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55136\ : std_logic;
signal \N__55133\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55116\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55104\ : std_logic;
signal \N__55101\ : std_logic;
signal \N__55098\ : std_logic;
signal \N__55095\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55071\ : std_logic;
signal \N__55066\ : std_logic;
signal \N__55063\ : std_logic;
signal \N__55060\ : std_logic;
signal \N__55059\ : std_logic;
signal \N__55058\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55056\ : std_logic;
signal \N__55053\ : std_logic;
signal \N__55050\ : std_logic;
signal \N__55047\ : std_logic;
signal \N__55042\ : std_logic;
signal \N__55037\ : std_logic;
signal \N__55036\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55034\ : std_logic;
signal \N__55029\ : std_logic;
signal \N__55026\ : std_logic;
signal \N__55023\ : std_logic;
signal \N__55022\ : std_logic;
signal \N__55019\ : std_logic;
signal \N__55012\ : std_logic;
signal \N__55009\ : std_logic;
signal \N__55006\ : std_logic;
signal \N__55003\ : std_logic;
signal \N__54996\ : std_logic;
signal \N__54993\ : std_logic;
signal \N__54990\ : std_logic;
signal \N__54985\ : std_logic;
signal \N__54980\ : std_logic;
signal \N__54979\ : std_logic;
signal \N__54978\ : std_logic;
signal \N__54975\ : std_logic;
signal \N__54968\ : std_logic;
signal \N__54965\ : std_logic;
signal \N__54962\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54956\ : std_logic;
signal \N__54953\ : std_logic;
signal \N__54950\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54944\ : std_logic;
signal \N__54941\ : std_logic;
signal \N__54930\ : std_logic;
signal \N__54925\ : std_logic;
signal \N__54922\ : std_logic;
signal \N__54917\ : std_logic;
signal \N__54914\ : std_logic;
signal \N__54913\ : std_logic;
signal \N__54910\ : std_logic;
signal \N__54907\ : std_logic;
signal \N__54904\ : std_logic;
signal \N__54895\ : std_logic;
signal \N__54892\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54874\ : std_logic;
signal \N__54869\ : std_logic;
signal \N__54868\ : std_logic;
signal \N__54865\ : std_logic;
signal \N__54860\ : std_logic;
signal \N__54857\ : std_logic;
signal \N__54852\ : std_logic;
signal \N__54849\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54837\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54832\ : std_logic;
signal \N__54827\ : std_logic;
signal \N__54818\ : std_logic;
signal \N__54815\ : std_logic;
signal \N__54808\ : std_logic;
signal \N__54805\ : std_logic;
signal \N__54800\ : std_logic;
signal \N__54791\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54765\ : std_logic;
signal \N__54764\ : std_logic;
signal \N__54763\ : std_logic;
signal \N__54762\ : std_logic;
signal \N__54761\ : std_logic;
signal \N__54760\ : std_logic;
signal \N__54759\ : std_logic;
signal \N__54758\ : std_logic;
signal \N__54757\ : std_logic;
signal \N__54756\ : std_logic;
signal \N__54755\ : std_logic;
signal \N__54754\ : std_logic;
signal \N__54753\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54749\ : std_logic;
signal \N__54748\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54746\ : std_logic;
signal \N__54745\ : std_logic;
signal \N__54744\ : std_logic;
signal \N__54741\ : std_logic;
signal \N__54738\ : std_logic;
signal \N__54733\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54723\ : std_logic;
signal \N__54720\ : std_logic;
signal \N__54719\ : std_logic;
signal \N__54716\ : std_logic;
signal \N__54713\ : std_logic;
signal \N__54712\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54708\ : std_logic;
signal \N__54707\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54698\ : std_logic;
signal \N__54697\ : std_logic;
signal \N__54696\ : std_logic;
signal \N__54695\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54693\ : std_logic;
signal \N__54692\ : std_logic;
signal \N__54691\ : std_logic;
signal \N__54688\ : std_logic;
signal \N__54687\ : std_logic;
signal \N__54686\ : std_logic;
signal \N__54683\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54677\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54665\ : std_logic;
signal \N__54662\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54654\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54648\ : std_logic;
signal \N__54645\ : std_logic;
signal \N__54644\ : std_logic;
signal \N__54641\ : std_logic;
signal \N__54638\ : std_logic;
signal \N__54635\ : std_logic;
signal \N__54632\ : std_logic;
signal \N__54631\ : std_logic;
signal \N__54628\ : std_logic;
signal \N__54625\ : std_logic;
signal \N__54622\ : std_logic;
signal \N__54619\ : std_logic;
signal \N__54614\ : std_logic;
signal \N__54611\ : std_logic;
signal \N__54608\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54602\ : std_logic;
signal \N__54601\ : std_logic;
signal \N__54598\ : std_logic;
signal \N__54595\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54579\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54570\ : std_logic;
signal \N__54569\ : std_logic;
signal \N__54566\ : std_logic;
signal \N__54563\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54555\ : std_logic;
signal \N__54554\ : std_logic;
signal \N__54551\ : std_logic;
signal \N__54546\ : std_logic;
signal \N__54539\ : std_logic;
signal \N__54532\ : std_logic;
signal \N__54529\ : std_logic;
signal \N__54526\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54505\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54493\ : std_logic;
signal \N__54490\ : std_logic;
signal \N__54481\ : std_logic;
signal \N__54478\ : std_logic;
signal \N__54459\ : std_logic;
signal \N__54456\ : std_logic;
signal \N__54453\ : std_logic;
signal \N__54450\ : std_logic;
signal \N__54449\ : std_logic;
signal \N__54446\ : std_logic;
signal \N__54443\ : std_logic;
signal \N__54438\ : std_logic;
signal \N__54437\ : std_logic;
signal \N__54436\ : std_logic;
signal \N__54435\ : std_logic;
signal \N__54434\ : std_logic;
signal \N__54433\ : std_logic;
signal \N__54432\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54430\ : std_logic;
signal \N__54429\ : std_logic;
signal \N__54428\ : std_logic;
signal \N__54427\ : std_logic;
signal \N__54426\ : std_logic;
signal \N__54425\ : std_logic;
signal \N__54424\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54421\ : std_logic;
signal \N__54420\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54418\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54415\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54413\ : std_logic;
signal \N__54412\ : std_logic;
signal \N__54411\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54409\ : std_logic;
signal \N__54408\ : std_logic;
signal \N__54407\ : std_logic;
signal \N__54406\ : std_logic;
signal \N__54405\ : std_logic;
signal \N__54404\ : std_logic;
signal \N__54403\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54400\ : std_logic;
signal \N__54399\ : std_logic;
signal \N__54398\ : std_logic;
signal \N__54397\ : std_logic;
signal \N__54396\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54394\ : std_logic;
signal \N__54393\ : std_logic;
signal \N__54392\ : std_logic;
signal \N__54391\ : std_logic;
signal \N__54390\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54388\ : std_logic;
signal \N__54387\ : std_logic;
signal \N__54386\ : std_logic;
signal \N__54385\ : std_logic;
signal \N__54384\ : std_logic;
signal \N__54383\ : std_logic;
signal \N__54382\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54380\ : std_logic;
signal \N__54379\ : std_logic;
signal \N__54378\ : std_logic;
signal \N__54377\ : std_logic;
signal \N__54376\ : std_logic;
signal \N__54375\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54372\ : std_logic;
signal \N__54371\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54369\ : std_logic;
signal \N__54368\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54366\ : std_logic;
signal \N__54365\ : std_logic;
signal \N__54364\ : std_logic;
signal \N__54363\ : std_logic;
signal \N__54362\ : std_logic;
signal \N__54361\ : std_logic;
signal \N__54360\ : std_logic;
signal \N__54359\ : std_logic;
signal \N__54358\ : std_logic;
signal \N__54357\ : std_logic;
signal \N__54356\ : std_logic;
signal \N__54355\ : std_logic;
signal \N__54354\ : std_logic;
signal \N__54353\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54350\ : std_logic;
signal \N__54349\ : std_logic;
signal \N__54348\ : std_logic;
signal \N__54347\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54345\ : std_logic;
signal \N__54344\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54342\ : std_logic;
signal \N__54341\ : std_logic;
signal \N__54340\ : std_logic;
signal \N__54339\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54335\ : std_logic;
signal \N__54334\ : std_logic;
signal \N__54333\ : std_logic;
signal \N__54332\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54330\ : std_logic;
signal \N__54329\ : std_logic;
signal \N__54328\ : std_logic;
signal \N__54327\ : std_logic;
signal \N__54326\ : std_logic;
signal \N__54325\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54322\ : std_logic;
signal \N__54321\ : std_logic;
signal \N__54320\ : std_logic;
signal \N__54319\ : std_logic;
signal \N__54318\ : std_logic;
signal \N__54317\ : std_logic;
signal \N__54316\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54314\ : std_logic;
signal \N__54313\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54311\ : std_logic;
signal \N__54310\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54307\ : std_logic;
signal \N__54306\ : std_logic;
signal \N__54305\ : std_logic;
signal \N__54304\ : std_logic;
signal \N__54303\ : std_logic;
signal \N__54302\ : std_logic;
signal \N__54301\ : std_logic;
signal \N__54300\ : std_logic;
signal \N__54299\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54296\ : std_logic;
signal \N__54295\ : std_logic;
signal \N__54294\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54292\ : std_logic;
signal \N__54291\ : std_logic;
signal \N__54290\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54287\ : std_logic;
signal \N__54286\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54284\ : std_logic;
signal \N__54283\ : std_logic;
signal \N__54282\ : std_logic;
signal \N__54281\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54279\ : std_logic;
signal \N__54278\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54276\ : std_logic;
signal \N__54275\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54273\ : std_logic;
signal \N__54272\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54270\ : std_logic;
signal \N__54269\ : std_logic;
signal \N__53928\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53924\ : std_logic;
signal \N__53921\ : std_logic;
signal \N__53918\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53914\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53901\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53892\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53886\ : std_logic;
signal \N__53883\ : std_logic;
signal \N__53880\ : std_logic;
signal \N__53877\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53868\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53850\ : std_logic;
signal \N__53847\ : std_logic;
signal \N__53844\ : std_logic;
signal \N__53841\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53831\ : std_logic;
signal \N__53828\ : std_logic;
signal \N__53825\ : std_logic;
signal \N__53822\ : std_logic;
signal \N__53819\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53810\ : std_logic;
signal \N__53807\ : std_logic;
signal \N__53804\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53798\ : std_logic;
signal \N__53797\ : std_logic;
signal \N__53796\ : std_logic;
signal \N__53795\ : std_logic;
signal \N__53794\ : std_logic;
signal \N__53793\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53790\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53787\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53784\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53781\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53778\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53772\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53768\ : std_logic;
signal \N__53767\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53764\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53762\ : std_logic;
signal \N__53761\ : std_logic;
signal \N__53758\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53755\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53751\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53749\ : std_logic;
signal \N__53746\ : std_logic;
signal \N__53739\ : std_logic;
signal \N__53730\ : std_logic;
signal \N__53729\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53724\ : std_logic;
signal \N__53723\ : std_logic;
signal \N__53722\ : std_logic;
signal \N__53721\ : std_logic;
signal \N__53720\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53707\ : std_logic;
signal \N__53704\ : std_logic;
signal \N__53699\ : std_logic;
signal \N__53696\ : std_logic;
signal \N__53693\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53687\ : std_logic;
signal \N__53684\ : std_logic;
signal \N__53683\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53681\ : std_logic;
signal \N__53680\ : std_logic;
signal \N__53679\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53673\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53671\ : std_logic;
signal \N__53670\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53668\ : std_logic;
signal \N__53667\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53659\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53642\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53634\ : std_logic;
signal \N__53631\ : std_logic;
signal \N__53628\ : std_logic;
signal \N__53621\ : std_logic;
signal \N__53618\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53614\ : std_logic;
signal \N__53613\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53611\ : std_logic;
signal \N__53608\ : std_logic;
signal \N__53605\ : std_logic;
signal \N__53602\ : std_logic;
signal \N__53597\ : std_logic;
signal \N__53590\ : std_logic;
signal \N__53585\ : std_logic;
signal \N__53580\ : std_logic;
signal \N__53577\ : std_logic;
signal \N__53568\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53559\ : std_logic;
signal \N__53556\ : std_logic;
signal \N__53555\ : std_logic;
signal \N__53554\ : std_logic;
signal \N__53553\ : std_logic;
signal \N__53552\ : std_logic;
signal \N__53549\ : std_logic;
signal \N__53548\ : std_logic;
signal \N__53545\ : std_logic;
signal \N__53536\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53513\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53507\ : std_logic;
signal \N__53502\ : std_logic;
signal \N__53499\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53489\ : std_logic;
signal \N__53486\ : std_logic;
signal \N__53483\ : std_logic;
signal \N__53480\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53472\ : std_logic;
signal \N__53469\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53459\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53454\ : std_logic;
signal \N__53447\ : std_logic;
signal \N__53444\ : std_logic;
signal \N__53441\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53423\ : std_logic;
signal \N__53420\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53397\ : std_logic;
signal \N__53388\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53355\ : std_logic;
signal \N__53352\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53348\ : std_logic;
signal \N__53345\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53334\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53328\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53324\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53315\ : std_logic;
signal \N__53312\ : std_logic;
signal \N__53309\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53301\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53299\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53294\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53288\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53279\ : std_logic;
signal \N__53278\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53276\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53269\ : std_logic;
signal \N__53266\ : std_logic;
signal \N__53265\ : std_logic;
signal \N__53262\ : std_logic;
signal \N__53261\ : std_logic;
signal \N__53260\ : std_logic;
signal \N__53257\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53254\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53234\ : std_logic;
signal \N__53231\ : std_logic;
signal \N__53228\ : std_logic;
signal \N__53225\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53214\ : std_logic;
signal \N__53211\ : std_logic;
signal \N__53208\ : std_logic;
signal \N__53207\ : std_logic;
signal \N__53204\ : std_logic;
signal \N__53201\ : std_logic;
signal \N__53198\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53191\ : std_logic;
signal \N__53188\ : std_logic;
signal \N__53183\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53173\ : std_logic;
signal \N__53168\ : std_logic;
signal \N__53163\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53155\ : std_logic;
signal \N__53152\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53139\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53106\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53100\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53076\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53047\ : std_logic;
signal \N__53044\ : std_logic;
signal \N__53041\ : std_logic;
signal \N__53040\ : std_logic;
signal \N__53039\ : std_logic;
signal \N__53038\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53036\ : std_logic;
signal \N__53035\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53027\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52995\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52980\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52950\ : std_logic;
signal \N__52949\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52945\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52923\ : std_logic;
signal \N__52920\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52914\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52907\ : std_logic;
signal \N__52906\ : std_logic;
signal \N__52901\ : std_logic;
signal \N__52898\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52893\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52887\ : std_logic;
signal \N__52882\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52859\ : std_logic;
signal \N__52856\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52841\ : std_logic;
signal \N__52840\ : std_logic;
signal \N__52837\ : std_logic;
signal \N__52834\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52821\ : std_logic;
signal \N__52818\ : std_logic;
signal \N__52815\ : std_logic;
signal \N__52812\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52807\ : std_logic;
signal \N__52802\ : std_logic;
signal \N__52797\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52787\ : std_logic;
signal \N__52784\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52778\ : std_logic;
signal \N__52775\ : std_logic;
signal \N__52774\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52765\ : std_logic;
signal \N__52762\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52752\ : std_logic;
signal \N__52749\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52734\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52725\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52704\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52695\ : std_logic;
signal \N__52692\ : std_logic;
signal \N__52689\ : std_logic;
signal \N__52686\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52680\ : std_logic;
signal \N__52677\ : std_logic;
signal \N__52674\ : std_logic;
signal \N__52671\ : std_logic;
signal \N__52668\ : std_logic;
signal \N__52665\ : std_logic;
signal \N__52662\ : std_logic;
signal \N__52659\ : std_logic;
signal \N__52656\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52644\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52639\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52627\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52617\ : std_logic;
signal \N__52614\ : std_logic;
signal \N__52611\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52601\ : std_logic;
signal \N__52598\ : std_logic;
signal \N__52589\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52547\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52528\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52518\ : std_logic;
signal \N__52515\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52502\ : std_logic;
signal \N__52499\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52482\ : std_logic;
signal \N__52473\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52452\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52442\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52428\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52422\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52412\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52389\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52374\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52370\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52359\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52355\ : std_logic;
signal \N__52354\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52346\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52339\ : std_logic;
signal \N__52336\ : std_logic;
signal \N__52333\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52331\ : std_logic;
signal \N__52330\ : std_logic;
signal \N__52321\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52299\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52287\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52262\ : std_logic;
signal \N__52259\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52212\ : std_logic;
signal \N__52209\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52197\ : std_logic;
signal \N__52194\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52187\ : std_logic;
signal \N__52184\ : std_logic;
signal \N__52181\ : std_logic;
signal \N__52178\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52146\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52128\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52117\ : std_logic;
signal \N__52114\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52112\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52079\ : std_logic;
signal \N__52076\ : std_logic;
signal \N__52073\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52060\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52052\ : std_logic;
signal \N__52049\ : std_logic;
signal \N__52046\ : std_logic;
signal \N__52043\ : std_logic;
signal \N__52032\ : std_logic;
signal \N__52029\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52026\ : std_logic;
signal \N__52023\ : std_logic;
signal \N__52022\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52019\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52013\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52011\ : std_logic;
signal \N__52010\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__52007\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51998\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51995\ : std_logic;
signal \N__51994\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51989\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51961\ : std_logic;
signal \N__51960\ : std_logic;
signal \N__51959\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51949\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51944\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51940\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51929\ : std_logic;
signal \N__51926\ : std_logic;
signal \N__51925\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51898\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51884\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51877\ : std_logic;
signal \N__51876\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51872\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51869\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51864\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51862\ : std_logic;
signal \N__51861\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51799\ : std_logic;
signal \N__51796\ : std_logic;
signal \N__51793\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51761\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51731\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51719\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51671\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51656\ : std_logic;
signal \N__51655\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51650\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51644\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51641\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51632\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51611\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51599\ : std_logic;
signal \N__51596\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51575\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51573\ : std_logic;
signal \N__51572\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51533\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51512\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51429\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51416\ : std_logic;
signal \N__51413\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51407\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51384\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51381\ : std_logic;
signal \N__51378\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51357\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51350\ : std_logic;
signal \N__51347\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51333\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51302\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51278\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51195\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51177\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51173\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51156\ : std_logic;
signal \N__51155\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51108\ : std_logic;
signal \N__51107\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51091\ : std_logic;
signal \N__51088\ : std_logic;
signal \N__51083\ : std_logic;
signal \N__51078\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51072\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51068\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51046\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51035\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51019\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50987\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50959\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50920\ : std_logic;
signal \N__50917\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50902\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50862\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50854\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50840\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50832\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50792\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50783\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50752\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50732\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50729\ : std_logic;
signal \N__50726\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50702\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50671\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50644\ : std_logic;
signal \N__50639\ : std_logic;
signal \N__50630\ : std_logic;
signal \N__50627\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50080\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49601\ : std_logic;
signal \N__49598\ : std_logic;
signal \N__49595\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49556\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49310\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49265\ : std_logic;
signal \N__49262\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49172\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48899\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \ICE_GPMO_2\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\ : std_logic;
signal \ICE_SYSCLK\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\ : std_logic;
signal \RTD_SCLK\ : std_logic;
signal \RTD.n8\ : std_logic;
signal \RTD_SDI\ : std_logic;
signal \RTD.n11718\ : std_logic;
signal \RTD.n21_cascade_\ : std_logic;
signal \n13176_cascade_\ : std_logic;
signal n18755 : std_logic;
signal n13176 : std_logic;
signal \n18755_cascade_\ : std_logic;
signal \RTD.n16\ : std_logic;
signal \RTD.cfg_buf_6\ : std_logic;
signal cfg_buf_0 : std_logic;
signal \RTD.n9_cascade_\ : std_logic;
signal \RTD.adress_7_N_1339_7_cascade_\ : std_logic;
signal \RTD.cfg_buf_5\ : std_logic;
signal \RTD.cfg_buf_3\ : std_logic;
signal \RTD.n11_adj_1405\ : std_logic;
signal \RTD.cfg_buf_4\ : std_logic;
signal \RTD.cfg_buf_2\ : std_logic;
signal \RTD.n10\ : std_logic;
signal \RTD.adress_7\ : std_logic;
signal \RTD.n7318\ : std_logic;
signal \RTD.n7318_cascade_\ : std_logic;
signal \RTD.n4_cascade_\ : std_logic;
signal \RTD.cfg_buf_7\ : std_logic;
signal cfg_buf_1 : std_logic;
signal \RTD.n12\ : std_logic;
signal \RTD.n11\ : std_logic;
signal \RTD.n11_adj_1403\ : std_logic;
signal \RTD.n32\ : std_logic;
signal \RTD.n32_cascade_\ : std_logic;
signal \RTD.n21555\ : std_logic;
signal \RTD.n6\ : std_logic;
signal \RTD_SDO\ : std_logic;
signal \n1_adj_1606_cascade_\ : std_logic;
signal \RTD.n20160\ : std_logic;
signal read_buf_3 : std_logic;
signal read_buf_2 : std_logic;
signal \DDS_MCLK1\ : std_logic;
signal \RTD_CS\ : std_logic;
signal \RTD.n11687\ : std_logic;
signal adress_5 : std_logic;
signal adress_6 : std_logic;
signal \RTD.n19_cascade_\ : std_logic;
signal adress_0 : std_logic;
signal \n13165_cascade_\ : std_logic;
signal adress_1 : std_logic;
signal \n14479_cascade_\ : std_logic;
signal adress_4 : std_logic;
signal \RTD.n21362_cascade_\ : std_logic;
signal \RTD.n1\ : std_logic;
signal n14479 : std_logic;
signal adress_2 : std_logic;
signal n13165 : std_logic;
signal adress_3 : std_logic;
signal \RTD.mode\ : std_logic;
signal \RTD_DRDY\ : std_logic;
signal \RTD.adress_7_N_1339_7\ : std_logic;
signal \RTD.n16638\ : std_logic;
signal \RTD.n16638_cascade_\ : std_logic;
signal \RTD.n20787\ : std_logic;
signal \RTD.n17835\ : std_logic;
signal \RTD.n7\ : std_logic;
signal \RTD.n11726\ : std_logic;
signal \RTD.n19787\ : std_logic;
signal \RTD.n14_cascade_\ : std_logic;
signal \RTD.n20832\ : std_logic;
signal \RTD.n11704_cascade_\ : std_logic;
signal \RTD.cfg_tmp_1\ : std_logic;
signal \RTD.cfg_tmp_2\ : std_logic;
signal \RTD.cfg_tmp_3\ : std_logic;
signal \RTD.cfg_tmp_4\ : std_logic;
signal \RTD.cfg_tmp_5\ : std_logic;
signal \RTD.cfg_tmp_6\ : std_logic;
signal \RTD.cfg_tmp_7\ : std_logic;
signal \RTD.cfg_tmp_0\ : std_logic;
signal \RTD.n11704\ : std_logic;
signal \RTD.n14999\ : std_logic;
signal read_buf_4 : std_logic;
signal read_buf_0 : std_logic;
signal read_buf_1 : std_logic;
signal read_buf_5 : std_logic;
signal read_buf_6 : std_logic;
signal read_buf_12 : std_logic;
signal read_buf_14 : std_logic;
signal \VAC_MISO\ : std_logic;
signal cmd_rdadctmp_0_adj_1450 : std_logic;
signal cmd_rdadctmp_1_adj_1449 : std_logic;
signal \DDS_CS1\ : std_logic;
signal \CLK_DDS.n9_adj_1394\ : std_logic;
signal buf_adcdata_vac_5 : std_logic;
signal buf_adcdata_iac_5 : std_logic;
signal \n19_adj_1629_cascade_\ : std_logic;
signal buf_data_iac_6 : std_logic;
signal buf_adcdata_vac_4 : std_logic;
signal \n19_adj_1632_cascade_\ : std_logic;
signal buf_adcdata_iac_4 : std_logic;
signal buf_adcdata_iac_6 : std_logic;
signal n22_adj_1627 : std_logic;
signal cmd_rdadctmp_12 : std_logic;
signal cmd_rdadctmp_13 : std_logic;
signal \RTD.n17799\ : std_logic;
signal \RTD.bit_cnt_3\ : std_logic;
signal \RTD.bit_cnt_1\ : std_logic;
signal \RTD.bit_cnt_2\ : std_logic;
signal \RTD.bit_cnt_0\ : std_logic;
signal \RTD.n11740\ : std_logic;
signal \CLK_DDS.n16894\ : std_logic;
signal read_buf_15 : std_logic;
signal read_buf_7 : std_logic;
signal \buf_readRTD_10\ : std_logic;
signal n1_adj_1606 : std_logic;
signal n13293 : std_logic;
signal read_buf_10 : std_logic;
signal read_buf_11 : std_logic;
signal read_buf_13 : std_logic;
signal \buf_readRTD_13\ : std_logic;
signal read_buf_9 : std_logic;
signal \buf_readRTD_9\ : std_logic;
signal \buf_cfgRTD_1\ : std_logic;
signal \n14_adj_1610_cascade_\ : std_logic;
signal \VAC_CS\ : std_logic;
signal cmd_rdadctmp_14 : std_logic;
signal cmd_rdadctmp_2_adj_1448 : std_logic;
signal cmd_rdadctmp_3_adj_1447 : std_logic;
signal cmd_rdadctmp_4_adj_1446 : std_logic;
signal n20864 : std_logic;
signal \n20864_cascade_\ : std_logic;
signal \ADC_VAC.n17_cascade_\ : std_logic;
signal \ADC_VAC.n12\ : std_logic;
signal \IAC_CS\ : std_logic;
signal n14_adj_1612 : std_logic;
signal n20867 : std_logic;
signal \n20867_cascade_\ : std_logic;
signal \IAC_MISO\ : std_logic;
signal \n12498_cascade_\ : std_logic;
signal cmd_rdadctmp_0 : std_logic;
signal cmd_rdadctmp_1 : std_logic;
signal cmd_rdadctmp_2 : std_logic;
signal \AC_ADC_SYNC\ : std_logic;
signal buf_adcdata_vdc_5 : std_logic;
signal n19_adj_1626 : std_logic;
signal cmd_rdadctmp_16_adj_1434 : std_logic;
signal buf_data_iac_4 : std_logic;
signal n22_adj_1633 : std_logic;
signal bit_cnt_3 : std_logic;
signal n21456 : std_logic;
signal bit_cnt_1 : std_logic;
signal bit_cnt_2 : std_logic;
signal n8_adj_1602 : std_logic;
signal \CLK_DDS.n9\ : std_logic;
signal cmd_rdadctmp_13_adj_1437 : std_logic;
signal buf_adcdata_vac_8 : std_logic;
signal buf_adcdata_vac_6 : std_logic;
signal cmd_rdadctmp_14_adj_1436 : std_logic;
signal cmd_rdadctmp_15_adj_1435 : std_logic;
signal \buf_cfgRTD_2\ : std_logic;
signal \buf_cfgRTD_5\ : std_logic;
signal cmd_rdadctmp_24_adj_1426 : std_logic;
signal \n22321_cascade_\ : std_logic;
signal read_buf_8 : std_logic;
signal n11714 : std_logic;
signal \VAC_SCLK\ : std_logic;
signal cmd_rdadctmp_5_adj_1445 : std_logic;
signal cmd_rdadctmp_6_adj_1444 : std_logic;
signal \ADC_VAC.n21312\ : std_logic;
signal \ADC_VAC.n20958_cascade_\ : std_logic;
signal \ADC_VAC.n20959\ : std_logic;
signal \ADC_VDC.n19_cascade_\ : std_logic;
signal \ADC_VDC.n18563_cascade_\ : std_logic;
signal \ADC_VDC.n18563\ : std_logic;
signal \ADC_VDC.n21384_cascade_\ : std_logic;
signal \ADC_VDC.n13034\ : std_logic;
signal \ADC_VDC.avg_cnt_0\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \ADC_VDC.n19698\ : std_logic;
signal \ADC_VDC.n19699\ : std_logic;
signal \ADC_VDC.n19700\ : std_logic;
signal \ADC_VDC.n19701\ : std_logic;
signal \ADC_VDC.n19702\ : std_logic;
signal \ADC_VDC.n19703\ : std_logic;
signal \ADC_VDC.n19704\ : std_logic;
signal \ADC_VDC.n19705\ : std_logic;
signal \ADC_VDC.avg_cnt_8\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \ADC_VDC.avg_cnt_9\ : std_logic;
signal \ADC_VDC.n19706\ : std_logic;
signal \ADC_VDC.avg_cnt_10\ : std_logic;
signal \ADC_VDC.n19707\ : std_logic;
signal \ADC_VDC.n19708\ : std_logic;
signal \ADC_VDC.n13010_cascade_\ : std_logic;
signal \n12871_cascade_\ : std_logic;
signal cmd_rdadctmp_0_adj_1479 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_0\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal cmd_rdadctmp_1_adj_1478 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_1\ : std_logic;
signal \ADC_VDC.n19663\ : std_logic;
signal cmd_rdadctmp_2_adj_1477 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_2\ : std_logic;
signal \ADC_VDC.n19664\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_3\ : std_logic;
signal \ADC_VDC.n19665\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_4\ : std_logic;
signal \ADC_VDC.n19666\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_5\ : std_logic;
signal \ADC_VDC.n19667\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_6\ : std_logic;
signal \ADC_VDC.n19668\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_7\ : std_logic;
signal \ADC_VDC.n19669\ : std_logic;
signal \ADC_VDC.n19670\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_8\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_9\ : std_logic;
signal \ADC_VDC.n19671\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_10\ : std_logic;
signal \ADC_VDC.n19672\ : std_logic;
signal cmd_rdadctmp_11_adj_1468 : std_logic;
signal \ADC_VDC.n19673\ : std_logic;
signal \ADC_VDC.n19674\ : std_logic;
signal \ADC_VDC.n19675\ : std_logic;
signal \ADC_VDC.n19676\ : std_logic;
signal \ADC_VDC.n19677\ : std_logic;
signal \ADC_VDC.n19678\ : std_logic;
signal cmd_rdadcbuf_16 : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal cmd_rdadctmp_17_adj_1462 : std_logic;
signal \ADC_VDC.n19679\ : std_logic;
signal \ADC_VDC.n19680\ : std_logic;
signal \ADC_VDC.n19681\ : std_logic;
signal cmd_rdadctmp_20_adj_1459 : std_logic;
signal \ADC_VDC.n19682\ : std_logic;
signal cmd_rdadctmp_21_adj_1458 : std_logic;
signal \ADC_VDC.n19683\ : std_logic;
signal \ADC_VDC.n19684\ : std_logic;
signal \ADC_VDC.n19685\ : std_logic;
signal \ADC_VDC.n19686\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \ADC_VDC.n19687\ : std_logic;
signal \ADC_VDC.n19688\ : std_logic;
signal \ADC_VDC.n19689\ : std_logic;
signal \ADC_VDC.n19690\ : std_logic;
signal \ADC_VDC.n19691\ : std_logic;
signal \ADC_VDC.n19692\ : std_logic;
signal \ADC_VDC.n19693\ : std_logic;
signal \ADC_VDC.n19694\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \ADC_VDC.n19695\ : std_logic;
signal \ADC_VDC.n13010\ : std_logic;
signal \ADC_VDC.n14915\ : std_logic;
signal \ADC_VDC.n19696\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_35_N_1138_34\ : std_logic;
signal buf_adcdata_vac_16 : std_logic;
signal cmd_rdadctmp_3 : std_logic;
signal cmd_rdadctmp_27_adj_1423 : std_logic;
signal cmd_rdadctmp_28_adj_1422 : std_logic;
signal cmd_rdadctmp_29_adj_1421 : std_logic;
signal cmd_rdadctmp_7_adj_1443 : std_logic;
signal cmd_rdadctmp_31_adj_1419 : std_logic;
signal cmd_rdadctmp_30_adj_1420 : std_logic;
signal n22405 : std_logic;
signal buf_adcdata_vac_21 : std_logic;
signal n21097 : std_logic;
signal \buf_cfgRTD_4\ : std_logic;
signal \buf_readRTD_12\ : std_logic;
signal \buf_readRTD_4\ : std_logic;
signal \AMPV_POW\ : std_logic;
signal \n23_adj_1540_cascade_\ : std_logic;
signal n21123 : std_logic;
signal \EIS_SYNCCLK\ : std_logic;
signal \IAC_CLK\ : std_logic;
signal cmd_rdadctmp_15 : std_logic;
signal n21082 : std_logic;
signal n21201 : std_logic;
signal \n22315_cascade_\ : std_logic;
signal n22318 : std_logic;
signal cmd_rdadctmp_22 : std_logic;
signal \buf_readRTD_8\ : std_logic;
signal \buf_cfgRTD_0\ : std_logic;
signal n21202 : std_logic;
signal \VAC_OSR1\ : std_logic;
signal cmd_rdadctmp_16 : std_logic;
signal cmd_rdadctmp_17 : std_logic;
signal \VAC_DRDY\ : std_logic;
signal cmd_rdadctmp_18 : std_logic;
signal \IAC_SCLK\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \ADC_IAC.n19649\ : std_logic;
signal \ADC_IAC.n19650\ : std_logic;
signal \ADC_IAC.n19651\ : std_logic;
signal \ADC_IAC.n19652\ : std_logic;
signal \ADC_IAC.n19653\ : std_logic;
signal \ADC_IAC.n19654\ : std_logic;
signal \ADC_IAC.n19655\ : std_logic;
signal \ADC_IAC.n14806\ : std_logic;
signal \ADC_IAC.n17_cascade_\ : std_logic;
signal \ADC_IAC.n12\ : std_logic;
signal \ADC_VDC.avg_cnt_4\ : std_logic;
signal \ADC_VDC.avg_cnt_7\ : std_logic;
signal \ADC_VDC.avg_cnt_3\ : std_logic;
signal \ADC_VDC.avg_cnt_5\ : std_logic;
signal \ADC_VDC.n20\ : std_logic;
signal \ADC_VDC.avg_cnt_11\ : std_logic;
signal \ADC_VDC.avg_cnt_2\ : std_logic;
signal \ADC_VDC.avg_cnt_1\ : std_logic;
signal \ADC_VDC.avg_cnt_6\ : std_logic;
signal \ADC_VDC.n21\ : std_logic;
signal cmd_rdadcbuf_27 : std_logic;
signal buf_adcdata_vdc_16 : std_logic;
signal cmd_rdadcbuf_19 : std_logic;
signal buf_adcdata_vdc_8 : std_logic;
signal cmd_rdadcbuf_12 : std_logic;
signal cmd_rdadcbuf_13 : std_logic;
signal cmd_rdadctmp_14_adj_1465 : std_logic;
signal cmd_rdadctmp_3_adj_1476 : std_logic;
signal cmd_rdadctmp_4_adj_1475 : std_logic;
signal cmd_rdadctmp_8_adj_1471 : std_logic;
signal cmd_rdadcbuf_18 : std_logic;
signal cmd_rdadctmp_5_adj_1474 : std_logic;
signal cmd_rdadctmp_6_adj_1473 : std_logic;
signal cmd_rdadctmp_7_adj_1472 : std_logic;
signal cmd_rdadcbuf_15 : std_logic;
signal buf_adcdata_vdc_4 : std_logic;
signal cmd_rdadctmp_12_adj_1467 : std_logic;
signal cmd_rdadctmp_13_adj_1466 : std_logic;
signal cmd_rdadctmp_9_adj_1470 : std_logic;
signal cmd_rdadctmp_10_adj_1469 : std_logic;
signal cmd_rdadcbuf_14 : std_logic;
signal cmd_rdadctmp_15_adj_1464 : std_logic;
signal cmd_rdadctmp_16_adj_1463 : std_logic;
signal n12871 : std_logic;
signal cmd_rdadctmp_18_adj_1461 : std_logic;
signal cmd_rdadctmp_19_adj_1460 : std_logic;
signal cmd_rdadcbuf_25 : std_logic;
signal cmd_rdadcbuf_24 : std_logic;
signal cmd_rdadcbuf_17 : std_logic;
signal buf_adcdata_vdc_6 : std_logic;
signal cmd_rdadcbuf_23 : std_logic;
signal buf_adcdata_vdc_7 : std_logic;
signal buf_adcdata_vac_7 : std_logic;
signal cmd_rdadcbuf_20 : std_logic;
signal cmd_rdadcbuf_22 : std_logic;
signal cmd_rdadcbuf_28 : std_logic;
signal cmd_rdadcbuf_34 : std_logic;
signal buf_adcdata_vdc_23 : std_logic;
signal buf_adcdata_vac_23 : std_logic;
signal cmd_rdadcbuf_32 : std_logic;
signal buf_adcdata_vdc_21 : std_logic;
signal cmd_rdadcbuf_31 : std_logic;
signal cmd_rdadcbuf_30 : std_logic;
signal cmd_rdadcbuf_29 : std_logic;
signal cmd_rdadctmp_23_adj_1427 : std_logic;
signal cmd_rdadctmp_26_adj_1424 : std_logic;
signal buf_adcdata_vdc_17 : std_logic;
signal n22441 : std_logic;
signal cmd_rdadctmp_25_adj_1425 : std_logic;
signal buf_adcdata_vac_17 : std_logic;
signal buf_adcdata_iac_7 : std_logic;
signal n19_adj_1623 : std_logic;
signal buf_data_iac_7 : std_logic;
signal \n22_adj_1624_cascade_\ : std_logic;
signal bit_cnt_0_adj_1456 : std_logic;
signal cmd_rdadctmp_7 : std_logic;
signal \DDS_MOSI1\ : std_logic;
signal \buf_cfgRTD_3\ : std_logic;
signal \buf_readRTD_11\ : std_logic;
signal buf_adcdata_vdc_12 : std_logic;
signal n19_adj_1511 : std_logic;
signal buf_adcdata_vdc_13 : std_logic;
signal cmd_rdadctmp_21_adj_1429 : std_logic;
signal buf_adcdata_vac_13 : std_logic;
signal cmd_rdadctmp_22_adj_1428 : std_logic;
signal cmd_rdadctmp_20_adj_1430 : std_logic;
signal buf_adcdata_vac_12 : std_logic;
signal cmd_rdadctmp_23 : std_logic;
signal n22417 : std_logic;
signal buf_adcdata_vac_20 : std_logic;
signal buf_adcdata_vdc_20 : std_logic;
signal cmd_rdadctmp_20 : std_logic;
signal n21139 : std_logic;
signal n22291 : std_logic;
signal \n21138_cascade_\ : std_logic;
signal buf_adcdata_iac_21 : std_logic;
signal buf_adcdata_vac_19 : std_logic;
signal n22435 : std_logic;
signal buf_adcdata_vdc_19 : std_logic;
signal cmd_rdadctmp_31 : std_logic;
signal cmd_rdadctmp_29 : std_logic;
signal cmd_rdadctmp_30 : std_logic;
signal buf_adcdata_iac_23 : std_logic;
signal \VAC_FLT1\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \ADC_VAC.n19656\ : std_logic;
signal \ADC_VAC.n19657\ : std_logic;
signal \ADC_VAC.n19658\ : std_logic;
signal \ADC_VAC.n19659\ : std_logic;
signal \ADC_VAC.bit_cnt_5\ : std_logic;
signal \ADC_VAC.n19660\ : std_logic;
signal \ADC_VAC.n19661\ : std_logic;
signal \ADC_VAC.n19662\ : std_logic;
signal \ADC_IAC.n20960_cascade_\ : std_logic;
signal \ADC_IAC.n20961\ : std_logic;
signal \ADC_IAC.bit_cnt_2\ : std_logic;
signal \ADC_IAC.bit_cnt_5\ : std_logic;
signal \ADC_IAC.bit_cnt_3\ : std_logic;
signal \ADC_IAC.bit_cnt_4\ : std_logic;
signal \ADC_IAC.bit_cnt_1\ : std_logic;
signal \ADC_IAC.bit_cnt_7\ : std_logic;
signal \ADC_IAC.n21295_cascade_\ : std_logic;
signal \ADC_IAC.n21294\ : std_logic;
signal \ADC_VAC.bit_cnt_4\ : std_logic;
signal \ADC_VAC.bit_cnt_3\ : std_logic;
signal \ADC_VAC.bit_cnt_1\ : std_logic;
signal \ADC_VAC.bit_cnt_2\ : std_logic;
signal \ADC_VAC.bit_cnt_0\ : std_logic;
signal \ADC_VAC.bit_cnt_6\ : std_logic;
signal \ADC_VAC.n21029_cascade_\ : std_logic;
signal \ADC_VAC.bit_cnt_7\ : std_logic;
signal \ADC_VAC.n21043\ : std_logic;
signal \ADC_IAC.bit_cnt_6\ : std_logic;
signal \ADC_IAC.bit_cnt_0\ : std_logic;
signal \ADC_IAC.n16\ : std_logic;
signal acadc_trig : std_logic;
signal \INVacadc_trig_300C_net\ : std_logic;
signal \IAC_DRDY\ : std_logic;
signal \ADC_IAC.n12473\ : std_logic;
signal \ADC_VDC.n11676_cascade_\ : std_logic;
signal \VDC_SCLK\ : std_logic;
signal \comm_spi.iclk_N_763\ : std_logic;
signal cmd_rdadcbuf_33 : std_logic;
signal cmd_rdadcbuf_11 : std_logic;
signal cmd_rdadcbuf_21 : std_logic;
signal n13087 : std_logic;
signal \n13087_cascade_\ : std_logic;
signal cmd_rdadcbuf_26 : std_logic;
signal cmd_rdadctmp_22_adj_1457 : std_logic;
signal \ADC_VDC.cmd_rdadctmp_23\ : std_logic;
signal \ADC_VDC.n12899\ : std_logic;
signal \ADC_VDC.n20656\ : std_logic;
signal \comm_spi.n22860\ : std_logic;
signal \comm_spi.n22860_cascade_\ : std_logic;
signal \comm_spi.n14597\ : std_logic;
signal buf_adcdata_vdc_0 : std_logic;
signal \n19_adj_1484_cascade_\ : std_logic;
signal \n22_adj_1483_cascade_\ : std_logic;
signal buf_data_iac_0 : std_logic;
signal buf_adcdata_iac_0 : std_logic;
signal cmd_rdadctmp_8_adj_1442 : std_logic;
signal buf_adcdata_vac_0 : std_logic;
signal cmd_rdadctmp_8 : std_logic;
signal \INVcomm_spi.bit_cnt_3767__i3C_net\ : std_logic;
signal adc_state_2_adj_1481 : std_logic;
signal \RTD.adc_state_1\ : std_logic;
signal \RTD.adc_state_3\ : std_logic;
signal \RTD.adc_state_0\ : std_logic;
signal \RTD.n15065\ : std_logic;
signal \DDS_SCK1\ : std_logic;
signal buf_adcdata_vdc_18 : std_logic;
signal buf_adcdata_vac_18 : std_logic;
signal n21081 : std_logic;
signal cmd_rdadctmp_6 : std_logic;
signal cmd_rdadctmp_4 : std_logic;
signal cmd_rdadctmp_5 : std_logic;
signal \THERMOSTAT\ : std_logic;
signal \n11347_cascade_\ : std_logic;
signal n11919 : std_logic;
signal buf_control_7 : std_logic;
signal \CLK_DDS.tmp_buf_10\ : std_logic;
signal \CLK_DDS.tmp_buf_11\ : std_logic;
signal \CLK_DDS.tmp_buf_12\ : std_logic;
signal tmp_buf_15_adj_1455 : std_logic;
signal \CLK_DDS.tmp_buf_7\ : std_logic;
signal buf_dds1_8 : std_logic;
signal buf_dds1_13 : std_logic;
signal cmd_rdadctmp_24 : std_logic;
signal buf_adcdata_iac_16 : std_logic;
signal cmd_rdadctmp_26 : std_logic;
signal n12395 : std_logic;
signal cmd_rdadctmp_27 : std_logic;
signal cmd_rdadctmp_28 : std_logic;
signal n19_adj_1527 : std_logic;
signal \n22279_cascade_\ : std_logic;
signal n17_adj_1526 : std_logic;
signal n23_adj_1529 : std_logic;
signal \n22363_cascade_\ : std_logic;
signal n21285 : std_logic;
signal n22282 : std_logic;
signal \n22366_cascade_\ : std_logic;
signal buf_dds1_15 : std_logic;
signal n16_adj_1525 : std_logic;
signal adc_state_1_adj_1417 : std_logic;
signal \IAC_OSR0\ : std_logic;
signal \n12367_cascade_\ : std_logic;
signal \n16563_cascade_\ : std_logic;
signal n22255 : std_logic;
signal \iac_raw_buf_N_734\ : std_logic;
signal \INVeis_state_i0C_net\ : std_logic;
signal \ADC_VDC.n21952\ : std_logic;
signal \INVcomm_spi.MISO_48_12186_12187_resetC_net\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal n19746 : std_logic;
signal n19747 : std_logic;
signal n19748 : std_logic;
signal n19749 : std_logic;
signal \ICE_SPI_SCLK\ : std_logic;
signal \comm_spi.n14596\ : std_logic;
signal \comm_spi.iclk_N_762\ : std_logic;
signal buf_adcdata_vdc_2 : std_logic;
signal \n19_adj_1639_cascade_\ : std_logic;
signal buf_data_iac_5 : std_logic;
signal n22_adj_1630 : std_logic;
signal buf_adcdata_iac_2 : std_logic;
signal cmd_rdadctmp_9 : std_logic;
signal cmd_rdadctmp_10 : std_logic;
signal n12498 : std_logic;
signal buf_adcdata_vac_2 : std_logic;
signal buf_adcdata_vdc_3 : std_logic;
signal \comm_spi.bit_cnt_1\ : std_logic;
signal \comm_spi.bit_cnt_2\ : std_logic;
signal \comm_spi.bit_cnt_0\ : std_logic;
signal cmd_rdadctmp_11 : std_logic;
signal buf_adcdata_vac_3 : std_logic;
signal cmd_rdadctmp_10_adj_1440 : std_logic;
signal cmd_rdadctmp_11_adj_1439 : std_logic;
signal cmd_rdadctmp_12_adj_1438 : std_logic;
signal n22_adj_1640 : std_logic;
signal buf_data_iac_2 : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal n19750 : std_logic;
signal n19751 : std_logic;
signal n19752 : std_logic;
signal n19753 : std_logic;
signal n19754 : std_logic;
signal n19755 : std_logic;
signal n19756 : std_logic;
signal n19757 : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal n19758 : std_logic;
signal n19759 : std_logic;
signal n19760 : std_logic;
signal n19761 : std_logic;
signal n19762 : std_logic;
signal n19763 : std_logic;
signal n19764 : std_logic;
signal n19765 : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal n19766 : std_logic;
signal n19767 : std_logic;
signal n19768 : std_logic;
signal n19769 : std_logic;
signal n19770 : std_logic;
signal n19771 : std_logic;
signal buf_dds1_14 : std_logic;
signal \CLK_DDS.tmp_buf_13\ : std_logic;
signal \CLK_DDS.tmp_buf_14\ : std_logic;
signal \CLK_DDS.tmp_buf_0\ : std_logic;
signal \CLK_DDS.tmp_buf_1\ : std_logic;
signal \CLK_DDS.tmp_buf_2\ : std_logic;
signal \CLK_DDS.tmp_buf_3\ : std_logic;
signal \CLK_DDS.tmp_buf_4\ : std_logic;
signal \CLK_DDS.tmp_buf_5\ : std_logic;
signal \CLK_DDS.tmp_buf_6\ : std_logic;
signal \CLK_DDS.tmp_buf_8\ : std_logic;
signal \CLK_DDS.tmp_buf_9\ : std_logic;
signal data_count_0 : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal data_count_1 : std_logic;
signal n19586 : std_logic;
signal data_count_2 : std_logic;
signal n19587 : std_logic;
signal data_count_3 : std_logic;
signal n19588 : std_logic;
signal data_count_4 : std_logic;
signal n19589 : std_logic;
signal data_count_5 : std_logic;
signal n19590 : std_logic;
signal data_count_6 : std_logic;
signal n19591 : std_logic;
signal data_count_7 : std_logic;
signal n19592 : std_logic;
signal n19593 : std_logic;
signal \INVdata_count_i0_i0C_net\ : std_logic;
signal data_count_8 : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal n19594 : std_logic;
signal data_count_9 : std_logic;
signal \INVdata_count_i0_i8C_net\ : std_logic;
signal \SIG_DDS.tmp_buf_10\ : std_logic;
signal buf_dds0_5 : std_logic;
signal buf_dds0_14 : std_logic;
signal \SIG_DDS.tmp_buf_13\ : std_logic;
signal \SIG_DDS.tmp_buf_11\ : std_logic;
signal \SIG_DDS.tmp_buf_12\ : std_logic;
signal \SIG_DDS.tmp_buf_9\ : std_logic;
signal \SIG_DDS.tmp_buf_5\ : std_logic;
signal n16554 : std_logic;
signal \iac_raw_buf_N_736_cascade_\ : std_logic;
signal n17_adj_1622 : std_logic;
signal \n20826_cascade_\ : std_logic;
signal \INVeis_end_299C_net\ : std_logic;
signal eis_end : std_logic;
signal n26_adj_1530 : std_logic;
signal n21234 : std_logic;
signal n21 : std_logic;
signal \n30_adj_1604_cascade_\ : std_logic;
signal n31 : std_logic;
signal \DTRIG_N_918\ : std_logic;
signal adc_state_1 : std_logic;
signal \n14_adj_1509_cascade_\ : std_logic;
signal n26_adj_1508 : std_logic;
signal n18_adj_1609 : std_logic;
signal n20915 : std_logic;
signal n20985 : std_logic;
signal n16571 : std_logic;
signal \n13_cascade_\ : std_logic;
signal n21337 : std_logic;
signal \INVeis_state_i2C_net\ : std_logic;
signal n17507 : std_logic;
signal eis_state_0 : std_logic;
signal \n11_adj_1621_cascade_\ : std_logic;
signal n11744 : std_logic;
signal \eis_end_N_724\ : std_logic;
signal \ADC_VDC.n10119_cascade_\ : std_logic;
signal \ADC_VDC.n12807\ : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal n19739 : std_logic;
signal n19740 : std_logic;
signal n19741 : std_logic;
signal n19742 : std_logic;
signal n19743 : std_logic;
signal n19744 : std_logic;
signal n19745 : std_logic;
signal \INVdds0_mclkcnt_i7_3772__i0C_net\ : std_logic;
signal clk_cnt_0 : std_logic;
signal clk_cnt_4 : std_logic;
signal clk_cnt_2 : std_logic;
signal clk_cnt_1 : std_logic;
signal \n6_cascade_\ : std_logic;
signal clk_cnt_3 : std_logic;
signal n14714 : std_logic;
signal \n14714_cascade_\ : std_logic;
signal \clk_RTD\ : std_logic;
signal dds0_mclkcnt_3 : std_logic;
signal dds0_mclkcnt_5 : std_logic;
signal dds0_mclkcnt_1 : std_logic;
signal dds0_mclkcnt_4 : std_logic;
signal dds0_mclkcnt_2 : std_logic;
signal dds0_mclkcnt_0 : std_logic;
signal \n12_adj_1480_cascade_\ : std_logic;
signal dds0_mclkcnt_7 : std_logic;
signal \n20799_cascade_\ : std_logic;
signal n10 : std_logic;
signal \INVcomm_spi.imiso_83_12192_12193_resetC_net\ : std_logic;
signal \comm_spi.n14611\ : std_logic;
signal \INVcomm_spi.MISO_48_12186_12187_setC_net\ : std_logic;
signal \ADC_VAC.n12594\ : std_logic;
signal \DTRIG_N_918_adj_1451\ : std_logic;
signal \ADC_VAC.n14844\ : std_logic;
signal dds0_mclkcnt_6 : std_logic;
signal n20799 : std_logic;
signal \INVdds0_mclk_294C_net\ : std_logic;
signal secclk_cnt_6 : std_logic;
signal secclk_cnt_14 : std_logic;
signal secclk_cnt_10 : std_logic;
signal secclk_cnt_3 : std_logic;
signal secclk_cnt_15 : std_logic;
signal secclk_cnt_8 : std_logic;
signal secclk_cnt_1 : std_logic;
signal secclk_cnt_5 : std_logic;
signal secclk_cnt_16 : std_logic;
signal secclk_cnt_2 : std_logic;
signal secclk_cnt_7 : std_logic;
signal secclk_cnt_13 : std_logic;
signal n27_adj_1597 : std_logic;
signal \n26_adj_1575_cascade_\ : std_logic;
signal n25_adj_1574 : std_logic;
signal \n19856_cascade_\ : std_logic;
signal secclk_cnt_20 : std_logic;
signal n14715 : std_logic;
signal secclk_cnt_0 : std_logic;
signal secclk_cnt_18 : std_logic;
signal secclk_cnt_11 : std_logic;
signal secclk_cnt_4 : std_logic;
signal n28_adj_1505 : std_logic;
signal buf_adcdata_iac_3 : std_logic;
signal n19_adj_1636 : std_logic;
signal secclk_cnt_17 : std_logic;
signal secclk_cnt_9 : std_logic;
signal n10_adj_1601 : std_logic;
signal buf_data_iac_3 : std_logic;
signal n22_adj_1637 : std_logic;
signal cmd_rdadctmp_17_adj_1433 : std_logic;
signal n12653 : std_logic;
signal cmd_rdadctmp_19_adj_1431 : std_logic;
signal secclk_cnt_21 : std_logic;
signal secclk_cnt_19 : std_logic;
signal secclk_cnt_12 : std_logic;
signal secclk_cnt_22 : std_logic;
signal n14_adj_1599 : std_logic;
signal \comm_spi.n14610\ : std_logic;
signal \INVcomm_spi.imiso_83_12192_12193_setC_net\ : std_logic;
signal \buf_readRTD_14\ : std_logic;
signal \buf_cfgRTD_6\ : std_logic;
signal \buf_readRTD_15\ : std_logic;
signal \buf_cfgRTD_7\ : std_logic;
signal n20_adj_1528 : std_logic;
signal cmd_rdadctmp_19 : std_logic;
signal cmd_rdadctmp_25 : std_logic;
signal buf_adcdata_iac_22 : std_logic;
signal \VAC_FLT0\ : std_logic;
signal \VDC_RNG0\ : std_logic;
signal \SIG_DDS.n10\ : std_logic;
signal buf_dds1_10 : std_logic;
signal \SELIRNG0\ : std_logic;
signal buf_dds0_1 : std_logic;
signal \SIG_DDS.tmp_buf_0\ : std_logic;
signal \SIG_DDS.tmp_buf_1\ : std_logic;
signal \SIG_DDS.tmp_buf_2\ : std_logic;
signal \SIG_DDS.tmp_buf_14\ : std_logic;
signal buf_dds0_15 : std_logic;
signal \SIG_DDS.tmp_buf_3\ : std_logic;
signal \SIG_DDS.tmp_buf_4\ : std_logic;
signal buf_dds0_8 : std_logic;
signal \SIG_DDS.tmp_buf_8\ : std_logic;
signal \SIG_DDS.tmp_buf_6\ : std_logic;
signal buf_dds0_7 : std_logic;
signal \SIG_DDS.tmp_buf_7\ : std_logic;
signal \acadc_skipCount_12\ : std_logic;
signal \acadc_skipCount_10\ : std_logic;
signal \acadc_skipCount_13\ : std_logic;
signal n20 : std_logic;
signal acadc_dtrig_v : std_logic;
signal acadc_dtrig_i : std_logic;
signal n4_adj_1546 : std_logic;
signal n23_adj_1501 : std_logic;
signal n24_adj_1642 : std_logic;
signal \acadc_skipCount_15\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \INVacadc_skipcnt_i0_i0C_net\ : std_logic;
signal n21037 : std_logic;
signal n19610 : std_logic;
signal \n19610_THRU_CRY_0_THRU_CO\ : std_logic;
signal \n19610_THRU_CRY_1_THRU_CO\ : std_logic;
signal \n19610_THRU_CRY_2_THRU_CO\ : std_logic;
signal \n19610_THRU_CRY_3_THRU_CO\ : std_logic;
signal \n19610_THRU_CRY_4_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n19610_THRU_CRY_5_THRU_CO\ : std_logic;
signal \n19610_THRU_CRY_6_THRU_CO\ : std_logic;
signal acadc_skipcnt_1 : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal n19611 : std_logic;
signal acadc_skipcnt_3 : std_logic;
signal n19612 : std_logic;
signal acadc_skipcnt_4 : std_logic;
signal n19613 : std_logic;
signal acadc_skipcnt_5 : std_logic;
signal n19614 : std_logic;
signal n19615 : std_logic;
signal n19616 : std_logic;
signal acadc_skipcnt_8 : std_logic;
signal n19617 : std_logic;
signal n19618 : std_logic;
signal \INVacadc_skipcnt_i0_i1C_net\ : std_logic;
signal acadc_skipcnt_9 : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal acadc_skipcnt_10 : std_logic;
signal n19619 : std_logic;
signal acadc_skipcnt_11 : std_logic;
signal n19620 : std_logic;
signal acadc_skipcnt_12 : std_logic;
signal n19621 : std_logic;
signal acadc_skipcnt_13 : std_logic;
signal n19622 : std_logic;
signal acadc_skipcnt_14 : std_logic;
signal n19623 : std_logic;
signal n19624 : std_logic;
signal acadc_skipcnt_15 : std_logic;
signal \INVacadc_skipcnt_i0_i9C_net\ : std_logic;
signal n11654 : std_logic;
signal n14671 : std_logic;
signal \ADC_VDC.n17\ : std_logic;
signal \ADC_VDC.n4\ : std_logic;
signal \ADC_VDC.n7_adj_1398\ : std_logic;
signal \ADC_VDC.n7_adj_1398_cascade_\ : std_logic;
signal \ADC_VDC.n77\ : std_logic;
signal \ADC_VDC.n77_cascade_\ : std_logic;
signal \ADC_VDC.n12\ : std_logic;
signal \ADC_VDC.n20899\ : std_logic;
signal \ADC_VDC.n72_cascade_\ : std_logic;
signal \ADC_VDC.n31_cascade_\ : std_logic;
signal \ADC_VDC.n22195_cascade_\ : std_logic;
signal \ADC_VDC.n22198_cascade_\ : std_logic;
signal \ADC_VDC.n18566\ : std_logic;
signal \ADC_VDC.n20811\ : std_logic;
signal \ADC_VDC.n6_adj_1399_cascade_\ : std_logic;
signal \ADC_VDC.n10536\ : std_logic;
signal \ADC_VDC.n21229\ : std_logic;
signal \ADC_VDC.n47\ : std_logic;
signal \comm_spi.n14608\ : std_logic;
signal buf_adcdata_vdc_1 : std_logic;
signal buf_adcdata_iac_1 : std_logic;
signal \n19_adj_1491_cascade_\ : std_logic;
signal buf_data_iac_1 : std_logic;
signal \n22_adj_1488_cascade_\ : std_logic;
signal n30_adj_1506 : std_logic;
signal comm_buf_2_1 : std_logic;
signal \n22249_cascade_\ : std_logic;
signal n30_adj_1482 : std_logic;
signal n30_adj_1625 : std_logic;
signal comm_buf_2_7 : std_logic;
signal n30_adj_1628 : std_logic;
signal n30_adj_1631 : std_logic;
signal n30_adj_1634 : std_logic;
signal n30_adj_1638 : std_logic;
signal n30_adj_1641 : std_logic;
signal \n4_adj_1594_cascade_\ : std_logic;
signal comm_buf_2_3 : std_logic;
signal \n22387_cascade_\ : std_logic;
signal n21193 : std_logic;
signal \n22390_cascade_\ : std_logic;
signal \n4_adj_1587_cascade_\ : std_logic;
signal \n21175_cascade_\ : std_logic;
signal \n2358_cascade_\ : std_logic;
signal \n20850_cascade_\ : std_logic;
signal \n31_adj_1613_cascade_\ : std_logic;
signal n12085 : std_logic;
signal \n12085_cascade_\ : std_logic;
signal n14764 : std_logic;
signal \n12228_cascade_\ : std_logic;
signal comm_buf_6_7 : std_logic;
signal n20850 : std_logic;
signal n20852 : std_logic;
signal comm_buf_6_3 : std_logic;
signal buf_dds1_1 : std_logic;
signal cmd_rdadctmp_9_adj_1441 : std_logic;
signal buf_adcdata_vac_1 : std_logic;
signal n20853 : std_logic;
signal adc_state_0_adj_1418 : std_logic;
signal cmd_rdadctmp_18_adj_1432 : std_logic;
signal n9_adj_1416 : std_logic;
signal buf_dds1_0 : std_logic;
signal n22_adj_1615 : std_logic;
signal \n10717_cascade_\ : std_logic;
signal n21344 : std_logic;
signal buf_dds1_5 : std_logic;
signal buf_dds1_7 : std_logic;
signal \acadc_skipCount_14\ : std_logic;
signal buf_dds0_4 : std_logic;
signal buf_dds1_4 : std_logic;
signal buf_dds0_0 : std_logic;
signal req_data_cnt_13 : std_logic;
signal n19_adj_1607 : std_logic;
signal \n29_cascade_\ : std_logic;
signal n16_adj_1603 : std_logic;
signal n24 : std_logic;
signal \n21_adj_1492_cascade_\ : std_logic;
signal n30_adj_1618 : std_logic;
signal n20_adj_1617 : std_logic;
signal n10717 : std_logic;
signal req_data_cnt_12 : std_logic;
signal \acadc_skipCount_9\ : std_logic;
signal \n8_adj_1573_cascade_\ : std_logic;
signal eis_stop : std_logic;
signal req_data_cnt_9 : std_logic;
signal n22375 : std_logic;
signal n22381 : std_logic;
signal n22384 : std_logic;
signal n11396 : std_logic;
signal \DDS_SCK\ : std_logic;
signal \comm_spi.n14605\ : std_logic;
signal \comm_spi.n14604\ : std_logic;
signal \ICE_SPI_MISO\ : std_logic;
signal \ADC_VDC.n19_adj_1401\ : std_logic;
signal \ADC_VDC.n21323_cascade_\ : std_logic;
signal \ADC_VDC.n21320\ : std_logic;
signal \ADC_VDC.n20965\ : std_logic;
signal \ADC_VDC.n10_cascade_\ : std_logic;
signal \ADC_VDC.n20812\ : std_logic;
signal \ADC_VDC.n20784\ : std_logic;
signal \ADC_VDC.n17509\ : std_logic;
signal \ADC_VDC.n11265\ : std_logic;
signal \ADC_VDC.n6\ : std_logic;
signal \ADC_VDC.n11265_cascade_\ : std_logic;
signal \ADC_VDC.n15\ : std_logic;
signal \ADC_VDC.n15_cascade_\ : std_logic;
signal \ADC_VDC.n20996\ : std_logic;
signal dds_state_1_adj_1453 : std_logic;
signal dds_state_2_adj_1452 : std_logic;
signal dds_state_0_adj_1454 : std_logic;
signal \CLK_DDS.n12784\ : std_logic;
signal \comm_spi.n14607\ : std_logic;
signal \n21122_cascade_\ : std_logic;
signal n21120 : std_logic;
signal n11361 : std_logic;
signal \n7_adj_1616_cascade_\ : std_logic;
signal \comm_spi.bit_cnt_3\ : std_logic;
signal \comm_spi.n17036\ : std_logic;
signal \INVcomm_spi.data_valid_85C_net\ : std_logic;
signal n20858 : std_logic;
signal adc_state_0 : std_logic;
signal cmd_rdadctmp_21 : std_logic;
signal buf_data_iac_21 : std_logic;
signal n21124 : std_logic;
signal \comm_spi.n14603\ : std_logic;
signal \comm_spi.data_tx_7__N_774\ : std_logic;
signal comm_tx_buf_7 : std_logic;
signal \comm_spi.data_tx_7__N_766\ : std_logic;
signal n12228 : std_logic;
signal buf_adcdata_vdc_9 : std_logic;
signal buf_adcdata_vac_9 : std_logic;
signal comm_tx_buf_3 : std_logic;
signal \n16891_cascade_\ : std_logic;
signal \SIG_DDS.n21571\ : std_logic;
signal buf_adcdata_vdc_10 : std_logic;
signal buf_adcdata_vac_10 : std_logic;
signal \ICE_GPMI_0\ : std_logic;
signal n11385 : std_logic;
signal \n10_adj_1554_cascade_\ : std_logic;
signal n11850 : std_logic;
signal \n20914_cascade_\ : std_logic;
signal n21014 : std_logic;
signal n17_adj_1489 : std_logic;
signal \SIG_DDS.n9\ : std_logic;
signal n22_adj_1499 : std_logic;
signal n18 : std_logic;
signal req_data_cnt_14 : std_logic;
signal n23_adj_1614 : std_logic;
signal n10520 : std_logic;
signal req_data_cnt_15 : std_logic;
signal \n8_adj_1532_cascade_\ : std_logic;
signal \data_index_9_N_216_0\ : std_logic;
signal n8_adj_1532 : std_logic;
signal n11338 : std_logic;
signal \n11338_cascade_\ : std_logic;
signal \n8813_cascade_\ : std_logic;
signal data_index_0 : std_logic;
signal n7 : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal data_index_1 : std_logic;
signal n19625 : std_logic;
signal n19626 : std_logic;
signal n19627 : std_logic;
signal n19628 : std_logic;
signal n19629 : std_logic;
signal n19630 : std_logic;
signal n19631 : std_logic;
signal n19632 : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal n10598 : std_logic;
signal n19633 : std_logic;
signal n7_adj_1572 : std_logic;
signal n8_adj_1573 : std_logic;
signal \data_index_9_N_216_1\ : std_logic;
signal \DDS_RNG_0\ : std_logic;
signal tmp_buf_15 : std_logic;
signal \DDS_MOSI\ : std_logic;
signal \DDS_CS\ : std_logic;
signal \SIG_DDS.n9_adj_1393\ : std_logic;
signal \comm_spi.data_tx_7__N_795\ : std_logic;
signal \ADC_VDC.bit_cnt_0\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \ADC_VDC.bit_cnt_1\ : std_logic;
signal \ADC_VDC.n19772\ : std_logic;
signal \ADC_VDC.bit_cnt_2\ : std_logic;
signal \ADC_VDC.n19773\ : std_logic;
signal \ADC_VDC.bit_cnt_3\ : std_logic;
signal \ADC_VDC.n19774\ : std_logic;
signal \ADC_VDC.bit_cnt_4\ : std_logic;
signal \ADC_VDC.n19775\ : std_logic;
signal \ADC_VDC.bit_cnt_5\ : std_logic;
signal \ADC_VDC.n19776\ : std_logic;
signal \ADC_VDC.bit_cnt_6\ : std_logic;
signal \ADC_VDC.n19777\ : std_logic;
signal \ADC_VDC.n19778\ : std_logic;
signal \ADC_VDC.bit_cnt_7\ : std_logic;
signal \ADC_VDC.n18550\ : std_logic;
signal \comm_spi.data_tx_7__N_786\ : std_logic;
signal \n20944_cascade_\ : std_logic;
signal n20964 : std_logic;
signal n20962 : std_logic;
signal n3 : std_logic;
signal n20801 : std_logic;
signal n4_adj_1586 : std_logic;
signal \n20801_cascade_\ : std_logic;
signal n19902 : std_logic;
signal n22423 : std_logic;
signal \n2_adj_1581_cascade_\ : std_logic;
signal \n21370_cascade_\ : std_logic;
signal n21369 : std_logic;
signal n22426 : std_logic;
signal n14 : std_logic;
signal \n1264_cascade_\ : std_logic;
signal n4_adj_1643 : std_logic;
signal n1264 : std_logic;
signal n8_adj_1582 : std_logic;
signal \comm_state_3_N_420_3\ : std_logic;
signal \comm_state_3_N_420_3_cascade_\ : std_logic;
signal \n21435_cascade_\ : std_logic;
signal n20829 : std_logic;
signal \n20937_cascade_\ : std_logic;
signal n20939 : std_logic;
signal n19_adj_1522 : std_logic;
signal \buf_readRTD_1\ : std_logic;
signal buf_adcdata_iac_9 : std_logic;
signal \n22261_cascade_\ : std_logic;
signal n16_adj_1521 : std_logic;
signal \n26_adj_1523_cascade_\ : std_logic;
signal \acadc_skipCount_1\ : std_logic;
signal \n22411_cascade_\ : std_logic;
signal req_data_cnt_1 : std_logic;
signal n22264 : std_logic;
signal \n22414_cascade_\ : std_logic;
signal \n30_adj_1524_cascade_\ : std_logic;
signal comm_buf_1_1 : std_logic;
signal \comm_spi.n14623\ : std_logic;
signal \comm_spi.data_tx_7__N_770\ : std_logic;
signal \comm_spi.n14622\ : std_logic;
signal \comm_spi.n22857\ : std_logic;
signal eis_state_1 : std_logic;
signal n26_adj_1644 : std_logic;
signal n20893 : std_logic;
signal n21521 : std_logic;
signal n14_adj_1533 : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal n14_adj_1556 : std_logic;
signal data_idxvec_1 : std_logic;
signal n19634 : std_logic;
signal n14_adj_1555 : std_logic;
signal n19635 : std_logic;
signal n19636 : std_logic;
signal n14_adj_1553 : std_logic;
signal n19637 : std_logic;
signal n14_adj_1584 : std_logic;
signal n19638 : std_logic;
signal n19639 : std_logic;
signal n14_adj_1551 : std_logic;
signal n19640 : std_logic;
signal n19641 : std_logic;
signal n14_adj_1550 : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal n14_adj_1580 : std_logic;
signal n19642 : std_logic;
signal n14_adj_1579 : std_logic;
signal n19643 : std_logic;
signal n19644 : std_logic;
signal n14_adj_1577 : std_logic;
signal data_idxvec_12 : std_logic;
signal n19645 : std_logic;
signal n14_adj_1583 : std_logic;
signal data_idxvec_13 : std_logic;
signal n19646 : std_logic;
signal n14_adj_1576 : std_logic;
signal data_idxvec_14 : std_logic;
signal n19647 : std_logic;
signal n14_adj_1549 : std_logic;
signal n19648 : std_logic;
signal data_idxvec_15 : std_logic;
signal n12280 : std_logic;
signal \iac_raw_buf_N_736\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal data_cntvec_1 : std_logic;
signal n19595 : std_logic;
signal n19596 : std_logic;
signal n19597 : std_logic;
signal n19598 : std_logic;
signal n19599 : std_logic;
signal n19600 : std_logic;
signal n19601 : std_logic;
signal n19602 : std_logic;
signal \INVdata_cntvec_i0_i0C_net\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal n19603 : std_logic;
signal n19604 : std_logic;
signal n19605 : std_logic;
signal data_cntvec_12 : std_logic;
signal n19606 : std_logic;
signal data_cntvec_13 : std_logic;
signal n19607 : std_logic;
signal data_cntvec_14 : std_logic;
signal n19608 : std_logic;
signal n19609 : std_logic;
signal data_cntvec_15 : std_logic;
signal \INVdata_cntvec_i0_i8C_net\ : std_logic;
signal n13457 : std_logic;
signal n14647 : std_logic;
signal acadc_skipcnt_0 : std_logic;
signal acadc_skipcnt_6 : std_logic;
signal n17 : std_logic;
signal \n8_adj_1565_cascade_\ : std_logic;
signal data_index_6 : std_logic;
signal \data_index_9_N_216_3\ : std_logic;
signal n8_adj_1565 : std_logic;
signal n7_adj_1564 : std_logic;
signal \data_index_9_N_216_6\ : std_logic;
signal data_index_9 : std_logic;
signal n8_adj_1559 : std_logic;
signal n7_adj_1558 : std_logic;
signal \n8_adj_1559_cascade_\ : std_logic;
signal \data_index_9_N_216_9\ : std_logic;
signal n7_adj_1560 : std_logic;
signal \data_index_9_N_216_8\ : std_logic;
signal \data_index_9_N_216_7\ : std_logic;
signal \clk_16MHz\ : std_logic;
signal dds0_mclk : std_logic;
signal buf_control_6 : std_logic;
signal \DDS_MCLK\ : std_logic;
signal \comm_spi.n14619\ : std_logic;
signal \comm_spi.n22884\ : std_logic;
signal \comm_spi.n22884_cascade_\ : std_logic;
signal \comm_spi.n14593\ : std_logic;
signal \comm_spi.n14618\ : std_logic;
signal \comm_spi.data_tx_7__N_772\ : std_logic;
signal \comm_spi.data_tx_7__N_792\ : std_logic;
signal \comm_spi.n22881\ : std_logic;
signal \comm_spi.data_tx_7__N_789\ : std_logic;
signal \comm_spi.data_tx_7__N_771\ : std_logic;
signal \comm_spi.n22878\ : std_logic;
signal wdtick_cnt_2 : std_logic;
signal wdtick_cnt_0 : std_logic;
signal wdtick_cnt_1 : std_logic;
signal \TEST_LED\ : std_logic;
signal \comm_spi.n14627\ : std_logic;
signal \comm_spi.n22875\ : std_logic;
signal \comm_spi.n14626\ : std_logic;
signal n11741 : std_logic;
signal n20992 : std_logic;
signal \n9255_cascade_\ : std_logic;
signal n14737 : std_logic;
signal flagcntwd : std_logic;
signal n11390 : std_logic;
signal \n12336_cascade_\ : std_logic;
signal n20378 : std_logic;
signal comm_buf_2_4 : std_logic;
signal comm_buf_6_4 : std_logic;
signal \n21538_cascade_\ : std_logic;
signal n1_adj_1591 : std_logic;
signal \n22369_cascade_\ : std_logic;
signal n2_adj_1592 : std_logic;
signal n4_adj_1593 : std_logic;
signal \comm_spi.data_tx_7__N_783\ : std_logic;
signal comm_tx_buf_4 : std_logic;
signal \comm_spi.data_tx_7__N_769\ : std_logic;
signal comm_buf_2_2 : std_logic;
signal \n22393_cascade_\ : std_logic;
signal comm_buf_6_2 : std_logic;
signal \n4_adj_1595_cascade_\ : std_logic;
signal n22396 : std_logic;
signal \n21196_cascade_\ : std_logic;
signal comm_tx_buf_2 : std_logic;
signal comm_buf_6_1 : std_logic;
signal \n4_adj_1596_cascade_\ : std_logic;
signal n22252 : std_logic;
signal \n21052_cascade_\ : std_logic;
signal comm_tx_buf_1 : std_logic;
signal buf_data_vac_0 : std_logic;
signal buf_data_vac_7 : std_logic;
signal comm_buf_5_7 : std_logic;
signal buf_data_vac_6 : std_logic;
signal buf_data_vac_5 : std_logic;
signal buf_data_vac_4 : std_logic;
signal comm_buf_5_4 : std_logic;
signal buf_data_vac_3 : std_logic;
signal comm_buf_5_3 : std_logic;
signal buf_data_vac_2 : std_logic;
signal comm_buf_5_2 : std_logic;
signal buf_data_vac_1 : std_logic;
signal comm_buf_5_1 : std_logic;
signal \IAC_OSR1\ : std_logic;
signal buf_adcdata_iac_17 : std_logic;
signal buf_dds0_9 : std_logic;
signal \n22237_cascade_\ : std_logic;
signal buf_dds1_9 : std_logic;
signal buf_data_iac_17 : std_logic;
signal n22378 : std_logic;
signal \n21062_cascade_\ : std_logic;
signal n22240 : std_logic;
signal n22444 : std_logic;
signal \n22447_cascade_\ : std_logic;
signal \n22450_cascade_\ : std_logic;
signal comm_buf_0_1 : std_logic;
signal n30 : std_logic;
signal n21272 : std_logic;
signal n23_adj_1538 : std_logic;
signal \n22273_cascade_\ : std_logic;
signal n21286 : std_logic;
signal n17_adj_1535 : std_logic;
signal n16_adj_1534 : std_logic;
signal \n22288_cascade_\ : std_logic;
signal n22276 : std_logic;
signal \n30_adj_1539_cascade_\ : std_logic;
signal buf_adcdata_vdc_22 : std_logic;
signal buf_adcdata_vac_22 : std_logic;
signal n20_adj_1537 : std_logic;
signal \n19_adj_1536_cascade_\ : std_logic;
signal n22285 : std_logic;
signal buf_adcdata_iac_20 : std_logic;
signal buf_dds0_12 : std_logic;
signal \n22303_cascade_\ : std_logic;
signal buf_dds1_12 : std_logic;
signal n21309 : std_logic;
signal n23_adj_1541 : std_logic;
signal n21568 : std_logic;
signal n22243 : std_logic;
signal n22306 : std_logic;
signal n22420 : std_logic;
signal n22246 : std_logic;
signal \n21092_cascade_\ : std_logic;
signal \n30_adj_1542_cascade_\ : std_logic;
signal n21087 : std_logic;
signal \n22357_cascade_\ : std_logic;
signal \n22360_cascade_\ : std_logic;
signal \n21137_cascade_\ : std_logic;
signal n21072 : std_logic;
signal n22327 : std_logic;
signal n22330 : std_logic;
signal data_idxvec_11 : std_logic;
signal data_cntvec_11 : std_logic;
signal buf_data_iac_19 : std_logic;
signal \n26_adj_1544_cascade_\ : std_logic;
signal acadc_rst : std_logic;
signal req_data_cnt_10 : std_logic;
signal n21088 : std_logic;
signal req_data_cnt_6 : std_logic;
signal buf_dds1_6 : std_logic;
signal buf_dds0_6 : std_logic;
signal buf_adcdata_iac_18 : std_logic;
signal n21073 : std_logic;
signal n16891 : std_logic;
signal data_index_5 : std_logic;
signal data_idxvec_10 : std_logic;
signal data_cntvec_10 : std_logic;
signal n21150 : std_logic;
signal data_idxvec_9 : std_logic;
signal data_cntvec_9 : std_logic;
signal n21060 : std_logic;
signal n8_adj_1569 : std_logic;
signal n7_adj_1568 : std_logic;
signal data_index_3 : std_logic;
signal data_idxvec_8 : std_logic;
signal data_cntvec_8 : std_logic;
signal req_data_cnt_11 : std_logic;
signal \n8_adj_1571_cascade_\ : std_logic;
signal data_index_2 : std_logic;
signal buf_dds0_10 : std_logic;
signal n20907 : std_logic;
signal n12429 : std_logic;
signal \n9306_cascade_\ : std_logic;
signal buf_dds0_13 : std_logic;
signal acadc_skipcnt_7 : std_logic;
signal acadc_skipcnt_2 : std_logic;
signal n22 : std_logic;
signal n9 : std_logic;
signal n20912 : std_logic;
signal comm_buf_0_4 : std_logic;
signal \n12381_cascade_\ : std_logic;
signal \VAC_OSR0\ : std_logic;
signal \acadc_skipCount_6\ : std_logic;
signal dds_state_0 : std_logic;
signal dds_state_2 : std_logic;
signal trig_dds0 : std_logic;
signal \SIG_DDS.n12722\ : std_logic;
signal data_index_8 : std_logic;
signal n8_adj_1561 : std_logic;
signal n8_adj_1563 : std_logic;
signal n7_adj_1562 : std_logic;
signal data_index_7 : std_logic;
signal \SELIRNG1\ : std_logic;
signal \acadc_skipCount_11\ : std_logic;
signal n23_adj_1543 : std_logic;
signal n11915 : std_logic;
signal buf_data_iac_22 : std_logic;
signal n21273 : std_logic;
signal buf_data_iac_20 : std_logic;
signal n21569 : std_logic;
signal \comm_spi.n14592\ : std_logic;
signal \comm_spi.n14639\ : std_logic;
signal \comm_spi.data_tx_7__N_777\ : std_logic;
signal \comm_spi.data_tx_7__N_780\ : std_logic;
signal comm_buf_5_6 : std_logic;
signal \n22183_cascade_\ : std_logic;
signal comm_buf_5_0 : std_logic;
signal n4 : std_logic;
signal comm_buf_6_0 : std_logic;
signal n21211 : std_logic;
signal n1 : std_logic;
signal comm_buf_2_0 : std_logic;
signal n2 : std_logic;
signal comm_tx_buf_0 : std_logic;
signal \comm_spi.data_tx_7__N_773\ : std_logic;
signal \n17479_cascade_\ : std_logic;
signal comm_buf_6_5 : std_logic;
signal comm_buf_2_5 : std_logic;
signal n17480 : std_logic;
signal comm_buf_5_5 : std_logic;
signal n21212 : std_logic;
signal \n17482_cascade_\ : std_logic;
signal n22189 : std_logic;
signal comm_tx_buf_5 : std_logic;
signal buf_data_vac_8 : std_logic;
signal comm_buf_4_0 : std_logic;
signal buf_data_vac_15 : std_logic;
signal comm_buf_4_7 : std_logic;
signal buf_data_vac_14 : std_logic;
signal comm_buf_4_6 : std_logic;
signal buf_data_vac_13 : std_logic;
signal comm_buf_4_5 : std_logic;
signal buf_data_vac_12 : std_logic;
signal comm_buf_4_4 : std_logic;
signal buf_data_vac_11 : std_logic;
signal comm_buf_4_3 : std_logic;
signal buf_data_vac_10 : std_logic;
signal comm_buf_4_2 : std_logic;
signal buf_data_vac_9 : std_logic;
signal comm_buf_4_1 : std_logic;
signal \SIG_DDS.bit_cnt_3\ : std_logic;
signal bit_cnt_0 : std_logic;
signal \SIG_DDS.bit_cnt_1\ : std_logic;
signal \SIG_DDS.bit_cnt_2\ : std_logic;
signal dds_state_1 : std_logic;
signal n14884 : std_logic;
signal n12220 : std_logic;
signal \n12220_cascade_\ : std_logic;
signal n14785 : std_logic;
signal n14778 : std_logic;
signal n30_adj_1531 : std_logic;
signal comm_buf_0_7 : std_logic;
signal n22324 : std_logic;
signal comm_buf_0_5 : std_logic;
signal buf_adcdata_iac_8 : std_logic;
signal n16_adj_1487 : std_logic;
signal n19_adj_1486 : std_logic;
signal \buf_readRTD_0\ : std_logic;
signal n22213 : std_logic;
signal data_idxvec_0 : std_logic;
signal data_cntvec_0 : std_logic;
signal \n26_cascade_\ : std_logic;
signal \acadc_skipCount_0\ : std_logic;
signal \n22201_cascade_\ : std_logic;
signal req_data_cnt_0 : std_logic;
signal n22216 : std_logic;
signal \n22204_cascade_\ : std_logic;
signal \n30_adj_1485_cascade_\ : std_logic;
signal comm_buf_1_0 : std_logic;
signal buf_adcdata_iac_19 : std_logic;
signal buf_dds0_11 : std_logic;
signal \n22297_cascade_\ : std_logic;
signal buf_dds1_11 : std_logic;
signal n21076 : std_logic;
signal n22300 : std_logic;
signal \n22312_cascade_\ : std_logic;
signal eis_start : std_logic;
signal req_data_cnt_8 : std_logic;
signal n22294 : std_logic;
signal \n21071_cascade_\ : std_logic;
signal comm_buf_0_0 : std_logic;
signal n14750 : std_logic;
signal n22219 : std_logic;
signal \acadc_skipCount_8\ : std_logic;
signal n14_adj_1578 : std_logic;
signal n9_adj_1415 : std_logic;
signal buf_data_iac_16 : std_logic;
signal n21165 : std_logic;
signal \n21167_cascade_\ : std_logic;
signal n22222 : std_logic;
signal n21070 : std_logic;
signal n21084 : std_logic;
signal n21085 : std_logic;
signal n22309 : std_logic;
signal n12399 : std_logic;
signal comm_buf_0_3 : std_logic;
signal \IAC_FLT1\ : std_logic;
signal n20914 : std_logic;
signal trig_dds1 : std_logic;
signal n8_adj_1571 : std_logic;
signal n7_adj_1570 : std_logic;
signal \data_index_9_N_216_2\ : std_logic;
signal n11819 : std_logic;
signal n12381 : std_logic;
signal comm_buf_0_2 : std_logic;
signal \IAC_FLT0\ : std_logic;
signal wdtick_flag : std_logic;
signal buf_control_0 : std_logic;
signal \CONT_SD\ : std_logic;
signal \comm_spi.imosi_N_753\ : std_logic;
signal \comm_spi.n22872\ : std_logic;
signal \comm_spi.n14630\ : std_logic;
signal \comm_spi.n14631\ : std_logic;
signal \comm_spi.data_tx_7__N_768\ : std_logic;
signal \comm_spi.n22869\ : std_logic;
signal \comm_spi.n14634\ : std_logic;
signal \comm_spi.n14635\ : std_logic;
signal \comm_spi.n14638\ : std_logic;
signal \ADC_VDC.genclk.n21446_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n26\ : std_logic;
signal \ADC_VDC.genclk.n27\ : std_logic;
signal \ADC_VDC.genclk.n28_adj_1397\ : std_logic;
signal \comm_spi.data_tx_7__N_767\ : std_logic;
signal comm_buf_0_6 : std_logic;
signal \n1_adj_1588_cascade_\ : std_logic;
signal comm_tx_buf_6 : std_logic;
signal n12336 : std_logic;
signal n14799 : std_logic;
signal comm_buf_2_6 : std_logic;
signal n2_adj_1589 : std_logic;
signal comm_buf_6_6 : std_logic;
signal n4_adj_1590 : std_logic;
signal \n21539_cascade_\ : std_logic;
signal n22339 : std_logic;
signal buf_data_vac_16 : std_logic;
signal comm_buf_3_0 : std_logic;
signal buf_data_vac_20 : std_logic;
signal comm_buf_3_4 : std_logic;
signal buf_data_vac_23 : std_logic;
signal comm_buf_3_7 : std_logic;
signal buf_data_vac_22 : std_logic;
signal comm_buf_3_6 : std_logic;
signal buf_data_vac_21 : std_logic;
signal comm_buf_3_5 : std_logic;
signal buf_data_vac_19 : std_logic;
signal comm_buf_3_3 : std_logic;
signal buf_data_vac_18 : std_logic;
signal comm_buf_3_2 : std_logic;
signal comm_rx_buf_1 : std_logic;
signal buf_data_vac_17 : std_logic;
signal comm_buf_3_1 : std_logic;
signal n20878 : std_logic;
signal \n21352_cascade_\ : std_logic;
signal \n12_cascade_\ : std_logic;
signal n12136 : std_logic;
signal \n12136_cascade_\ : std_logic;
signal n14771 : std_logic;
signal n19783 : std_logic;
signal \n18991_cascade_\ : std_logic;
signal \n4_adj_1545_cascade_\ : std_logic;
signal n11961 : std_logic;
signal \n18993_cascade_\ : std_logic;
signal n12_adj_1605 : std_logic;
signal \n11991_cascade_\ : std_logic;
signal n14506 : std_logic;
signal n11896 : std_logic;
signal n10697 : std_logic;
signal n18993 : std_logic;
signal n20843 : std_logic;
signal \n12_adj_1635_cascade_\ : std_logic;
signal n20917 : std_logic;
signal n12178 : std_logic;
signal n21177 : std_logic;
signal \n22225_cascade_\ : std_logic;
signal data_idxvec_6 : std_logic;
signal data_cntvec_6 : std_logic;
signal buf_data_iac_14 : std_logic;
signal \n26_adj_1507_cascade_\ : std_logic;
signal n21178 : std_logic;
signal comm_rx_buf_6 : std_logic;
signal n22228 : std_logic;
signal buf_adcdata_vdc_14 : std_logic;
signal buf_adcdata_vac_14 : std_logic;
signal \n19_cascade_\ : std_logic;
signal \buf_readRTD_6\ : std_logic;
signal n21046 : std_logic;
signal n16_adj_1510 : std_logic;
signal buf_adcdata_iac_12 : std_logic;
signal n22231 : std_logic;
signal data_idxvec_4 : std_logic;
signal data_cntvec_4 : std_logic;
signal \n26_adj_1512_cascade_\ : std_logic;
signal \acadc_skipCount_4\ : std_logic;
signal \n22351_cascade_\ : std_logic;
signal req_data_cnt_4 : std_logic;
signal n22234 : std_logic;
signal \n22354_cascade_\ : std_logic;
signal comm_rx_buf_4 : std_logic;
signal \n30_adj_1513_cascade_\ : std_logic;
signal n19_adj_1518 : std_logic;
signal \buf_readRTD_2\ : std_logic;
signal buf_adcdata_iac_10 : std_logic;
signal \n22207_cascade_\ : std_logic;
signal req_data_cnt_2 : std_logic;
signal \n22429_cascade_\ : std_logic;
signal \acadc_skipCount_2\ : std_logic;
signal n22210 : std_logic;
signal \n22432_cascade_\ : std_logic;
signal comm_rx_buf_2 : std_logic;
signal \n30_adj_1520_cascade_\ : std_logic;
signal data_idxvec_2 : std_logic;
signal data_cntvec_2 : std_logic;
signal n26_adj_1519 : std_logic;
signal n14_adj_1585 : std_logic;
signal n8 : std_logic;
signal buf_adcdata_iac_14 : std_logic;
signal n16 : std_logic;
signal n21045 : std_logic;
signal req_data_cnt_7 : std_logic;
signal \acadc_skipCount_7\ : std_logic;
signal buf_dds1_3 : std_logic;
signal buf_dds0_3 : std_logic;
signal buf_dds1_2 : std_logic;
signal n16_adj_1517 : std_logic;
signal comm_buf_1_2 : std_logic;
signal n12367 : std_logic;
signal buf_dds0_2 : std_logic;
signal comm_buf_1_6 : std_logic;
signal n14_adj_1552 : std_logic;
signal comm_buf_1_4 : std_logic;
signal data_index_4 : std_logic;
signal n8813 : std_logic;
signal n8_adj_1567 : std_logic;
signal n7_adj_1566 : std_logic;
signal \data_index_9_N_216_4\ : std_logic;
signal \ADC_VDC.n11750\ : std_logic;
signal \VDC_SDO\ : std_logic;
signal \ADC_VDC.adc_state_0\ : std_logic;
signal \ADC_VDC.n62\ : std_logic;
signal adc_state_2 : std_logic;
signal adc_state_3 : std_logic;
signal \ADC_VDC.n62_cascade_\ : std_logic;
signal \ADC_VDC.adc_state_1\ : std_logic;
signal \ADC_VDC.n11\ : std_logic;
signal \ADC_VDC.genclk.t0off_0\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal \ADC_VDC.genclk.t0off_1\ : std_logic;
signal \ADC_VDC.genclk.n19709\ : std_logic;
signal \ADC_VDC.genclk.t0off_2\ : std_logic;
signal \ADC_VDC.genclk.n19710\ : std_logic;
signal \ADC_VDC.genclk.t0off_3\ : std_logic;
signal \ADC_VDC.genclk.n19711\ : std_logic;
signal \ADC_VDC.genclk.t0off_4\ : std_logic;
signal \ADC_VDC.genclk.n19712\ : std_logic;
signal \ADC_VDC.genclk.t0off_5\ : std_logic;
signal \ADC_VDC.genclk.n19713\ : std_logic;
signal \ADC_VDC.genclk.t0off_6\ : std_logic;
signal \ADC_VDC.genclk.n19714\ : std_logic;
signal \ADC_VDC.genclk.t0off_7\ : std_logic;
signal \ADC_VDC.genclk.n19715\ : std_logic;
signal \ADC_VDC.genclk.n19716\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i0C_net\ : std_logic;
signal \ADC_VDC.genclk.t0off_8\ : std_logic;
signal \bfn_19_8_0_\ : std_logic;
signal \ADC_VDC.genclk.t0off_9\ : std_logic;
signal \ADC_VDC.genclk.n19717\ : std_logic;
signal \ADC_VDC.genclk.t0off_10\ : std_logic;
signal \ADC_VDC.genclk.n19718\ : std_logic;
signal \ADC_VDC.genclk.t0off_11\ : std_logic;
signal \ADC_VDC.genclk.n19719\ : std_logic;
signal \ADC_VDC.genclk.t0off_12\ : std_logic;
signal \ADC_VDC.genclk.n19720\ : std_logic;
signal \ADC_VDC.genclk.t0off_13\ : std_logic;
signal \ADC_VDC.genclk.n19721\ : std_logic;
signal \ADC_VDC.genclk.t0off_14\ : std_logic;
signal \ADC_VDC.genclk.n19722\ : std_logic;
signal \ADC_VDC.genclk.n19723\ : std_logic;
signal \ADC_VDC.genclk.t0off_15\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.n11735\ : std_logic;
signal n14529 : std_logic;
signal n17815 : std_logic;
signal n23_adj_1620 : std_logic;
signal \n21_adj_1598_cascade_\ : std_logic;
signal n17564 : std_logic;
signal n2358 : std_logic;
signal n20856 : std_logic;
signal \n15_cascade_\ : std_logic;
signal n18_adj_1619 : std_logic;
signal n14130 : std_logic;
signal n20880 : std_logic;
signal \n20880_cascade_\ : std_logic;
signal n12_adj_1548 : std_logic;
signal \ICE_SPI_CE0\ : std_logic;
signal comm_data_vld : std_logic;
signal n18984 : std_logic;
signal comm_cmd_4 : std_logic;
signal comm_cmd_6 : std_logic;
signal comm_cmd_5 : std_logic;
signal n21546 : std_logic;
signal n12092 : std_logic;
signal n12219 : std_logic;
signal n9255 : std_logic;
signal \n11853_cascade_\ : std_logic;
signal n12226 : std_logic;
signal comm_state_0 : std_logic;
signal n18991 : std_logic;
signal n20804 : std_logic;
signal n21341 : std_logic;
signal \n21339_cascade_\ : std_logic;
signal n38_adj_1608 : std_logic;
signal n21054 : std_logic;
signal \n22267_cascade_\ : std_logic;
signal data_idxvec_7 : std_logic;
signal data_cntvec_7 : std_logic;
signal buf_data_iac_15 : std_logic;
signal \n26_adj_1502_cascade_\ : std_logic;
signal n21055 : std_logic;
signal comm_rx_buf_7 : std_logic;
signal n22270 : std_logic;
signal comm_buf_1_7 : std_logic;
signal buf_adcdata_vdc_15 : std_logic;
signal buf_adcdata_vac_15 : std_logic;
signal \n19_adj_1503_cascade_\ : std_logic;
signal \buf_readRTD_7\ : std_logic;
signal n21049 : std_logic;
signal \buf_readRTD_3\ : std_logic;
signal req_data_cnt_3 : std_logic;
signal \acadc_skipCount_3\ : std_logic;
signal \n21132_cascade_\ : std_logic;
signal n21127 : std_logic;
signal \n22333_cascade_\ : std_logic;
signal comm_rx_buf_3 : std_logic;
signal \n22336_cascade_\ : std_logic;
signal comm_buf_1_3 : std_logic;
signal buf_adcdata_vdc_11 : std_logic;
signal buf_adcdata_vac_11 : std_logic;
signal n19_adj_1515 : std_logic;
signal data_idxvec_3 : std_logic;
signal data_cntvec_3 : std_logic;
signal buf_data_iac_11 : std_logic;
signal \n26_adj_1516_cascade_\ : std_logic;
signal n21133 : std_logic;
signal \n21316_cascade_\ : std_logic;
signal comm_length_2 : std_logic;
signal comm_index_0 : std_logic;
signal comm_index_2 : std_logic;
signal n4_adj_1600 : std_logic;
signal \n4_adj_1600_cascade_\ : std_logic;
signal comm_index_1 : std_logic;
signal \n5_cascade_\ : std_logic;
signal comm_cmd_7 : std_logic;
signal n21888 : std_logic;
signal n21317 : std_logic;
signal buf_adcdata_iac_15 : std_logic;
signal n16_adj_1504 : std_logic;
signal n21048 : std_logic;
signal comm_rx_buf_5 : std_logic;
signal comm_state_1 : std_logic;
signal comm_buf_1_5 : std_logic;
signal n11991 : std_logic;
signal n14757 : std_logic;
signal n19_adj_1497 : std_logic;
signal \buf_readRTD_5\ : std_logic;
signal data_idxvec_5 : std_logic;
signal data_cntvec_5 : std_logic;
signal \n26_adj_1498_cascade_\ : std_logic;
signal req_data_cnt_5 : std_logic;
signal \n22345_cascade_\ : std_logic;
signal \acadc_skipCount_5\ : std_logic;
signal \n22348_cascade_\ : std_logic;
signal n30_adj_1500 : std_logic;
signal buf_adcdata_iac_11 : std_logic;
signal n16_adj_1514 : std_logic;
signal n21126 : std_logic;
signal buf_data_iac_10 : std_logic;
signal n21564 : std_logic;
signal buf_data_iac_8 : std_logic;
signal n21218 : std_logic;
signal buf_data_iac_23 : std_logic;
signal n21364 : std_logic;
signal \INVADC_VDC.genclk.div_state_i1C_net\ : std_logic;
signal \ADC_VDC.genclk.n6\ : std_logic;
signal \comm_spi.iclk\ : std_logic;
signal \ADC_VDC.genclk.n21444\ : std_logic;
signal \comm_spi.DOUT_7__N_747\ : std_logic;
signal \VDC_CLK\ : std_logic;
signal \INVADC_VDC.genclk.div_state_i0C_net\ : std_logic;
signal \comm_spi.n14614\ : std_logic;
signal \comm_spi.n14615\ : std_logic;
signal comm_rx_buf_0 : std_logic;
signal \comm_spi.n22866\ : std_logic;
signal \comm_spi.n22866_cascade_\ : std_logic;
signal \comm_spi.n14601\ : std_logic;
signal \comm_spi.imosi_cascade_\ : std_logic;
signal \comm_spi.DOUT_7__N_746\ : std_logic;
signal \ADC_VDC.genclk.div_state_0\ : std_logic;
signal \comm_spi.imosi\ : std_logic;
signal \comm_spi.n22863\ : std_logic;
signal \comm_spi.n14600\ : std_logic;
signal comm_clear : std_logic;
signal \ICE_SPI_MOSI\ : std_logic;
signal \comm_spi.imosi_N_752\ : std_logic;
signal comm_state_2 : std_logic;
signal comm_length_0 : std_logic;
signal comm_cmd_1 : std_logic;
signal comm_cmd_3 : std_logic;
signal comm_length_1 : std_logic;
signal \clk_32MHz\ : std_logic;
signal n11860 : std_logic;
signal n14655 : std_logic;
signal buf_data_iac_12 : std_logic;
signal n21451 : std_logic;
signal buf_data_iac_18 : std_logic;
signal n21151 : std_logic;
signal n16_adj_1496 : std_logic;
signal n22399 : std_logic;
signal buf_adcdata_iac_13 : std_logic;
signal comm_cmd_2 : std_logic;
signal n22402 : std_logic;
signal buf_data_iac_13 : std_logic;
signal n21350 : std_logic;
signal buf_data_iac_9 : std_logic;
signal comm_cmd_0 : std_logic;
signal n21529 : std_logic;
signal comm_state_3 : std_logic;
signal n17489 : std_logic;
signal n9306 : std_logic;
signal n17487 : std_logic;
signal \data_index_9_N_216_5\ : std_logic;
signal \bfn_22_7_0_\ : std_logic;
signal \ADC_VDC.genclk.n19724\ : std_logic;
signal \ADC_VDC.genclk.n19725\ : std_logic;
signal \ADC_VDC.genclk.n19726\ : std_logic;
signal \ADC_VDC.genclk.n19727\ : std_logic;
signal \ADC_VDC.genclk.n19728\ : std_logic;
signal \ADC_VDC.genclk.n19729\ : std_logic;
signal \ADC_VDC.genclk.n19730\ : std_logic;
signal \ADC_VDC.genclk.n19731\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i0C_net\ : std_logic;
signal \bfn_22_8_0_\ : std_logic;
signal \ADC_VDC.genclk.n19732\ : std_logic;
signal \ADC_VDC.genclk.n19733\ : std_logic;
signal \ADC_VDC.genclk.n19734\ : std_logic;
signal \ADC_VDC.genclk.n19735\ : std_logic;
signal \ADC_VDC.genclk.n19736\ : std_logic;
signal \ADC_VDC.genclk.n19737\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ADC_VDC.genclk.n19738\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.n15051\ : std_logic;
signal \ADC_VDC.genclk.t0on_6\ : std_logic;
signal \ADC_VDC.genclk.t0on_1\ : std_logic;
signal \ADC_VDC.genclk.t0on_4\ : std_logic;
signal \ADC_VDC.genclk.t0on_0\ : std_logic;
signal \ADC_VDC.genclk.n21449_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n21443\ : std_logic;
signal \ADC_VDC.genclk.t0on_12\ : std_logic;
signal \ADC_VDC.genclk.t0on_2\ : std_logic;
signal \ADC_VDC.genclk.t0on_7\ : std_logic;
signal \ADC_VDC.genclk.t0on_10\ : std_logic;
signal \ADC_VDC.genclk.n27_adj_1396\ : std_logic;
signal \ADC_VDC.genclk.t0on_3\ : std_logic;
signal \ADC_VDC.genclk.t0on_13\ : std_logic;
signal \ADC_VDC.genclk.t0on_5\ : std_logic;
signal \ADC_VDC.genclk.t0on_8\ : std_logic;
signal \ADC_VDC.genclk.n26_adj_1395\ : std_logic;
signal \ADC_VDC.genclk.div_state_1\ : std_logic;
signal \ADC_VDC.genclk.div_state_1__N_1274\ : std_logic;
signal \ADC_VDC.genclk.t0on_14\ : std_logic;
signal \ADC_VDC.genclk.t0on_9\ : std_logic;
signal \ADC_VDC.genclk.t0on_15\ : std_logic;
signal \ADC_VDC.genclk.t0on_11\ : std_logic;
signal \ADC_VDC.genclk.n28\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VAC_DRDY_wire\ : std_logic;
signal \IAC_FLT1_wire\ : std_logic;
signal \DDS_SCK_wire\ : std_logic;
signal \ICE_IOR_166_wire\ : std_logic;
signal \ICE_IOR_119_wire\ : std_logic;
signal \DDS_MOSI_wire\ : std_logic;
signal \VAC_MISO_wire\ : std_logic;
signal \DDS_MOSI1_wire\ : std_logic;
signal \ICE_IOR_146_wire\ : std_logic;
signal \VDC_CLK_wire\ : std_logic;
signal \ICE_IOT_222_wire\ : std_logic;
signal \IAC_CS_wire\ : std_logic;
signal \ICE_IOL_18B_wire\ : std_logic;
signal \ICE_IOL_13A_wire\ : std_logic;
signal \ICE_IOB_81_wire\ : std_logic;
signal \VAC_OSR1_wire\ : std_logic;
signal \IAC_MOSI_wire\ : std_logic;
signal \DDS_CS1_wire\ : std_logic;
signal \ICE_IOL_4B_wire\ : std_logic;
signal \ICE_IOB_94_wire\ : std_logic;
signal \VAC_CS_wire\ : std_logic;
signal \VAC_CLK_wire\ : std_logic;
signal \ICE_SPI_CE0_wire\ : std_logic;
signal \ICE_IOR_167_wire\ : std_logic;
signal \ICE_IOR_118_wire\ : std_logic;
signal \RTD_SDO_wire\ : std_logic;
signal \IAC_OSR0_wire\ : std_logic;
signal \VDC_SCLK_wire\ : std_logic;
signal \VAC_FLT1_wire\ : std_logic;
signal \ICE_SPI_MOSI_wire\ : std_logic;
signal \ICE_IOR_165_wire\ : std_logic;
signal \ICE_IOR_147_wire\ : std_logic;
signal \ICE_IOL_14A_wire\ : std_logic;
signal \ICE_IOL_13B_wire\ : std_logic;
signal \ICE_IOB_91_wire\ : std_logic;
signal \ICE_GPMO_0_wire\ : std_logic;
signal \DDS_RNG_0_wire\ : std_logic;
signal \VDC_RNG0_wire\ : std_logic;
signal \ICE_SPI_SCLK_wire\ : std_logic;
signal \ICE_IOR_152_wire\ : std_logic;
signal \ICE_IOL_12A_wire\ : std_logic;
signal \RTD_DRDY_wire\ : std_logic;
signal \ICE_SPI_MISO_wire\ : std_logic;
signal \ICE_IOT_177_wire\ : std_logic;
signal \ICE_IOR_141_wire\ : std_logic;
signal \ICE_IOB_80_wire\ : std_logic;
signal \ICE_IOB_102_wire\ : std_logic;
signal \ICE_GPMO_2_wire\ : std_logic;
signal \ICE_GPMI_0_wire\ : std_logic;
signal \IAC_MISO_wire\ : std_logic;
signal \VAC_OSR0_wire\ : std_logic;
signal \VAC_MOSI_wire\ : std_logic;
signal \TEST_LED_wire\ : std_logic;
signal \ICE_IOR_148_wire\ : std_logic;
signal \STAT_COMM_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \ICE_IOR_161_wire\ : std_logic;
signal \ICE_IOB_95_wire\ : std_logic;
signal \ICE_IOB_82_wire\ : std_logic;
signal \ICE_IOB_104_wire\ : std_logic;
signal \IAC_CLK_wire\ : std_logic;
signal \DDS_CS_wire\ : std_logic;
signal \SELIRNG0_wire\ : std_logic;
signal \RTD_SDI_wire\ : std_logic;
signal \ICE_IOT_221_wire\ : std_logic;
signal \ICE_IOT_197_wire\ : std_logic;
signal \DDS_MCLK_wire\ : std_logic;
signal \RTD_SCLK_wire\ : std_logic;
signal \RTD_CS_wire\ : std_logic;
signal \ICE_IOR_137_wire\ : std_logic;
signal \IAC_OSR1_wire\ : std_logic;
signal \VAC_FLT0_wire\ : std_logic;
signal \ICE_IOR_144_wire\ : std_logic;
signal \ICE_IOR_128_wire\ : std_logic;
signal \ICE_GPMO_1_wire\ : std_logic;
signal \IAC_SCLK_wire\ : std_logic;
signal \EIS_SYNCCLK_wire\ : std_logic;
signal \ICE_IOR_139_wire\ : std_logic;
signal \ICE_IOL_4A_wire\ : std_logic;
signal \VAC_SCLK_wire\ : std_logic;
signal \THERMOSTAT_wire\ : std_logic;
signal \ICE_IOR_164_wire\ : std_logic;
signal \ICE_IOB_103_wire\ : std_logic;
signal \AMPV_POW_wire\ : std_logic;
signal \VDC_SDO_wire\ : std_logic;
signal \ICE_IOT_174_wire\ : std_logic;
signal \ICE_IOR_140_wire\ : std_logic;
signal \ICE_IOB_96_wire\ : std_logic;
signal \CONT_SD_wire\ : std_logic;
signal \AC_ADC_SYNC_wire\ : std_logic;
signal \SELIRNG1_wire\ : std_logic;
signal \ICE_IOL_12B_wire\ : std_logic;
signal \ICE_IOR_160_wire\ : std_logic;
signal \ICE_IOR_136_wire\ : std_logic;
signal \DDS_MCLK1_wire\ : std_logic;
signal \ICE_IOT_198_wire\ : std_logic;
signal \ICE_IOT_173_wire\ : std_logic;
signal \IAC_DRDY_wire\ : std_logic;
signal \ICE_IOT_178_wire\ : std_logic;
signal \ICE_IOR_138_wire\ : std_logic;
signal \ICE_IOR_120_wire\ : std_logic;
signal \IAC_FLT0_wire\ : std_logic;
signal \DDS_SCK1_wire\ : std_logic;
signal \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \VAC_DRDY_wire\ <= VAC_DRDY;
    IAC_FLT1 <= \IAC_FLT1_wire\;
    DDS_SCK <= \DDS_SCK_wire\;
    \ICE_IOR_166_wire\ <= ICE_IOR_166;
    \ICE_IOR_119_wire\ <= ICE_IOR_119;
    DDS_MOSI <= \DDS_MOSI_wire\;
    \VAC_MISO_wire\ <= VAC_MISO;
    DDS_MOSI1 <= \DDS_MOSI1_wire\;
    \ICE_IOR_146_wire\ <= ICE_IOR_146;
    VDC_CLK <= \VDC_CLK_wire\;
    \ICE_IOT_222_wire\ <= ICE_IOT_222;
    IAC_CS <= \IAC_CS_wire\;
    \ICE_IOL_18B_wire\ <= ICE_IOL_18B;
    \ICE_IOL_13A_wire\ <= ICE_IOL_13A;
    \ICE_IOB_81_wire\ <= ICE_IOB_81;
    VAC_OSR1 <= \VAC_OSR1_wire\;
    IAC_MOSI <= \IAC_MOSI_wire\;
    DDS_CS1 <= \DDS_CS1_wire\;
    \ICE_IOL_4B_wire\ <= ICE_IOL_4B;
    \ICE_IOB_94_wire\ <= ICE_IOB_94;
    VAC_CS <= \VAC_CS_wire\;
    VAC_CLK <= \VAC_CLK_wire\;
    \ICE_SPI_CE0_wire\ <= ICE_SPI_CE0;
    \ICE_IOR_167_wire\ <= ICE_IOR_167;
    \ICE_IOR_118_wire\ <= ICE_IOR_118;
    \RTD_SDO_wire\ <= RTD_SDO;
    IAC_OSR0 <= \IAC_OSR0_wire\;
    VDC_SCLK <= \VDC_SCLK_wire\;
    VAC_FLT1 <= \VAC_FLT1_wire\;
    \ICE_SPI_MOSI_wire\ <= ICE_SPI_MOSI;
    \ICE_IOR_165_wire\ <= ICE_IOR_165;
    \ICE_IOR_147_wire\ <= ICE_IOR_147;
    \ICE_IOL_14A_wire\ <= ICE_IOL_14A;
    \ICE_IOL_13B_wire\ <= ICE_IOL_13B;
    \ICE_IOB_91_wire\ <= ICE_IOB_91;
    \ICE_GPMO_0_wire\ <= ICE_GPMO_0;
    DDS_RNG_0 <= \DDS_RNG_0_wire\;
    VDC_RNG0 <= \VDC_RNG0_wire\;
    \ICE_SPI_SCLK_wire\ <= ICE_SPI_SCLK;
    \ICE_IOR_152_wire\ <= ICE_IOR_152;
    \ICE_IOL_12A_wire\ <= ICE_IOL_12A;
    \RTD_DRDY_wire\ <= RTD_DRDY;
    ICE_SPI_MISO <= \ICE_SPI_MISO_wire\;
    \ICE_IOT_177_wire\ <= ICE_IOT_177;
    \ICE_IOR_141_wire\ <= ICE_IOR_141;
    \ICE_IOB_80_wire\ <= ICE_IOB_80;
    \ICE_IOB_102_wire\ <= ICE_IOB_102;
    \ICE_GPMO_2_wire\ <= ICE_GPMO_2;
    ICE_GPMI_0 <= \ICE_GPMI_0_wire\;
    \IAC_MISO_wire\ <= IAC_MISO;
    VAC_OSR0 <= \VAC_OSR0_wire\;
    VAC_MOSI <= \VAC_MOSI_wire\;
    TEST_LED <= \TEST_LED_wire\;
    \ICE_IOR_148_wire\ <= ICE_IOR_148;
    STAT_COMM <= \STAT_COMM_wire\;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    \ICE_IOR_161_wire\ <= ICE_IOR_161;
    \ICE_IOB_95_wire\ <= ICE_IOB_95;
    \ICE_IOB_82_wire\ <= ICE_IOB_82;
    \ICE_IOB_104_wire\ <= ICE_IOB_104;
    IAC_CLK <= \IAC_CLK_wire\;
    DDS_CS <= \DDS_CS_wire\;
    SELIRNG0 <= \SELIRNG0_wire\;
    RTD_SDI <= \RTD_SDI_wire\;
    \ICE_IOT_221_wire\ <= ICE_IOT_221;
    \ICE_IOT_197_wire\ <= ICE_IOT_197;
    DDS_MCLK <= \DDS_MCLK_wire\;
    RTD_SCLK <= \RTD_SCLK_wire\;
    RTD_CS <= \RTD_CS_wire\;
    \ICE_IOR_137_wire\ <= ICE_IOR_137;
    IAC_OSR1 <= \IAC_OSR1_wire\;
    VAC_FLT0 <= \VAC_FLT0_wire\;
    \ICE_IOR_144_wire\ <= ICE_IOR_144;
    \ICE_IOR_128_wire\ <= ICE_IOR_128;
    \ICE_GPMO_1_wire\ <= ICE_GPMO_1;
    IAC_SCLK <= \IAC_SCLK_wire\;
    \EIS_SYNCCLK_wire\ <= EIS_SYNCCLK;
    \ICE_IOR_139_wire\ <= ICE_IOR_139;
    \ICE_IOL_4A_wire\ <= ICE_IOL_4A;
    VAC_SCLK <= \VAC_SCLK_wire\;
    \THERMOSTAT_wire\ <= THERMOSTAT;
    \ICE_IOR_164_wire\ <= ICE_IOR_164;
    \ICE_IOB_103_wire\ <= ICE_IOB_103;
    AMPV_POW <= \AMPV_POW_wire\;
    \VDC_SDO_wire\ <= VDC_SDO;
    \ICE_IOT_174_wire\ <= ICE_IOT_174;
    \ICE_IOR_140_wire\ <= ICE_IOR_140;
    \ICE_IOB_96_wire\ <= ICE_IOB_96;
    CONT_SD <= \CONT_SD_wire\;
    AC_ADC_SYNC <= \AC_ADC_SYNC_wire\;
    SELIRNG1 <= \SELIRNG1_wire\;
    \ICE_IOL_12B_wire\ <= ICE_IOL_12B;
    \ICE_IOR_160_wire\ <= ICE_IOR_160;
    \ICE_IOR_136_wire\ <= ICE_IOR_136;
    DDS_MCLK1 <= \DDS_MCLK1_wire\;
    \ICE_IOT_198_wire\ <= ICE_IOT_198;
    \ICE_IOT_173_wire\ <= ICE_IOT_173;
    \IAC_DRDY_wire\ <= IAC_DRDY;
    \ICE_IOT_178_wire\ <= ICE_IOT_178;
    \ICE_IOR_138_wire\ <= ICE_IOR_138;
    \ICE_IOR_120_wire\ <= ICE_IOR_120;
    IAC_FLT0 <= \IAC_FLT0_wire\;
    DDS_SCK1 <= \DDS_SCK1_wire\;
    \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    buf_data_iac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(13);
    buf_data_vac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(9);
    buf_data_iac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(5);
    buf_data_vac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ <= '0'&\N__39015\&\N__38916\&\N__38829\&\N__38232\&\N__55983\&\N__47577\&\N__38352\&\N__45051\&\N__36435\&\N__36177\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ <= '0'&\N__29544\&\N__29655\&\N__29754\&\N__28701\&\N__28809\&\N__28920\&\N__29025\&\N__29133\&\N__29241\&\N__29352\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ <= '0'&'0'&\N__43230\&'0'&'0'&'0'&\N__25290\&'0'&'0'&'0'&\N__40716\&'0'&'0'&'0'&\N__27084\&'0';
    buf_data_iac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(13);
    buf_data_vac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(9);
    buf_data_iac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(5);
    buf_data_vac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ <= '0'&\N__38972\&\N__38873\&\N__38786\&\N__38192\&\N__55940\&\N__47531\&\N__38315\&\N__45008\&\N__36395\&\N__36137\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ <= '0'&\N__29507\&\N__29618\&\N__29714\&\N__28658\&\N__28769\&\N__28883\&\N__28994\&\N__29099\&\N__29204\&\N__29318\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ <= '0'&'0'&\N__37176\&'0'&'0'&'0'&\N__34941\&'0'&'0'&'0'&\N__43517\&'0'&'0'&'0'&\N__21576\&'0';
    buf_data_iac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(13);
    buf_data_vac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(9);
    buf_data_iac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(5);
    buf_data_vac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ <= '0'&\N__39033\&\N__38934\&\N__38847\&\N__38250\&\N__56001\&\N__47595\&\N__38370\&\N__45069\&\N__36453\&\N__36195\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ <= '0'&\N__29562\&\N__29673\&\N__29772\&\N__28719\&\N__28827\&\N__28938\&\N__29043\&\N__29151\&\N__29259\&\N__29370\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ <= '0'&'0'&\N__25002\&'0'&'0'&'0'&\N__22830\&'0'&'0'&'0'&\N__40386\&'0'&'0'&'0'&\N__25098\&'0';
    buf_data_iac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(13);
    buf_data_vac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(9);
    buf_data_iac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(5);
    buf_data_vac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ <= '0'&\N__38984\&\N__38885\&\N__38798\&\N__38204\&\N__55952\&\N__47543\&\N__38327\&\N__45020\&\N__36407\&\N__36149\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ <= '0'&\N__29519\&\N__29630\&\N__29726\&\N__28670\&\N__28781\&\N__28895\&\N__29001\&\N__29109\&\N__29216\&\N__29328\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ <= '0'&'0'&\N__52788\&'0'&'0'&'0'&\N__50921\&'0'&'0'&'0'&\N__46647\&'0'&'0'&'0'&\N__35961\&'0';
    buf_data_iac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(13);
    buf_data_vac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(9);
    buf_data_iac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(5);
    buf_data_vac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ <= '0'&\N__39039\&\N__38940\&\N__38853\&\N__38256\&\N__56007\&\N__47601\&\N__38376\&\N__45075\&\N__36459\&\N__36201\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ <= '0'&\N__29568\&\N__29679\&\N__29778\&\N__28725\&\N__28833\&\N__28944\&\N__29049\&\N__29157\&\N__29265\&\N__29376\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ <= '0'&'0'&\N__25164\&'0'&'0'&'0'&\N__24192\&'0'&'0'&'0'&\N__31938\&'0'&'0'&'0'&\N__40434\&'0';
    buf_data_iac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(13);
    buf_data_vac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(9);
    buf_data_iac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(5);
    buf_data_vac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ <= '0'&\N__38996\&\N__38897\&\N__38810\&\N__38214\&\N__55964\&\N__47555\&\N__38334\&\N__45032\&\N__36417\&\N__36159\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ <= '0'&\N__29526\&\N__29637\&\N__29736\&\N__28682\&\N__28791\&\N__28902\&\N__29007\&\N__29115\&\N__29223\&\N__29334\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ <= '0'&'0'&\N__53832\&'0'&'0'&'0'&\N__24927\&'0'&'0'&'0'&\N__46268\&'0'&'0'&'0'&\N__24861\&'0';
    buf_data_iac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(13);
    buf_data_vac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(9);
    buf_data_iac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(5);
    buf_data_vac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ <= '0'&\N__38987\&\N__38888\&\N__38801\&\N__38201\&\N__55955\&\N__47552\&\N__38318\&\N__45023\&\N__36404\&\N__36146\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ <= '0'&\N__29510\&\N__29621\&\N__29723\&\N__28673\&\N__28778\&\N__28886\&\N__28985\&\N__29096\&\N__29207\&\N__29315\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ <= '0'&'0'&\N__20463\&'0'&'0'&'0'&\N__20484\&'0'&'0'&'0'&\N__20406\&'0'&'0'&'0'&\N__20430\&'0';
    buf_data_iac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(13);
    buf_data_vac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(9);
    buf_data_iac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(5);
    buf_data_vac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ <= '0'&\N__39003\&\N__38904\&\N__38817\&\N__38220\&\N__55971\&\N__47565\&\N__38340\&\N__45039\&\N__36423\&\N__36165\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ <= '0'&\N__29532\&\N__29643\&\N__29742\&\N__28689\&\N__28797\&\N__28908\&\N__29013\&\N__29121\&\N__29229\&\N__29340\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ <= '0'&'0'&\N__52188\&'0'&'0'&'0'&\N__50220\&'0'&'0'&'0'&\N__47046\&'0'&'0'&'0'&\N__46353\&'0';
    buf_data_iac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(13);
    buf_data_vac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(9);
    buf_data_iac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(5);
    buf_data_vac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ <= '0'&\N__38999\&\N__38900\&\N__38813\&\N__38213\&\N__55967\&\N__47564\&\N__38330\&\N__45035\&\N__36416\&\N__36158\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ <= '0'&\N__29522\&\N__29633\&\N__29735\&\N__28685\&\N__28790\&\N__28898\&\N__28997\&\N__29108\&\N__29219\&\N__29327\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ <= '0'&'0'&\N__24834\&'0'&'0'&'0'&\N__24297\&'0'&'0'&'0'&\N__20649\&'0'&'0'&'0'&\N__21546\&'0';
    buf_data_iac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(13);
    buf_data_vac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(9);
    buf_data_iac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(5);
    buf_data_vac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ <= '0'&\N__39027\&\N__38928\&\N__38841\&\N__38244\&\N__55995\&\N__47589\&\N__38364\&\N__45063\&\N__36447\&\N__36189\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ <= '0'&\N__29556\&\N__29667\&\N__29766\&\N__28713\&\N__28821\&\N__28932\&\N__29037\&\N__29145\&\N__29253\&\N__29364\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ <= '0'&'0'&\N__31050\&'0'&'0'&'0'&\N__28371\&'0'&'0'&'0'&\N__28179\&'0'&'0'&'0'&\N__27897\&'0';
    buf_data_iac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(13);
    buf_data_vac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(9);
    buf_data_iac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(5);
    buf_data_vac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ <= '0'&\N__39009\&\N__38910\&\N__38823\&\N__38226\&\N__55977\&\N__47571\&\N__38346\&\N__45045\&\N__36429\&\N__36171\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ <= '0'&\N__29538\&\N__29649\&\N__29748\&\N__28695\&\N__28803\&\N__28914\&\N__29019\&\N__29127\&\N__29235\&\N__29346\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ <= '0'&'0'&\N__39768\&'0'&'0'&'0'&\N__24393\&'0'&'0'&'0'&\N__27348\&'0'&'0'&'0'&\N__22683\&'0';
    buf_data_iac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(13);
    buf_data_vac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(9);
    buf_data_iac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(5);
    buf_data_vac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ <= '0'&\N__39021\&\N__38922\&\N__38835\&\N__38238\&\N__55989\&\N__47583\&\N__38358\&\N__45057\&\N__36441\&\N__36183\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ <= '0'&\N__29550\&\N__29661\&\N__29760\&\N__28707\&\N__28815\&\N__28926\&\N__29031\&\N__29139\&\N__29247\&\N__29358\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ <= '0'&'0'&\N__32847\&'0'&'0'&'0'&\N__33717\&'0'&'0'&'0'&\N__26973\&'0'&'0'&'0'&\N__26907\&'0';

    \pll_main.zim_pll_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "101",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => OPEN,
            REFERENCECLK => \N__19206\,
            RESETB => \N__58564\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => \clk_16MHz\,
            DYNAMICDELAY => \pll_main.zim_pll_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \clk_32MHz\,
            SCLK => \GNDG0\
        );

    \iac_raw_buf_vac_raw_buf_merged2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54379\,
            RE => \N__58508\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            WE => \N__27730\
        );

    \iac_raw_buf_vac_raw_buf_merged7_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54437\,
            RE => \N__58607\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            WE => \N__27707\
        );

    \iac_raw_buf_vac_raw_buf_merged1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54299\,
            RE => \N__58359\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            WE => \N__27758\
        );

    \iac_raw_buf_vac_raw_buf_merged6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54435\,
            RE => \N__58585\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            WE => \N__27706\
        );

    \iac_raw_buf_vac_raw_buf_merged0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54284\,
            RE => \N__58507\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            WE => \N__27759\
        );

    \iac_raw_buf_vac_raw_buf_merged5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54433\,
            RE => \N__58566\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            WE => \N__27708\
        );

    \iac_raw_buf_vac_raw_buf_merged9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54337\,
            RE => \N__58584\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            WE => \N__27756\
        );

    \iac_raw_buf_vac_raw_buf_merged4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54425\,
            RE => \N__58565\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            WE => \N__27709\
        );

    \iac_raw_buf_vac_raw_buf_merged8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54311\,
            RE => \N__58560\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            WE => \N__27757\
        );

    \iac_raw_buf_vac_raw_buf_merged10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54325\,
            RE => \N__58424\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            WE => \N__27749\
        );

    \iac_raw_buf_vac_raw_buf_merged3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54406\,
            RE => \N__58509\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            WE => \N__27729\
        );

    \iac_raw_buf_vac_raw_buf_merged11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__54351\,
            RE => \N__58428\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            WE => \N__27748\
        );

    \ipInertedIOPad_VAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59563\,
            DIN => \N__59562\,
            DOUT => \N__59561\,
            PACKAGEPIN => \VAC_DRDY_wire\
        );

    \ipInertedIOPad_VAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59563\,
            PADOUT => \N__59562\,
            PADIN => \N__59561\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59554\,
            DIN => \N__59553\,
            DOUT => \N__59552\,
            PACKAGEPIN => \IAC_FLT1_wire\
        );

    \ipInertedIOPad_IAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59554\,
            PADOUT => \N__59553\,
            PADIN => \N__59552\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44121\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59545\,
            DIN => \N__59544\,
            DOUT => \N__59543\,
            PACKAGEPIN => \DDS_SCK_wire\
        );

    \ipInertedIOPad_DDS_SCK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59545\,
            PADOUT => \N__59544\,
            PADIN => \N__59543\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34197\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_166_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59536\,
            DIN => \N__59535\,
            DOUT => \N__59534\,
            PACKAGEPIN => \ICE_IOR_166_wire\
        );

    \ipInertedIOPad_ICE_IOR_166_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59536\,
            PADOUT => \N__59535\,
            PADIN => \N__59534\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_119_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59527\,
            DIN => \N__59526\,
            DOUT => \N__59525\,
            PACKAGEPIN => \ICE_IOR_119_wire\
        );

    \ipInertedIOPad_ICE_IOR_119_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59527\,
            PADOUT => \N__59526\,
            PADIN => \N__59525\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59518\,
            DIN => \N__59517\,
            DOUT => \N__59516\,
            PACKAGEPIN => \DDS_MOSI_wire\
        );

    \ipInertedIOPad_DDS_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59518\,
            PADOUT => \N__59517\,
            PADIN => \N__59516\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36762\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59509\,
            DIN => \N__59508\,
            DOUT => \N__59507\,
            PACKAGEPIN => \VAC_MISO_wire\
        );

    \ipInertedIOPad_VAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59509\,
            PADOUT => \N__59508\,
            PADIN => \N__59507\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59500\,
            DIN => \N__59499\,
            DOUT => \N__59498\,
            PACKAGEPIN => \DDS_MOSI1_wire\
        );

    \ipInertedIOPad_DDS_MOSI1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59500\,
            PADOUT => \N__59499\,
            PADIN => \N__59498\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24726\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_146_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59491\,
            DIN => \N__59490\,
            DOUT => \N__59489\,
            PACKAGEPIN => \ICE_IOR_146_wire\
        );

    \ipInertedIOPad_ICE_IOR_146_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59491\,
            PADOUT => \N__59490\,
            PADIN => \N__59489\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59482\,
            DIN => \N__59481\,
            DOUT => \N__59480\,
            PACKAGEPIN => \VDC_CLK_wire\
        );

    \ipInertedIOPad_VDC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59482\,
            PADOUT => \N__59481\,
            PADIN => \N__59480\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__53324\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_222_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59473\,
            DIN => \N__59472\,
            DOUT => \N__59471\,
            PACKAGEPIN => \ICE_IOT_222_wire\
        );

    \ipInertedIOPad_ICE_IOT_222_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59473\,
            PADOUT => \N__59472\,
            PADIN => \N__59471\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59464\,
            DIN => \N__59463\,
            DOUT => \N__59462\,
            PACKAGEPIN => \IAC_CS_wire\
        );

    \ipInertedIOPad_IAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59464\,
            PADOUT => \N__59463\,
            PADIN => \N__59462\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21213\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_18B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59455\,
            DIN => \N__59454\,
            DOUT => \N__59453\,
            PACKAGEPIN => \ICE_IOL_18B_wire\
        );

    \ipInertedIOPad_ICE_IOL_18B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59455\,
            PADOUT => \N__59454\,
            PADIN => \N__59453\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59446\,
            DIN => \N__59445\,
            DOUT => \N__59444\,
            PACKAGEPIN => \ICE_IOL_13A_wire\
        );

    \ipInertedIOPad_ICE_IOL_13A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59446\,
            PADOUT => \N__59445\,
            PADIN => \N__59444\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_81_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59437\,
            DIN => \N__59436\,
            DOUT => \N__59435\,
            PACKAGEPIN => \ICE_IOB_81_wire\
        );

    \ipInertedIOPad_ICE_IOB_81_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59437\,
            PADOUT => \N__59436\,
            PADIN => \N__59435\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59428\,
            DIN => \N__59427\,
            DOUT => \N__59426\,
            PACKAGEPIN => \VAC_OSR1_wire\
        );

    \ipInertedIOPad_VAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59428\,
            PADOUT => \N__59427\,
            PADIN => \N__59426\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23187\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59419\,
            DIN => \N__59418\,
            DOUT => \N__59417\,
            PACKAGEPIN => \IAC_MOSI_wire\
        );

    \ipInertedIOPad_IAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59419\,
            PADOUT => \N__59418\,
            PADIN => \N__59417\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59410\,
            DIN => \N__59409\,
            DOUT => \N__59408\,
            PACKAGEPIN => \DDS_CS1_wire\
        );

    \ipInertedIOPad_DDS_CS1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59410\,
            PADOUT => \N__59409\,
            PADIN => \N__59408\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20304\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59401\,
            DIN => \N__59400\,
            DOUT => \N__59399\,
            PACKAGEPIN => \ICE_IOL_4B_wire\
        );

    \ipInertedIOPad_ICE_IOL_4B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59401\,
            PADOUT => \N__59400\,
            PADIN => \N__59399\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_94_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59392\,
            DIN => \N__59391\,
            DOUT => \N__59390\,
            PACKAGEPIN => \ICE_IOB_94_wire\
        );

    \ipInertedIOPad_ICE_IOB_94_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59392\,
            PADOUT => \N__59391\,
            PADIN => \N__59390\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59383\,
            DIN => \N__59382\,
            DOUT => \N__59381\,
            PACKAGEPIN => \VAC_CS_wire\
        );

    \ipInertedIOPad_VAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59383\,
            PADOUT => \N__59382\,
            PADIN => \N__59381\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21126\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59374\,
            DIN => \N__59373\,
            DOUT => \N__59372\,
            PACKAGEPIN => \VAC_CLK_wire\
        );

    \ipInertedIOPad_VAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59374\,
            PADOUT => \N__59373\,
            PADIN => \N__59372\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22998\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_CE0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59365\,
            DIN => \N__59364\,
            DOUT => \N__59363\,
            PACKAGEPIN => \ICE_SPI_CE0_wire\
        );

    \ipInertedIOPad_ICE_SPI_CE0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59365\,
            PADOUT => \N__59364\,
            PADIN => \N__59363\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_CE0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_167_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59356\,
            DIN => \N__59355\,
            DOUT => \N__59354\,
            PACKAGEPIN => \ICE_IOR_167_wire\
        );

    \ipInertedIOPad_ICE_IOR_167_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59356\,
            PADOUT => \N__59355\,
            PADIN => \N__59354\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_118_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59347\,
            DIN => \N__59346\,
            DOUT => \N__59345\,
            PACKAGEPIN => \ICE_IOR_118_wire\
        );

    \ipInertedIOPad_ICE_IOR_118_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59347\,
            PADOUT => \N__59346\,
            PADIN => \N__59345\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDO_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59338\,
            DIN => \N__59337\,
            DOUT => \N__59336\,
            PACKAGEPIN => \RTD_SDO_wire\
        );

    \ipInertedIOPad_RTD_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59338\,
            PADOUT => \N__59337\,
            PADIN => \N__59336\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59329\,
            DIN => \N__59328\,
            DOUT => \N__59327\,
            PACKAGEPIN => \IAC_OSR0_wire\
        );

    \ipInertedIOPad_IAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59329\,
            PADOUT => \N__59328\,
            PADIN => \N__59327\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27636\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59320\,
            DIN => \N__59319\,
            DOUT => \N__59318\,
            PACKAGEPIN => \VDC_SCLK_wire\
        );

    \ipInertedIOPad_VDC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59320\,
            PADOUT => \N__59319\,
            PADIN => \N__59318\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25851\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59311\,
            DIN => \N__59310\,
            DOUT => \N__59309\,
            PACKAGEPIN => \VAC_FLT1_wire\
        );

    \ipInertedIOPad_VAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59311\,
            PADOUT => \N__59310\,
            PADIN => \N__59309\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25365\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MOSI_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59302\,
            DIN => \N__59301\,
            DOUT => \N__59300\,
            PACKAGEPIN => \ICE_SPI_MOSI_wire\
        );

    \ipInertedIOPad_ICE_SPI_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59302\,
            PADOUT => \N__59301\,
            PADIN => \N__59300\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_MOSI\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_165_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59293\,
            DIN => \N__59292\,
            DOUT => \N__59291\,
            PACKAGEPIN => \ICE_IOR_165_wire\
        );

    \ipInertedIOPad_ICE_IOR_165_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59293\,
            PADOUT => \N__59292\,
            PADIN => \N__59291\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_147_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59284\,
            DIN => \N__59283\,
            DOUT => \N__59282\,
            PACKAGEPIN => \ICE_IOR_147_wire\
        );

    \ipInertedIOPad_ICE_IOR_147_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59284\,
            PADOUT => \N__59283\,
            PADIN => \N__59282\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_14A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59275\,
            DIN => \N__59274\,
            DOUT => \N__59273\,
            PACKAGEPIN => \ICE_IOL_14A_wire\
        );

    \ipInertedIOPad_ICE_IOL_14A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59275\,
            PADOUT => \N__59274\,
            PADIN => \N__59273\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59266\,
            DIN => \N__59265\,
            DOUT => \N__59264\,
            PACKAGEPIN => \ICE_IOL_13B_wire\
        );

    \ipInertedIOPad_ICE_IOL_13B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59266\,
            PADOUT => \N__59265\,
            PADIN => \N__59264\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_91_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59257\,
            DIN => \N__59256\,
            DOUT => \N__59255\,
            PACKAGEPIN => \ICE_IOB_91_wire\
        );

    \ipInertedIOPad_ICE_IOB_91_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59257\,
            PADOUT => \N__59256\,
            PADIN => \N__59255\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59248\,
            DIN => \N__59247\,
            DOUT => \N__59246\,
            PACKAGEPIN => \ICE_GPMO_0_wire\
        );

    \ipInertedIOPad_ICE_GPMO_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59248\,
            PADOUT => \N__59247\,
            PADIN => \N__59246\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_RNG_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59239\,
            DIN => \N__59238\,
            DOUT => \N__59237\,
            PACKAGEPIN => \DDS_RNG_0_wire\
        );

    \ipInertedIOPad_DDS_RNG_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59239\,
            PADOUT => \N__59238\,
            PADIN => \N__59237\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36365\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_RNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59230\,
            DIN => \N__59229\,
            DOUT => \N__59228\,
            PACKAGEPIN => \VDC_RNG0_wire\
        );

    \ipInertedIOPad_VDC_RNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59230\,
            PADOUT => \N__59229\,
            PADIN => \N__59228\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31866\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_SCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59221\,
            DIN => \N__59220\,
            DOUT => \N__59219\,
            PACKAGEPIN => \ICE_SPI_SCLK_wire\
        );

    \ipInertedIOPad_ICE_SPI_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59221\,
            PADOUT => \N__59220\,
            PADIN => \N__59219\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_SCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_152_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59212\,
            DIN => \N__59211\,
            DOUT => \N__59210\,
            PACKAGEPIN => \ICE_IOR_152_wire\
        );

    \ipInertedIOPad_ICE_IOR_152_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59212\,
            PADOUT => \N__59211\,
            PADIN => \N__59210\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59203\,
            DIN => \N__59202\,
            DOUT => \N__59201\,
            PACKAGEPIN => \ICE_IOL_12A_wire\
        );

    \ipInertedIOPad_ICE_IOL_12A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59203\,
            PADOUT => \N__59202\,
            PADIN => \N__59201\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_DRDY_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59194\,
            DIN => \N__59193\,
            DOUT => \N__59192\,
            PACKAGEPIN => \RTD_DRDY_wire\
        );

    \ipInertedIOPad_RTD_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59194\,
            PADOUT => \N__59193\,
            PADIN => \N__59192\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59185\,
            DIN => \N__59184\,
            DOUT => \N__59183\,
            PACKAGEPIN => \ICE_SPI_MISO_wire\
        );

    \ipInertedIOPad_ICE_SPI_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59185\,
            PADOUT => \N__59184\,
            PADIN => \N__59183\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34143\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_177_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59176\,
            DIN => \N__59175\,
            DOUT => \N__59174\,
            PACKAGEPIN => \ICE_IOT_177_wire\
        );

    \ipInertedIOPad_ICE_IOT_177_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59176\,
            PADOUT => \N__59175\,
            PADIN => \N__59174\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_141_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59167\,
            DIN => \N__59166\,
            DOUT => \N__59165\,
            PACKAGEPIN => \ICE_IOR_141_wire\
        );

    \ipInertedIOPad_ICE_IOR_141_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59167\,
            PADOUT => \N__59166\,
            PADIN => \N__59165\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_80_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59158\,
            DIN => \N__59157\,
            DOUT => \N__59156\,
            PACKAGEPIN => \ICE_IOB_80_wire\
        );

    \ipInertedIOPad_ICE_IOB_80_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59158\,
            PADOUT => \N__59157\,
            PADIN => \N__59156\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_102_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59149\,
            DIN => \N__59148\,
            DOUT => \N__59147\,
            PACKAGEPIN => \ICE_IOB_102_wire\
        );

    \ipInertedIOPad_ICE_IOB_102_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59149\,
            PADOUT => \N__59148\,
            PADIN => \N__59147\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59140\,
            DIN => \N__59139\,
            DOUT => \N__59138\,
            PACKAGEPIN => \ICE_GPMO_2_wire\
        );

    \ipInertedIOPad_ICE_GPMO_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59140\,
            PADOUT => \N__59139\,
            PADIN => \N__59138\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMI_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59131\,
            DIN => \N__59130\,
            DOUT => \N__59129\,
            PACKAGEPIN => \ICE_GPMI_0_wire\
        );

    \ipInertedIOPad_ICE_GPMI_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59131\,
            PADOUT => \N__59130\,
            PADIN => \N__59129\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__35928\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59122\,
            DIN => \N__59121\,
            DOUT => \N__59120\,
            PACKAGEPIN => \IAC_MISO_wire\
        );

    \ipInertedIOPad_IAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59122\,
            PADOUT => \N__59121\,
            PADIN => \N__59120\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59113\,
            DIN => \N__59112\,
            DOUT => \N__59111\,
            PACKAGEPIN => \VAC_OSR0_wire\
        );

    \ipInertedIOPad_VAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59113\,
            PADOUT => \N__59112\,
            PADIN => \N__59111\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__41400\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59104\,
            DIN => \N__59103\,
            DOUT => \N__59102\,
            PACKAGEPIN => \VAC_MOSI_wire\
        );

    \ipInertedIOPad_VAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59104\,
            PADOUT => \N__59103\,
            PADIN => \N__59102\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TEST_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59095\,
            DIN => \N__59094\,
            DOUT => \N__59093\,
            PACKAGEPIN => \TEST_LED_wire\
        );

    \ipInertedIOPad_TEST_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59095\,
            PADOUT => \N__59094\,
            PADIN => \N__59093\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__39207\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_148_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59086\,
            DIN => \N__59085\,
            DOUT => \N__59084\,
            PACKAGEPIN => \ICE_IOR_148_wire\
        );

    \ipInertedIOPad_ICE_IOR_148_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59086\,
            PADOUT => \N__59085\,
            PADIN => \N__59084\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_STAT_COMM_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59077\,
            DIN => \N__59076\,
            DOUT => \N__59075\,
            PACKAGEPIN => \STAT_COMM_wire\
        );

    \ipInertedIOPad_STAT_COMM_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59077\,
            PADOUT => \N__59076\,
            PADIN => \N__59075\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19191\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SYSCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59068\,
            DIN => \N__59067\,
            DOUT => \N__59066\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ipInertedIOPad_ICE_SYSCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59068\,
            PADOUT => \N__59067\,
            PADIN => \N__59066\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SYSCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_161_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59059\,
            DIN => \N__59058\,
            DOUT => \N__59057\,
            PACKAGEPIN => \ICE_IOR_161_wire\
        );

    \ipInertedIOPad_ICE_IOR_161_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59059\,
            PADOUT => \N__59058\,
            PADIN => \N__59057\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_95_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59050\,
            DIN => \N__59049\,
            DOUT => \N__59048\,
            PACKAGEPIN => \ICE_IOB_95_wire\
        );

    \ipInertedIOPad_ICE_IOB_95_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59050\,
            PADOUT => \N__59049\,
            PADIN => \N__59048\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_82_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59041\,
            DIN => \N__59040\,
            DOUT => \N__59039\,
            PACKAGEPIN => \ICE_IOB_82_wire\
        );

    \ipInertedIOPad_ICE_IOB_82_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59041\,
            PADOUT => \N__59040\,
            PADIN => \N__59039\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_104_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59032\,
            DIN => \N__59031\,
            DOUT => \N__59030\,
            PACKAGEPIN => \ICE_IOB_104_wire\
        );

    \ipInertedIOPad_ICE_IOB_104_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59032\,
            PADOUT => \N__59031\,
            PADIN => \N__59030\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59023\,
            DIN => \N__59022\,
            DOUT => \N__59021\,
            PACKAGEPIN => \IAC_CLK_wire\
        );

    \ipInertedIOPad_IAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59023\,
            PADOUT => \N__59022\,
            PADIN => \N__59021\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22994\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59014\,
            DIN => \N__59013\,
            DOUT => \N__59012\,
            PACKAGEPIN => \DDS_CS_wire\
        );

    \ipInertedIOPad_DDS_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59014\,
            PADOUT => \N__59013\,
            PADIN => \N__59012\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36741\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59005\,
            DIN => \N__59004\,
            DOUT => \N__59003\,
            PACKAGEPIN => \SELIRNG0_wire\
        );

    \ipInertedIOPad_SELIRNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59005\,
            PADOUT => \N__59004\,
            PADIN => \N__59003\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31782\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58996\,
            DIN => \N__58995\,
            DOUT => \N__58994\,
            PACKAGEPIN => \RTD_SDI_wire\
        );

    \ipInertedIOPad_RTD_SDI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58996\,
            PADOUT => \N__58995\,
            PADIN => \N__58994\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19254\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_221_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58987\,
            DIN => \N__58986\,
            DOUT => \N__58985\,
            PACKAGEPIN => \ICE_IOT_221_wire\
        );

    \ipInertedIOPad_ICE_IOT_221_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58987\,
            PADOUT => \N__58986\,
            PADIN => \N__58985\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_197_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58978\,
            DIN => \N__58977\,
            DOUT => \N__58976\,
            PACKAGEPIN => \ICE_IOT_197_wire\
        );

    \ipInertedIOPad_ICE_IOT_197_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58978\,
            PADOUT => \N__58977\,
            PADIN => \N__58976\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58969\,
            DIN => \N__58968\,
            DOUT => \N__58967\,
            PACKAGEPIN => \DDS_MCLK_wire\
        );

    \ipInertedIOPad_DDS_MCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58969\,
            PADOUT => \N__58968\,
            PADIN => \N__58967\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__38649\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58960\,
            DIN => \N__58959\,
            DOUT => \N__58958\,
            PACKAGEPIN => \RTD_SCLK_wire\
        );

    \ipInertedIOPad_RTD_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58960\,
            PADOUT => \N__58959\,
            PADIN => \N__58958\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19224\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58951\,
            DIN => \N__58950\,
            DOUT => \N__58949\,
            PACKAGEPIN => \RTD_CS_wire\
        );

    \ipInertedIOPad_RTD_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58951\,
            PADOUT => \N__58950\,
            PADIN => \N__58949\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19581\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_137_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58942\,
            DIN => \N__58941\,
            DOUT => \N__58940\,
            PACKAGEPIN => \ICE_IOR_137_wire\
        );

    \ipInertedIOPad_ICE_IOR_137_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58942\,
            PADOUT => \N__58941\,
            PADIN => \N__58940\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58933\,
            DIN => \N__58932\,
            DOUT => \N__58931\,
            PACKAGEPIN => \IAC_OSR1_wire\
        );

    \ipInertedIOPad_IAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58933\,
            PADOUT => \N__58932\,
            PADIN => \N__58931\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__39807\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58924\,
            DIN => \N__58923\,
            DOUT => \N__58922\,
            PACKAGEPIN => \VAC_FLT0_wire\
        );

    \ipInertedIOPad_VAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58924\,
            PADOUT => \N__58923\,
            PADIN => \N__58922\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31902\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_144_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58915\,
            DIN => \N__58914\,
            DOUT => \N__58913\,
            PACKAGEPIN => \ICE_IOR_144_wire\
        );

    \ipInertedIOPad_ICE_IOR_144_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58915\,
            PADOUT => \N__58914\,
            PADIN => \N__58913\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_128_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58906\,
            DIN => \N__58905\,
            DOUT => \N__58904\,
            PACKAGEPIN => \ICE_IOR_128_wire\
        );

    \ipInertedIOPad_ICE_IOR_128_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58906\,
            PADOUT => \N__58905\,
            PADIN => \N__58904\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58897\,
            DIN => \N__58896\,
            DOUT => \N__58895\,
            PACKAGEPIN => \ICE_GPMO_1_wire\
        );

    \ipInertedIOPad_ICE_GPMO_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58897\,
            PADOUT => \N__58896\,
            PADIN => \N__58895\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58888\,
            DIN => \N__58887\,
            DOUT => \N__58886\,
            PACKAGEPIN => \IAC_SCLK_wire\
        );

    \ipInertedIOPad_IAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58888\,
            PADOUT => \N__58887\,
            PADIN => \N__58886\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23322\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_EIS_SYNCCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58879\,
            DIN => \N__58878\,
            DOUT => \N__58877\,
            PACKAGEPIN => \EIS_SYNCCLK_wire\
        );

    \ipInertedIOPad_EIS_SYNCCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58879\,
            PADOUT => \N__58878\,
            PADIN => \N__58877\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \EIS_SYNCCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_139_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58870\,
            DIN => \N__58869\,
            DOUT => \N__58868\,
            PACKAGEPIN => \ICE_IOR_139_wire\
        );

    \ipInertedIOPad_ICE_IOR_139_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58870\,
            PADOUT => \N__58869\,
            PADIN => \N__58868\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58861\,
            DIN => \N__58860\,
            DOUT => \N__58859\,
            PACKAGEPIN => \ICE_IOL_4A_wire\
        );

    \ipInertedIOPad_ICE_IOL_4A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58861\,
            PADOUT => \N__58860\,
            PADIN => \N__58859\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58852\,
            DIN => \N__58851\,
            DOUT => \N__58850\,
            PACKAGEPIN => \VAC_SCLK_wire\
        );

    \ipInertedIOPad_VAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58852\,
            PADOUT => \N__58851\,
            PADIN => \N__58850\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21957\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_THERMOSTAT_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58843\,
            DIN => \N__58842\,
            DOUT => \N__58841\,
            PACKAGEPIN => \THERMOSTAT_wire\
        );

    \ipInertedIOPad_THERMOSTAT_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58843\,
            PADOUT => \N__58842\,
            PADIN => \N__58841\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \THERMOSTAT\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_164_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58834\,
            DIN => \N__58833\,
            DOUT => \N__58832\,
            PACKAGEPIN => \ICE_IOR_164_wire\
        );

    \ipInertedIOPad_ICE_IOR_164_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58834\,
            PADOUT => \N__58833\,
            PADIN => \N__58832\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_103_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58825\,
            DIN => \N__58824\,
            DOUT => \N__58823\,
            PACKAGEPIN => \ICE_IOB_103_wire\
        );

    \ipInertedIOPad_ICE_IOB_103_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58825\,
            PADOUT => \N__58824\,
            PADIN => \N__58823\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AMPV_POW_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58816\,
            DIN => \N__58815\,
            DOUT => \N__58814\,
            PACKAGEPIN => \AMPV_POW_wire\
        );

    \ipInertedIOPad_AMPV_POW_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58816\,
            PADOUT => \N__58815\,
            PADIN => \N__58814\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23058\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SDO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58807\,
            DIN => \N__58806\,
            DOUT => \N__58805\,
            PACKAGEPIN => \VDC_SDO_wire\
        );

    \ipInertedIOPad_VDC_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58807\,
            PADOUT => \N__58806\,
            PADIN => \N__58805\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VDC_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_174_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58798\,
            DIN => \N__58797\,
            DOUT => \N__58796\,
            PACKAGEPIN => \ICE_IOT_174_wire\
        );

    \ipInertedIOPad_ICE_IOT_174_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58798\,
            PADOUT => \N__58797\,
            PADIN => \N__58796\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_140_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58789\,
            DIN => \N__58788\,
            DOUT => \N__58787\,
            PACKAGEPIN => \ICE_IOR_140_wire\
        );

    \ipInertedIOPad_ICE_IOR_140_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58789\,
            PADOUT => \N__58788\,
            PADIN => \N__58787\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_96_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58780\,
            DIN => \N__58779\,
            DOUT => \N__58778\,
            PACKAGEPIN => \ICE_IOB_96_wire\
        );

    \ipInertedIOPad_ICE_IOB_96_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58780\,
            PADOUT => \N__58779\,
            PADIN => \N__58778\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CONT_SD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58771\,
            DIN => \N__58770\,
            DOUT => \N__58769\,
            PACKAGEPIN => \CONT_SD_wire\
        );

    \ipInertedIOPad_CONT_SD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58771\,
            PADOUT => \N__58770\,
            PADIN => \N__58769\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44592\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AC_ADC_SYNC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58762\,
            DIN => \N__58761\,
            DOUT => \N__58760\,
            PACKAGEPIN => \AC_ADC_SYNC_wire\
        );

    \ipInertedIOPad_AC_ADC_SYNC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58762\,
            PADOUT => \N__58761\,
            PADIN => \N__58760\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21282\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58753\,
            DIN => \N__58752\,
            DOUT => \N__58751\,
            PACKAGEPIN => \SELIRNG1_wire\
        );

    \ipInertedIOPad_SELIRNG1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58753\,
            PADOUT => \N__58752\,
            PADIN => \N__58751\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__41964\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58744\,
            DIN => \N__58743\,
            DOUT => \N__58742\,
            PACKAGEPIN => \ICE_IOL_12B_wire\
        );

    \ipInertedIOPad_ICE_IOL_12B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58744\,
            PADOUT => \N__58743\,
            PADIN => \N__58742\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_160_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58735\,
            DIN => \N__58734\,
            DOUT => \N__58733\,
            PACKAGEPIN => \ICE_IOR_160_wire\
        );

    \ipInertedIOPad_ICE_IOR_160_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58735\,
            PADOUT => \N__58734\,
            PADIN => \N__58733\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_136_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58726\,
            DIN => \N__58725\,
            DOUT => \N__58724\,
            PACKAGEPIN => \ICE_IOR_136_wire\
        );

    \ipInertedIOPad_ICE_IOR_136_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58726\,
            PADOUT => \N__58725\,
            PADIN => \N__58724\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58717\,
            DIN => \N__58716\,
            DOUT => \N__58715\,
            PACKAGEPIN => \DDS_MCLK1_wire\
        );

    \ipInertedIOPad_DDS_MCLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58717\,
            PADOUT => \N__58716\,
            PADIN => \N__58715\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19596\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_198_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58708\,
            DIN => \N__58707\,
            DOUT => \N__58706\,
            PACKAGEPIN => \ICE_IOT_198_wire\
        );

    \ipInertedIOPad_ICE_IOT_198_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58708\,
            PADOUT => \N__58707\,
            PADIN => \N__58706\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_173_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58699\,
            DIN => \N__58698\,
            DOUT => \N__58697\,
            PACKAGEPIN => \ICE_IOT_173_wire\
        );

    \ipInertedIOPad_ICE_IOT_173_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58699\,
            PADOUT => \N__58698\,
            PADIN => \N__58697\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58690\,
            DIN => \N__58689\,
            DOUT => \N__58688\,
            PACKAGEPIN => \IAC_DRDY_wire\
        );

    \ipInertedIOPad_IAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58690\,
            PADOUT => \N__58689\,
            PADIN => \N__58688\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_178_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58681\,
            DIN => \N__58680\,
            DOUT => \N__58679\,
            PACKAGEPIN => \ICE_IOT_178_wire\
        );

    \ipInertedIOPad_ICE_IOT_178_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58681\,
            PADOUT => \N__58680\,
            PADIN => \N__58679\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_138_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58672\,
            DIN => \N__58671\,
            DOUT => \N__58670\,
            PACKAGEPIN => \ICE_IOR_138_wire\
        );

    \ipInertedIOPad_ICE_IOR_138_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58672\,
            PADOUT => \N__58671\,
            PADIN => \N__58670\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_120_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58663\,
            DIN => \N__58662\,
            DOUT => \N__58661\,
            PACKAGEPIN => \ICE_IOR_120_wire\
        );

    \ipInertedIOPad_ICE_IOR_120_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58663\,
            PADOUT => \N__58662\,
            PADIN => \N__58661\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58654\,
            DIN => \N__58653\,
            DOUT => \N__58652\,
            PACKAGEPIN => \IAC_FLT0_wire\
        );

    \ipInertedIOPad_IAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58654\,
            PADOUT => \N__58653\,
            PADIN => \N__58652\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44685\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58645\,
            DIN => \N__58644\,
            DOUT => \N__58643\,
            PACKAGEPIN => \DDS_SCK1_wire\
        );

    \ipInertedIOPad_DDS_SCK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58645\,
            PADOUT => \N__58644\,
            PADIN => \N__58643\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27132\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__14719\ : InMux
    port map (
            O => \N__58626\,
            I => \ADC_VDC.genclk.n19737\
        );

    \I__14718\ : CascadeMux
    port map (
            O => \N__58623\,
            I => \N__58617\
        );

    \I__14717\ : CascadeMux
    port map (
            O => \N__58622\,
            I => \N__58613\
        );

    \I__14716\ : CascadeMux
    port map (
            O => \N__58621\,
            I => \N__58609\
        );

    \I__14715\ : InMux
    port map (
            O => \N__58620\,
            I => \N__58592\
        );

    \I__14714\ : InMux
    port map (
            O => \N__58617\,
            I => \N__58592\
        );

    \I__14713\ : InMux
    port map (
            O => \N__58616\,
            I => \N__58592\
        );

    \I__14712\ : InMux
    port map (
            O => \N__58613\,
            I => \N__58592\
        );

    \I__14711\ : InMux
    port map (
            O => \N__58612\,
            I => \N__58592\
        );

    \I__14710\ : InMux
    port map (
            O => \N__58609\,
            I => \N__58592\
        );

    \I__14709\ : InMux
    port map (
            O => \N__58608\,
            I => \N__58592\
        );

    \I__14708\ : SRMux
    port map (
            O => \N__58607\,
            I => \N__58589\
        );

    \I__14707\ : LocalMux
    port map (
            O => \N__58592\,
            I => \N__58586\
        );

    \I__14706\ : LocalMux
    port map (
            O => \N__58589\,
            I => \N__58581\
        );

    \I__14705\ : Span4Mux_v
    port map (
            O => \N__58586\,
            I => \N__58570\
        );

    \I__14704\ : SRMux
    port map (
            O => \N__58585\,
            I => \N__58567\
        );

    \I__14703\ : SRMux
    port map (
            O => \N__58584\,
            I => \N__58561\
        );

    \I__14702\ : Span4Mux_h
    port map (
            O => \N__58581\,
            I => \N__58557\
        );

    \I__14701\ : CascadeMux
    port map (
            O => \N__58580\,
            I => \N__58554\
        );

    \I__14700\ : CascadeMux
    port map (
            O => \N__58579\,
            I => \N__58550\
        );

    \I__14699\ : CascadeMux
    port map (
            O => \N__58578\,
            I => \N__58546\
        );

    \I__14698\ : CascadeMux
    port map (
            O => \N__58577\,
            I => \N__58542\
        );

    \I__14697\ : CascadeMux
    port map (
            O => \N__58576\,
            I => \N__58538\
        );

    \I__14696\ : CascadeMux
    port map (
            O => \N__58575\,
            I => \N__58534\
        );

    \I__14695\ : CascadeMux
    port map (
            O => \N__58574\,
            I => \N__58530\
        );

    \I__14694\ : CascadeMux
    port map (
            O => \N__58573\,
            I => \N__58526\
        );

    \I__14693\ : Span4Mux_h
    port map (
            O => \N__58570\,
            I => \N__58519\
        );

    \I__14692\ : LocalMux
    port map (
            O => \N__58567\,
            I => \N__58516\
        );

    \I__14691\ : SRMux
    port map (
            O => \N__58566\,
            I => \N__58513\
        );

    \I__14690\ : SRMux
    port map (
            O => \N__58565\,
            I => \N__58510\
        );

    \I__14689\ : IoInMux
    port map (
            O => \N__58564\,
            I => \N__58504\
        );

    \I__14688\ : LocalMux
    port map (
            O => \N__58561\,
            I => \N__58497\
        );

    \I__14687\ : SRMux
    port map (
            O => \N__58560\,
            I => \N__58494\
        );

    \I__14686\ : Span4Mux_v
    port map (
            O => \N__58557\,
            I => \N__58491\
        );

    \I__14685\ : InMux
    port map (
            O => \N__58554\,
            I => \N__58476\
        );

    \I__14684\ : InMux
    port map (
            O => \N__58553\,
            I => \N__58476\
        );

    \I__14683\ : InMux
    port map (
            O => \N__58550\,
            I => \N__58476\
        );

    \I__14682\ : InMux
    port map (
            O => \N__58549\,
            I => \N__58476\
        );

    \I__14681\ : InMux
    port map (
            O => \N__58546\,
            I => \N__58476\
        );

    \I__14680\ : InMux
    port map (
            O => \N__58545\,
            I => \N__58476\
        );

    \I__14679\ : InMux
    port map (
            O => \N__58542\,
            I => \N__58476\
        );

    \I__14678\ : InMux
    port map (
            O => \N__58541\,
            I => \N__58459\
        );

    \I__14677\ : InMux
    port map (
            O => \N__58538\,
            I => \N__58459\
        );

    \I__14676\ : InMux
    port map (
            O => \N__58537\,
            I => \N__58459\
        );

    \I__14675\ : InMux
    port map (
            O => \N__58534\,
            I => \N__58459\
        );

    \I__14674\ : InMux
    port map (
            O => \N__58533\,
            I => \N__58459\
        );

    \I__14673\ : InMux
    port map (
            O => \N__58530\,
            I => \N__58459\
        );

    \I__14672\ : InMux
    port map (
            O => \N__58529\,
            I => \N__58459\
        );

    \I__14671\ : InMux
    port map (
            O => \N__58526\,
            I => \N__58459\
        );

    \I__14670\ : CascadeMux
    port map (
            O => \N__58525\,
            I => \N__58456\
        );

    \I__14669\ : CascadeMux
    port map (
            O => \N__58524\,
            I => \N__58452\
        );

    \I__14668\ : CascadeMux
    port map (
            O => \N__58523\,
            I => \N__58448\
        );

    \I__14667\ : CascadeMux
    port map (
            O => \N__58522\,
            I => \N__58444\
        );

    \I__14666\ : Span4Mux_h
    port map (
            O => \N__58519\,
            I => \N__58435\
        );

    \I__14665\ : Span4Mux_v
    port map (
            O => \N__58516\,
            I => \N__58435\
        );

    \I__14664\ : LocalMux
    port map (
            O => \N__58513\,
            I => \N__58435\
        );

    \I__14663\ : LocalMux
    port map (
            O => \N__58510\,
            I => \N__58435\
        );

    \I__14662\ : SRMux
    port map (
            O => \N__58509\,
            I => \N__58432\
        );

    \I__14661\ : SRMux
    port map (
            O => \N__58508\,
            I => \N__58429\
        );

    \I__14660\ : SRMux
    port map (
            O => \N__58507\,
            I => \N__58425\
        );

    \I__14659\ : LocalMux
    port map (
            O => \N__58504\,
            I => \N__58421\
        );

    \I__14658\ : CascadeMux
    port map (
            O => \N__58503\,
            I => \N__58417\
        );

    \I__14657\ : CascadeMux
    port map (
            O => \N__58502\,
            I => \N__58413\
        );

    \I__14656\ : CascadeMux
    port map (
            O => \N__58501\,
            I => \N__58409\
        );

    \I__14655\ : CascadeMux
    port map (
            O => \N__58500\,
            I => \N__58405\
        );

    \I__14654\ : Span4Mux_h
    port map (
            O => \N__58497\,
            I => \N__58400\
        );

    \I__14653\ : LocalMux
    port map (
            O => \N__58494\,
            I => \N__58400\
        );

    \I__14652\ : Span4Mux_v
    port map (
            O => \N__58491\,
            I => \N__58397\
        );

    \I__14651\ : LocalMux
    port map (
            O => \N__58476\,
            I => \N__58394\
        );

    \I__14650\ : LocalMux
    port map (
            O => \N__58459\,
            I => \N__58391\
        );

    \I__14649\ : InMux
    port map (
            O => \N__58456\,
            I => \N__58376\
        );

    \I__14648\ : InMux
    port map (
            O => \N__58455\,
            I => \N__58376\
        );

    \I__14647\ : InMux
    port map (
            O => \N__58452\,
            I => \N__58376\
        );

    \I__14646\ : InMux
    port map (
            O => \N__58451\,
            I => \N__58376\
        );

    \I__14645\ : InMux
    port map (
            O => \N__58448\,
            I => \N__58376\
        );

    \I__14644\ : InMux
    port map (
            O => \N__58447\,
            I => \N__58376\
        );

    \I__14643\ : InMux
    port map (
            O => \N__58444\,
            I => \N__58376\
        );

    \I__14642\ : Span4Mux_v
    port map (
            O => \N__58435\,
            I => \N__58369\
        );

    \I__14641\ : LocalMux
    port map (
            O => \N__58432\,
            I => \N__58369\
        );

    \I__14640\ : LocalMux
    port map (
            O => \N__58429\,
            I => \N__58369\
        );

    \I__14639\ : SRMux
    port map (
            O => \N__58428\,
            I => \N__58366\
        );

    \I__14638\ : LocalMux
    port map (
            O => \N__58425\,
            I => \N__58363\
        );

    \I__14637\ : SRMux
    port map (
            O => \N__58424\,
            I => \N__58360\
        );

    \I__14636\ : IoSpan4Mux
    port map (
            O => \N__58421\,
            I => \N__58356\
        );

    \I__14635\ : InMux
    port map (
            O => \N__58420\,
            I => \N__58339\
        );

    \I__14634\ : InMux
    port map (
            O => \N__58417\,
            I => \N__58339\
        );

    \I__14633\ : InMux
    port map (
            O => \N__58416\,
            I => \N__58339\
        );

    \I__14632\ : InMux
    port map (
            O => \N__58413\,
            I => \N__58339\
        );

    \I__14631\ : InMux
    port map (
            O => \N__58412\,
            I => \N__58339\
        );

    \I__14630\ : InMux
    port map (
            O => \N__58409\,
            I => \N__58339\
        );

    \I__14629\ : InMux
    port map (
            O => \N__58408\,
            I => \N__58339\
        );

    \I__14628\ : InMux
    port map (
            O => \N__58405\,
            I => \N__58339\
        );

    \I__14627\ : Span4Mux_v
    port map (
            O => \N__58400\,
            I => \N__58336\
        );

    \I__14626\ : Span4Mux_v
    port map (
            O => \N__58397\,
            I => \N__58326\
        );

    \I__14625\ : Span4Mux_h
    port map (
            O => \N__58394\,
            I => \N__58326\
        );

    \I__14624\ : Span4Mux_v
    port map (
            O => \N__58391\,
            I => \N__58326\
        );

    \I__14623\ : LocalMux
    port map (
            O => \N__58376\,
            I => \N__58326\
        );

    \I__14622\ : Span4Mux_v
    port map (
            O => \N__58369\,
            I => \N__58317\
        );

    \I__14621\ : LocalMux
    port map (
            O => \N__58366\,
            I => \N__58317\
        );

    \I__14620\ : Span4Mux_v
    port map (
            O => \N__58363\,
            I => \N__58317\
        );

    \I__14619\ : LocalMux
    port map (
            O => \N__58360\,
            I => \N__58317\
        );

    \I__14618\ : SRMux
    port map (
            O => \N__58359\,
            I => \N__58314\
        );

    \I__14617\ : Span4Mux_s0_v
    port map (
            O => \N__58356\,
            I => \N__58311\
        );

    \I__14616\ : LocalMux
    port map (
            O => \N__58339\,
            I => \N__58308\
        );

    \I__14615\ : Sp12to4
    port map (
            O => \N__58336\,
            I => \N__58305\
        );

    \I__14614\ : InMux
    port map (
            O => \N__58335\,
            I => \N__58302\
        );

    \I__14613\ : Span4Mux_v
    port map (
            O => \N__58326\,
            I => \N__58299\
        );

    \I__14612\ : Span4Mux_v
    port map (
            O => \N__58317\,
            I => \N__58294\
        );

    \I__14611\ : LocalMux
    port map (
            O => \N__58314\,
            I => \N__58294\
        );

    \I__14610\ : Sp12to4
    port map (
            O => \N__58311\,
            I => \N__58288\
        );

    \I__14609\ : Span12Mux_s10_h
    port map (
            O => \N__58308\,
            I => \N__58288\
        );

    \I__14608\ : Span12Mux_h
    port map (
            O => \N__58305\,
            I => \N__58283\
        );

    \I__14607\ : LocalMux
    port map (
            O => \N__58302\,
            I => \N__58283\
        );

    \I__14606\ : Sp12to4
    port map (
            O => \N__58299\,
            I => \N__58278\
        );

    \I__14605\ : Sp12to4
    port map (
            O => \N__58294\,
            I => \N__58278\
        );

    \I__14604\ : InMux
    port map (
            O => \N__58293\,
            I => \N__58275\
        );

    \I__14603\ : Odrv12
    port map (
            O => \N__58288\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14602\ : Odrv12
    port map (
            O => \N__58283\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14601\ : Odrv12
    port map (
            O => \N__58278\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14600\ : LocalMux
    port map (
            O => \N__58275\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14599\ : InMux
    port map (
            O => \N__58266\,
            I => \ADC_VDC.genclk.n19738\
        );

    \I__14598\ : SRMux
    port map (
            O => \N__58263\,
            I => \N__58260\
        );

    \I__14597\ : LocalMux
    port map (
            O => \N__58260\,
            I => \N__58255\
        );

    \I__14596\ : SRMux
    port map (
            O => \N__58259\,
            I => \N__58252\
        );

    \I__14595\ : SRMux
    port map (
            O => \N__58258\,
            I => \N__58249\
        );

    \I__14594\ : Span4Mux_v
    port map (
            O => \N__58255\,
            I => \N__58244\
        );

    \I__14593\ : LocalMux
    port map (
            O => \N__58252\,
            I => \N__58244\
        );

    \I__14592\ : LocalMux
    port map (
            O => \N__58249\,
            I => \N__58240\
        );

    \I__14591\ : Span4Mux_h
    port map (
            O => \N__58244\,
            I => \N__58237\
        );

    \I__14590\ : SRMux
    port map (
            O => \N__58243\,
            I => \N__58234\
        );

    \I__14589\ : Span4Mux_v
    port map (
            O => \N__58240\,
            I => \N__58231\
        );

    \I__14588\ : Sp12to4
    port map (
            O => \N__58237\,
            I => \N__58226\
        );

    \I__14587\ : LocalMux
    port map (
            O => \N__58234\,
            I => \N__58226\
        );

    \I__14586\ : Odrv4
    port map (
            O => \N__58231\,
            I => \ADC_VDC.genclk.n15051\
        );

    \I__14585\ : Odrv12
    port map (
            O => \N__58226\,
            I => \ADC_VDC.genclk.n15051\
        );

    \I__14584\ : CascadeMux
    port map (
            O => \N__58221\,
            I => \N__58218\
        );

    \I__14583\ : InMux
    port map (
            O => \N__58218\,
            I => \N__58214\
        );

    \I__14582\ : InMux
    port map (
            O => \N__58217\,
            I => \N__58211\
        );

    \I__14581\ : LocalMux
    port map (
            O => \N__58214\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__14580\ : LocalMux
    port map (
            O => \N__58211\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__14579\ : InMux
    port map (
            O => \N__58206\,
            I => \N__58202\
        );

    \I__14578\ : InMux
    port map (
            O => \N__58205\,
            I => \N__58199\
        );

    \I__14577\ : LocalMux
    port map (
            O => \N__58202\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__14576\ : LocalMux
    port map (
            O => \N__58199\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__14575\ : CascadeMux
    port map (
            O => \N__58194\,
            I => \N__58190\
        );

    \I__14574\ : CascadeMux
    port map (
            O => \N__58193\,
            I => \N__58187\
        );

    \I__14573\ : InMux
    port map (
            O => \N__58190\,
            I => \N__58184\
        );

    \I__14572\ : InMux
    port map (
            O => \N__58187\,
            I => \N__58181\
        );

    \I__14571\ : LocalMux
    port map (
            O => \N__58184\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__14570\ : LocalMux
    port map (
            O => \N__58181\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__14569\ : InMux
    port map (
            O => \N__58176\,
            I => \N__58172\
        );

    \I__14568\ : InMux
    port map (
            O => \N__58175\,
            I => \N__58169\
        );

    \I__14567\ : LocalMux
    port map (
            O => \N__58172\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__14566\ : LocalMux
    port map (
            O => \N__58169\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__14565\ : CascadeMux
    port map (
            O => \N__58164\,
            I => \ADC_VDC.genclk.n21449_cascade_\
        );

    \I__14564\ : CascadeMux
    port map (
            O => \N__58161\,
            I => \N__58157\
        );

    \I__14563\ : CascadeMux
    port map (
            O => \N__58160\,
            I => \N__58154\
        );

    \I__14562\ : InMux
    port map (
            O => \N__58157\,
            I => \N__58151\
        );

    \I__14561\ : InMux
    port map (
            O => \N__58154\,
            I => \N__58148\
        );

    \I__14560\ : LocalMux
    port map (
            O => \N__58151\,
            I => \N__58145\
        );

    \I__14559\ : LocalMux
    port map (
            O => \N__58148\,
            I => \N__58142\
        );

    \I__14558\ : Span4Mux_h
    port map (
            O => \N__58145\,
            I => \N__58139\
        );

    \I__14557\ : Span4Mux_h
    port map (
            O => \N__58142\,
            I => \N__58136\
        );

    \I__14556\ : Odrv4
    port map (
            O => \N__58139\,
            I => \ADC_VDC.genclk.n21443\
        );

    \I__14555\ : Odrv4
    port map (
            O => \N__58136\,
            I => \ADC_VDC.genclk.n21443\
        );

    \I__14554\ : InMux
    port map (
            O => \N__58131\,
            I => \N__58127\
        );

    \I__14553\ : InMux
    port map (
            O => \N__58130\,
            I => \N__58124\
        );

    \I__14552\ : LocalMux
    port map (
            O => \N__58127\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__14551\ : LocalMux
    port map (
            O => \N__58124\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__14550\ : CascadeMux
    port map (
            O => \N__58119\,
            I => \N__58116\
        );

    \I__14549\ : InMux
    port map (
            O => \N__58116\,
            I => \N__58112\
        );

    \I__14548\ : InMux
    port map (
            O => \N__58115\,
            I => \N__58109\
        );

    \I__14547\ : LocalMux
    port map (
            O => \N__58112\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__14546\ : LocalMux
    port map (
            O => \N__58109\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__14545\ : CascadeMux
    port map (
            O => \N__58104\,
            I => \N__58100\
        );

    \I__14544\ : InMux
    port map (
            O => \N__58103\,
            I => \N__58097\
        );

    \I__14543\ : InMux
    port map (
            O => \N__58100\,
            I => \N__58094\
        );

    \I__14542\ : LocalMux
    port map (
            O => \N__58097\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__14541\ : LocalMux
    port map (
            O => \N__58094\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__14540\ : InMux
    port map (
            O => \N__58089\,
            I => \N__58085\
        );

    \I__14539\ : InMux
    port map (
            O => \N__58088\,
            I => \N__58082\
        );

    \I__14538\ : LocalMux
    port map (
            O => \N__58085\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__14537\ : LocalMux
    port map (
            O => \N__58082\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__14536\ : InMux
    port map (
            O => \N__58077\,
            I => \N__58074\
        );

    \I__14535\ : LocalMux
    port map (
            O => \N__58074\,
            I => \ADC_VDC.genclk.n27_adj_1396\
        );

    \I__14534\ : InMux
    port map (
            O => \N__58071\,
            I => \N__58067\
        );

    \I__14533\ : InMux
    port map (
            O => \N__58070\,
            I => \N__58064\
        );

    \I__14532\ : LocalMux
    port map (
            O => \N__58067\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__14531\ : LocalMux
    port map (
            O => \N__58064\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__14530\ : CascadeMux
    port map (
            O => \N__58059\,
            I => \N__58056\
        );

    \I__14529\ : InMux
    port map (
            O => \N__58056\,
            I => \N__58052\
        );

    \I__14528\ : InMux
    port map (
            O => \N__58055\,
            I => \N__58049\
        );

    \I__14527\ : LocalMux
    port map (
            O => \N__58052\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__14526\ : LocalMux
    port map (
            O => \N__58049\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__14525\ : CascadeMux
    port map (
            O => \N__58044\,
            I => \N__58040\
        );

    \I__14524\ : InMux
    port map (
            O => \N__58043\,
            I => \N__58037\
        );

    \I__14523\ : InMux
    port map (
            O => \N__58040\,
            I => \N__58034\
        );

    \I__14522\ : LocalMux
    port map (
            O => \N__58037\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__14521\ : LocalMux
    port map (
            O => \N__58034\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__14520\ : InMux
    port map (
            O => \N__58029\,
            I => \N__58025\
        );

    \I__14519\ : InMux
    port map (
            O => \N__58028\,
            I => \N__58022\
        );

    \I__14518\ : LocalMux
    port map (
            O => \N__58025\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__14517\ : LocalMux
    port map (
            O => \N__58022\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__14516\ : InMux
    port map (
            O => \N__58017\,
            I => \N__58014\
        );

    \I__14515\ : LocalMux
    port map (
            O => \N__58014\,
            I => \ADC_VDC.genclk.n26_adj_1395\
        );

    \I__14514\ : InMux
    port map (
            O => \N__58011\,
            I => \N__58007\
        );

    \I__14513\ : InMux
    port map (
            O => \N__58010\,
            I => \N__57999\
        );

    \I__14512\ : LocalMux
    port map (
            O => \N__58007\,
            I => \N__57996\
        );

    \I__14511\ : InMux
    port map (
            O => \N__58006\,
            I => \N__57993\
        );

    \I__14510\ : InMux
    port map (
            O => \N__58005\,
            I => \N__57986\
        );

    \I__14509\ : InMux
    port map (
            O => \N__58004\,
            I => \N__57986\
        );

    \I__14508\ : InMux
    port map (
            O => \N__58003\,
            I => \N__57986\
        );

    \I__14507\ : InMux
    port map (
            O => \N__58002\,
            I => \N__57983\
        );

    \I__14506\ : LocalMux
    port map (
            O => \N__57999\,
            I => \N__57978\
        );

    \I__14505\ : Span4Mux_h
    port map (
            O => \N__57996\,
            I => \N__57978\
        );

    \I__14504\ : LocalMux
    port map (
            O => \N__57993\,
            I => \N__57975\
        );

    \I__14503\ : LocalMux
    port map (
            O => \N__57986\,
            I => \N__57972\
        );

    \I__14502\ : LocalMux
    port map (
            O => \N__57983\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__14501\ : Odrv4
    port map (
            O => \N__57978\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__14500\ : Odrv4
    port map (
            O => \N__57975\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__14499\ : Odrv4
    port map (
            O => \N__57972\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__14498\ : CEMux
    port map (
            O => \N__57963\,
            I => \N__57960\
        );

    \I__14497\ : LocalMux
    port map (
            O => \N__57960\,
            I => \N__57956\
        );

    \I__14496\ : CEMux
    port map (
            O => \N__57959\,
            I => \N__57953\
        );

    \I__14495\ : Span4Mux_v
    port map (
            O => \N__57956\,
            I => \N__57950\
        );

    \I__14494\ : LocalMux
    port map (
            O => \N__57953\,
            I => \N__57947\
        );

    \I__14493\ : Span4Mux_h
    port map (
            O => \N__57950\,
            I => \N__57944\
        );

    \I__14492\ : Span4Mux_h
    port map (
            O => \N__57947\,
            I => \N__57941\
        );

    \I__14491\ : Odrv4
    port map (
            O => \N__57944\,
            I => \ADC_VDC.genclk.div_state_1__N_1274\
        );

    \I__14490\ : Odrv4
    port map (
            O => \N__57941\,
            I => \ADC_VDC.genclk.div_state_1__N_1274\
        );

    \I__14489\ : InMux
    port map (
            O => \N__57936\,
            I => \N__57932\
        );

    \I__14488\ : InMux
    port map (
            O => \N__57935\,
            I => \N__57929\
        );

    \I__14487\ : LocalMux
    port map (
            O => \N__57932\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__14486\ : LocalMux
    port map (
            O => \N__57929\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__14485\ : CascadeMux
    port map (
            O => \N__57924\,
            I => \N__57921\
        );

    \I__14484\ : InMux
    port map (
            O => \N__57921\,
            I => \N__57917\
        );

    \I__14483\ : InMux
    port map (
            O => \N__57920\,
            I => \N__57914\
        );

    \I__14482\ : LocalMux
    port map (
            O => \N__57917\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__14481\ : LocalMux
    port map (
            O => \N__57914\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__14480\ : CascadeMux
    port map (
            O => \N__57909\,
            I => \N__57905\
        );

    \I__14479\ : InMux
    port map (
            O => \N__57908\,
            I => \N__57902\
        );

    \I__14478\ : InMux
    port map (
            O => \N__57905\,
            I => \N__57899\
        );

    \I__14477\ : LocalMux
    port map (
            O => \N__57902\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__14476\ : LocalMux
    port map (
            O => \N__57899\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__14475\ : CascadeMux
    port map (
            O => \N__57894\,
            I => \N__57891\
        );

    \I__14474\ : InMux
    port map (
            O => \N__57891\,
            I => \N__57887\
        );

    \I__14473\ : InMux
    port map (
            O => \N__57890\,
            I => \N__57884\
        );

    \I__14472\ : LocalMux
    port map (
            O => \N__57887\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__14471\ : LocalMux
    port map (
            O => \N__57884\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__14470\ : InMux
    port map (
            O => \N__57879\,
            I => \N__57876\
        );

    \I__14469\ : LocalMux
    port map (
            O => \N__57876\,
            I => \N__57873\
        );

    \I__14468\ : Odrv4
    port map (
            O => \N__57873\,
            I => \ADC_VDC.genclk.n28\
        );

    \I__14467\ : InMux
    port map (
            O => \N__57870\,
            I => \ADC_VDC.genclk.n19728\
        );

    \I__14466\ : InMux
    port map (
            O => \N__57867\,
            I => \ADC_VDC.genclk.n19729\
        );

    \I__14465\ : InMux
    port map (
            O => \N__57864\,
            I => \ADC_VDC.genclk.n19730\
        );

    \I__14464\ : InMux
    port map (
            O => \N__57861\,
            I => \bfn_22_8_0_\
        );

    \I__14463\ : InMux
    port map (
            O => \N__57858\,
            I => \ADC_VDC.genclk.n19732\
        );

    \I__14462\ : InMux
    port map (
            O => \N__57855\,
            I => \ADC_VDC.genclk.n19733\
        );

    \I__14461\ : InMux
    port map (
            O => \N__57852\,
            I => \ADC_VDC.genclk.n19734\
        );

    \I__14460\ : InMux
    port map (
            O => \N__57849\,
            I => \ADC_VDC.genclk.n19735\
        );

    \I__14459\ : InMux
    port map (
            O => \N__57846\,
            I => \ADC_VDC.genclk.n19736\
        );

    \I__14458\ : InMux
    port map (
            O => \N__57843\,
            I => \N__57840\
        );

    \I__14457\ : LocalMux
    port map (
            O => \N__57840\,
            I => buf_data_iac_13
        );

    \I__14456\ : InMux
    port map (
            O => \N__57837\,
            I => \N__57834\
        );

    \I__14455\ : LocalMux
    port map (
            O => \N__57834\,
            I => n21350
        );

    \I__14454\ : InMux
    port map (
            O => \N__57831\,
            I => \N__57828\
        );

    \I__14453\ : LocalMux
    port map (
            O => \N__57828\,
            I => buf_data_iac_9
        );

    \I__14452\ : CascadeMux
    port map (
            O => \N__57825\,
            I => \N__57809\
        );

    \I__14451\ : InMux
    port map (
            O => \N__57824\,
            I => \N__57797\
        );

    \I__14450\ : InMux
    port map (
            O => \N__57823\,
            I => \N__57789\
        );

    \I__14449\ : InMux
    port map (
            O => \N__57822\,
            I => \N__57773\
        );

    \I__14448\ : InMux
    port map (
            O => \N__57821\,
            I => \N__57770\
        );

    \I__14447\ : InMux
    port map (
            O => \N__57820\,
            I => \N__57767\
        );

    \I__14446\ : CascadeMux
    port map (
            O => \N__57819\,
            I => \N__57764\
        );

    \I__14445\ : InMux
    port map (
            O => \N__57818\,
            I => \N__57760\
        );

    \I__14444\ : InMux
    port map (
            O => \N__57817\,
            I => \N__57751\
        );

    \I__14443\ : InMux
    port map (
            O => \N__57816\,
            I => \N__57744\
        );

    \I__14442\ : InMux
    port map (
            O => \N__57815\,
            I => \N__57741\
        );

    \I__14441\ : InMux
    port map (
            O => \N__57814\,
            I => \N__57729\
        );

    \I__14440\ : InMux
    port map (
            O => \N__57813\,
            I => \N__57729\
        );

    \I__14439\ : InMux
    port map (
            O => \N__57812\,
            I => \N__57729\
        );

    \I__14438\ : InMux
    port map (
            O => \N__57809\,
            I => \N__57724\
        );

    \I__14437\ : InMux
    port map (
            O => \N__57808\,
            I => \N__57724\
        );

    \I__14436\ : InMux
    port map (
            O => \N__57807\,
            I => \N__57717\
        );

    \I__14435\ : InMux
    port map (
            O => \N__57806\,
            I => \N__57717\
        );

    \I__14434\ : InMux
    port map (
            O => \N__57805\,
            I => \N__57717\
        );

    \I__14433\ : InMux
    port map (
            O => \N__57804\,
            I => \N__57714\
        );

    \I__14432\ : InMux
    port map (
            O => \N__57803\,
            I => \N__57705\
        );

    \I__14431\ : InMux
    port map (
            O => \N__57802\,
            I => \N__57705\
        );

    \I__14430\ : InMux
    port map (
            O => \N__57801\,
            I => \N__57705\
        );

    \I__14429\ : InMux
    port map (
            O => \N__57800\,
            I => \N__57705\
        );

    \I__14428\ : LocalMux
    port map (
            O => \N__57797\,
            I => \N__57702\
        );

    \I__14427\ : InMux
    port map (
            O => \N__57796\,
            I => \N__57695\
        );

    \I__14426\ : InMux
    port map (
            O => \N__57795\,
            I => \N__57690\
        );

    \I__14425\ : InMux
    port map (
            O => \N__57794\,
            I => \N__57690\
        );

    \I__14424\ : InMux
    port map (
            O => \N__57793\,
            I => \N__57685\
        );

    \I__14423\ : InMux
    port map (
            O => \N__57792\,
            I => \N__57685\
        );

    \I__14422\ : LocalMux
    port map (
            O => \N__57789\,
            I => \N__57682\
        );

    \I__14421\ : InMux
    port map (
            O => \N__57788\,
            I => \N__57675\
        );

    \I__14420\ : InMux
    port map (
            O => \N__57787\,
            I => \N__57675\
        );

    \I__14419\ : InMux
    port map (
            O => \N__57786\,
            I => \N__57675\
        );

    \I__14418\ : InMux
    port map (
            O => \N__57785\,
            I => \N__57672\
        );

    \I__14417\ : InMux
    port map (
            O => \N__57784\,
            I => \N__57669\
        );

    \I__14416\ : InMux
    port map (
            O => \N__57783\,
            I => \N__57662\
        );

    \I__14415\ : InMux
    port map (
            O => \N__57782\,
            I => \N__57658\
        );

    \I__14414\ : InMux
    port map (
            O => \N__57781\,
            I => \N__57655\
        );

    \I__14413\ : InMux
    port map (
            O => \N__57780\,
            I => \N__57648\
        );

    \I__14412\ : InMux
    port map (
            O => \N__57779\,
            I => \N__57643\
        );

    \I__14411\ : InMux
    port map (
            O => \N__57778\,
            I => \N__57643\
        );

    \I__14410\ : InMux
    port map (
            O => \N__57777\,
            I => \N__57638\
        );

    \I__14409\ : InMux
    port map (
            O => \N__57776\,
            I => \N__57635\
        );

    \I__14408\ : LocalMux
    port map (
            O => \N__57773\,
            I => \N__57632\
        );

    \I__14407\ : LocalMux
    port map (
            O => \N__57770\,
            I => \N__57627\
        );

    \I__14406\ : LocalMux
    port map (
            O => \N__57767\,
            I => \N__57627\
        );

    \I__14405\ : InMux
    port map (
            O => \N__57764\,
            I => \N__57619\
        );

    \I__14404\ : InMux
    port map (
            O => \N__57763\,
            I => \N__57619\
        );

    \I__14403\ : LocalMux
    port map (
            O => \N__57760\,
            I => \N__57611\
        );

    \I__14402\ : InMux
    port map (
            O => \N__57759\,
            I => \N__57608\
        );

    \I__14401\ : InMux
    port map (
            O => \N__57758\,
            I => \N__57605\
        );

    \I__14400\ : InMux
    port map (
            O => \N__57757\,
            I => \N__57600\
        );

    \I__14399\ : InMux
    port map (
            O => \N__57756\,
            I => \N__57597\
        );

    \I__14398\ : InMux
    port map (
            O => \N__57755\,
            I => \N__57594\
        );

    \I__14397\ : InMux
    port map (
            O => \N__57754\,
            I => \N__57585\
        );

    \I__14396\ : LocalMux
    port map (
            O => \N__57751\,
            I => \N__57582\
        );

    \I__14395\ : InMux
    port map (
            O => \N__57750\,
            I => \N__57579\
        );

    \I__14394\ : InMux
    port map (
            O => \N__57749\,
            I => \N__57576\
        );

    \I__14393\ : InMux
    port map (
            O => \N__57748\,
            I => \N__57573\
        );

    \I__14392\ : InMux
    port map (
            O => \N__57747\,
            I => \N__57569\
        );

    \I__14391\ : LocalMux
    port map (
            O => \N__57744\,
            I => \N__57564\
        );

    \I__14390\ : LocalMux
    port map (
            O => \N__57741\,
            I => \N__57564\
        );

    \I__14389\ : InMux
    port map (
            O => \N__57740\,
            I => \N__57561\
        );

    \I__14388\ : InMux
    port map (
            O => \N__57739\,
            I => \N__57558\
        );

    \I__14387\ : InMux
    port map (
            O => \N__57738\,
            I => \N__57555\
        );

    \I__14386\ : InMux
    port map (
            O => \N__57737\,
            I => \N__57550\
        );

    \I__14385\ : InMux
    port map (
            O => \N__57736\,
            I => \N__57547\
        );

    \I__14384\ : LocalMux
    port map (
            O => \N__57729\,
            I => \N__57544\
        );

    \I__14383\ : LocalMux
    port map (
            O => \N__57724\,
            I => \N__57539\
        );

    \I__14382\ : LocalMux
    port map (
            O => \N__57717\,
            I => \N__57539\
        );

    \I__14381\ : LocalMux
    port map (
            O => \N__57714\,
            I => \N__57532\
        );

    \I__14380\ : LocalMux
    port map (
            O => \N__57705\,
            I => \N__57532\
        );

    \I__14379\ : Span4Mux_h
    port map (
            O => \N__57702\,
            I => \N__57532\
        );

    \I__14378\ : InMux
    port map (
            O => \N__57701\,
            I => \N__57527\
        );

    \I__14377\ : InMux
    port map (
            O => \N__57700\,
            I => \N__57527\
        );

    \I__14376\ : InMux
    port map (
            O => \N__57699\,
            I => \N__57524\
        );

    \I__14375\ : InMux
    port map (
            O => \N__57698\,
            I => \N__57521\
        );

    \I__14374\ : LocalMux
    port map (
            O => \N__57695\,
            I => \N__57508\
        );

    \I__14373\ : LocalMux
    port map (
            O => \N__57690\,
            I => \N__57508\
        );

    \I__14372\ : LocalMux
    port map (
            O => \N__57685\,
            I => \N__57508\
        );

    \I__14371\ : Span4Mux_h
    port map (
            O => \N__57682\,
            I => \N__57508\
        );

    \I__14370\ : LocalMux
    port map (
            O => \N__57675\,
            I => \N__57508\
        );

    \I__14369\ : LocalMux
    port map (
            O => \N__57672\,
            I => \N__57508\
        );

    \I__14368\ : LocalMux
    port map (
            O => \N__57669\,
            I => \N__57505\
        );

    \I__14367\ : InMux
    port map (
            O => \N__57668\,
            I => \N__57500\
        );

    \I__14366\ : InMux
    port map (
            O => \N__57667\,
            I => \N__57500\
        );

    \I__14365\ : InMux
    port map (
            O => \N__57666\,
            I => \N__57493\
        );

    \I__14364\ : InMux
    port map (
            O => \N__57665\,
            I => \N__57493\
        );

    \I__14363\ : LocalMux
    port map (
            O => \N__57662\,
            I => \N__57490\
        );

    \I__14362\ : InMux
    port map (
            O => \N__57661\,
            I => \N__57487\
        );

    \I__14361\ : LocalMux
    port map (
            O => \N__57658\,
            I => \N__57484\
        );

    \I__14360\ : LocalMux
    port map (
            O => \N__57655\,
            I => \N__57481\
        );

    \I__14359\ : InMux
    port map (
            O => \N__57654\,
            I => \N__57478\
        );

    \I__14358\ : InMux
    port map (
            O => \N__57653\,
            I => \N__57467\
        );

    \I__14357\ : InMux
    port map (
            O => \N__57652\,
            I => \N__57467\
        );

    \I__14356\ : InMux
    port map (
            O => \N__57651\,
            I => \N__57467\
        );

    \I__14355\ : LocalMux
    port map (
            O => \N__57648\,
            I => \N__57462\
        );

    \I__14354\ : LocalMux
    port map (
            O => \N__57643\,
            I => \N__57462\
        );

    \I__14353\ : InMux
    port map (
            O => \N__57642\,
            I => \N__57459\
        );

    \I__14352\ : InMux
    port map (
            O => \N__57641\,
            I => \N__57456\
        );

    \I__14351\ : LocalMux
    port map (
            O => \N__57638\,
            I => \N__57451\
        );

    \I__14350\ : LocalMux
    port map (
            O => \N__57635\,
            I => \N__57451\
        );

    \I__14349\ : Span4Mux_v
    port map (
            O => \N__57632\,
            I => \N__57446\
        );

    \I__14348\ : Span4Mux_h
    port map (
            O => \N__57627\,
            I => \N__57446\
        );

    \I__14347\ : InMux
    port map (
            O => \N__57626\,
            I => \N__57443\
        );

    \I__14346\ : InMux
    port map (
            O => \N__57625\,
            I => \N__57440\
        );

    \I__14345\ : InMux
    port map (
            O => \N__57624\,
            I => \N__57437\
        );

    \I__14344\ : LocalMux
    port map (
            O => \N__57619\,
            I => \N__57434\
        );

    \I__14343\ : InMux
    port map (
            O => \N__57618\,
            I => \N__57423\
        );

    \I__14342\ : InMux
    port map (
            O => \N__57617\,
            I => \N__57423\
        );

    \I__14341\ : InMux
    port map (
            O => \N__57616\,
            I => \N__57423\
        );

    \I__14340\ : InMux
    port map (
            O => \N__57615\,
            I => \N__57423\
        );

    \I__14339\ : InMux
    port map (
            O => \N__57614\,
            I => \N__57423\
        );

    \I__14338\ : Span4Mux_h
    port map (
            O => \N__57611\,
            I => \N__57416\
        );

    \I__14337\ : LocalMux
    port map (
            O => \N__57608\,
            I => \N__57416\
        );

    \I__14336\ : LocalMux
    port map (
            O => \N__57605\,
            I => \N__57416\
        );

    \I__14335\ : InMux
    port map (
            O => \N__57604\,
            I => \N__57411\
        );

    \I__14334\ : InMux
    port map (
            O => \N__57603\,
            I => \N__57411\
        );

    \I__14333\ : LocalMux
    port map (
            O => \N__57600\,
            I => \N__57404\
        );

    \I__14332\ : LocalMux
    port map (
            O => \N__57597\,
            I => \N__57404\
        );

    \I__14331\ : LocalMux
    port map (
            O => \N__57594\,
            I => \N__57404\
        );

    \I__14330\ : InMux
    port map (
            O => \N__57593\,
            I => \N__57399\
        );

    \I__14329\ : InMux
    port map (
            O => \N__57592\,
            I => \N__57399\
        );

    \I__14328\ : InMux
    port map (
            O => \N__57591\,
            I => \N__57394\
        );

    \I__14327\ : InMux
    port map (
            O => \N__57590\,
            I => \N__57394\
        );

    \I__14326\ : InMux
    port map (
            O => \N__57589\,
            I => \N__57389\
        );

    \I__14325\ : InMux
    port map (
            O => \N__57588\,
            I => \N__57389\
        );

    \I__14324\ : LocalMux
    port map (
            O => \N__57585\,
            I => \N__57370\
        );

    \I__14323\ : Sp12to4
    port map (
            O => \N__57582\,
            I => \N__57370\
        );

    \I__14322\ : LocalMux
    port map (
            O => \N__57579\,
            I => \N__57370\
        );

    \I__14321\ : LocalMux
    port map (
            O => \N__57576\,
            I => \N__57370\
        );

    \I__14320\ : LocalMux
    port map (
            O => \N__57573\,
            I => \N__57370\
        );

    \I__14319\ : InMux
    port map (
            O => \N__57572\,
            I => \N__57367\
        );

    \I__14318\ : LocalMux
    port map (
            O => \N__57569\,
            I => \N__57362\
        );

    \I__14317\ : Sp12to4
    port map (
            O => \N__57564\,
            I => \N__57362\
        );

    \I__14316\ : LocalMux
    port map (
            O => \N__57561\,
            I => \N__57355\
        );

    \I__14315\ : LocalMux
    port map (
            O => \N__57558\,
            I => \N__57355\
        );

    \I__14314\ : LocalMux
    port map (
            O => \N__57555\,
            I => \N__57355\
        );

    \I__14313\ : InMux
    port map (
            O => \N__57554\,
            I => \N__57352\
        );

    \I__14312\ : InMux
    port map (
            O => \N__57553\,
            I => \N__57349\
        );

    \I__14311\ : LocalMux
    port map (
            O => \N__57550\,
            I => \N__57346\
        );

    \I__14310\ : LocalMux
    port map (
            O => \N__57547\,
            I => \N__57335\
        );

    \I__14309\ : Span4Mux_h
    port map (
            O => \N__57544\,
            I => \N__57335\
        );

    \I__14308\ : Span4Mux_h
    port map (
            O => \N__57539\,
            I => \N__57335\
        );

    \I__14307\ : Span4Mux_v
    port map (
            O => \N__57532\,
            I => \N__57335\
        );

    \I__14306\ : LocalMux
    port map (
            O => \N__57527\,
            I => \N__57335\
        );

    \I__14305\ : LocalMux
    port map (
            O => \N__57524\,
            I => \N__57330\
        );

    \I__14304\ : LocalMux
    port map (
            O => \N__57521\,
            I => \N__57330\
        );

    \I__14303\ : Span4Mux_v
    port map (
            O => \N__57508\,
            I => \N__57323\
        );

    \I__14302\ : Span4Mux_h
    port map (
            O => \N__57505\,
            I => \N__57323\
        );

    \I__14301\ : LocalMux
    port map (
            O => \N__57500\,
            I => \N__57323\
        );

    \I__14300\ : InMux
    port map (
            O => \N__57499\,
            I => \N__57320\
        );

    \I__14299\ : InMux
    port map (
            O => \N__57498\,
            I => \N__57317\
        );

    \I__14298\ : LocalMux
    port map (
            O => \N__57493\,
            I => \N__57312\
        );

    \I__14297\ : Span4Mux_v
    port map (
            O => \N__57490\,
            I => \N__57312\
        );

    \I__14296\ : LocalMux
    port map (
            O => \N__57487\,
            I => \N__57303\
        );

    \I__14295\ : Span4Mux_h
    port map (
            O => \N__57484\,
            I => \N__57303\
        );

    \I__14294\ : Span4Mux_h
    port map (
            O => \N__57481\,
            I => \N__57303\
        );

    \I__14293\ : LocalMux
    port map (
            O => \N__57478\,
            I => \N__57303\
        );

    \I__14292\ : InMux
    port map (
            O => \N__57477\,
            I => \N__57300\
        );

    \I__14291\ : InMux
    port map (
            O => \N__57476\,
            I => \N__57293\
        );

    \I__14290\ : InMux
    port map (
            O => \N__57475\,
            I => \N__57293\
        );

    \I__14289\ : InMux
    port map (
            O => \N__57474\,
            I => \N__57293\
        );

    \I__14288\ : LocalMux
    port map (
            O => \N__57467\,
            I => \N__57288\
        );

    \I__14287\ : Span4Mux_v
    port map (
            O => \N__57462\,
            I => \N__57288\
        );

    \I__14286\ : LocalMux
    port map (
            O => \N__57459\,
            I => \N__57281\
        );

    \I__14285\ : LocalMux
    port map (
            O => \N__57456\,
            I => \N__57281\
        );

    \I__14284\ : Span4Mux_v
    port map (
            O => \N__57451\,
            I => \N__57281\
        );

    \I__14283\ : Span4Mux_v
    port map (
            O => \N__57446\,
            I => \N__57278\
        );

    \I__14282\ : LocalMux
    port map (
            O => \N__57443\,
            I => \N__57263\
        );

    \I__14281\ : LocalMux
    port map (
            O => \N__57440\,
            I => \N__57263\
        );

    \I__14280\ : LocalMux
    port map (
            O => \N__57437\,
            I => \N__57263\
        );

    \I__14279\ : Span4Mux_h
    port map (
            O => \N__57434\,
            I => \N__57263\
        );

    \I__14278\ : LocalMux
    port map (
            O => \N__57423\,
            I => \N__57263\
        );

    \I__14277\ : Span4Mux_v
    port map (
            O => \N__57416\,
            I => \N__57263\
        );

    \I__14276\ : LocalMux
    port map (
            O => \N__57411\,
            I => \N__57263\
        );

    \I__14275\ : Span4Mux_h
    port map (
            O => \N__57404\,
            I => \N__57258\
        );

    \I__14274\ : LocalMux
    port map (
            O => \N__57399\,
            I => \N__57251\
        );

    \I__14273\ : LocalMux
    port map (
            O => \N__57394\,
            I => \N__57251\
        );

    \I__14272\ : LocalMux
    port map (
            O => \N__57389\,
            I => \N__57251\
        );

    \I__14271\ : InMux
    port map (
            O => \N__57388\,
            I => \N__57246\
        );

    \I__14270\ : InMux
    port map (
            O => \N__57387\,
            I => \N__57246\
        );

    \I__14269\ : InMux
    port map (
            O => \N__57386\,
            I => \N__57241\
        );

    \I__14268\ : InMux
    port map (
            O => \N__57385\,
            I => \N__57241\
        );

    \I__14267\ : InMux
    port map (
            O => \N__57384\,
            I => \N__57232\
        );

    \I__14266\ : InMux
    port map (
            O => \N__57383\,
            I => \N__57232\
        );

    \I__14265\ : InMux
    port map (
            O => \N__57382\,
            I => \N__57232\
        );

    \I__14264\ : InMux
    port map (
            O => \N__57381\,
            I => \N__57232\
        );

    \I__14263\ : Span12Mux_v
    port map (
            O => \N__57370\,
            I => \N__57225\
        );

    \I__14262\ : LocalMux
    port map (
            O => \N__57367\,
            I => \N__57225\
        );

    \I__14261\ : Span12Mux_v
    port map (
            O => \N__57362\,
            I => \N__57225\
        );

    \I__14260\ : Span12Mux_h
    port map (
            O => \N__57355\,
            I => \N__57222\
        );

    \I__14259\ : LocalMux
    port map (
            O => \N__57352\,
            I => \N__57215\
        );

    \I__14258\ : LocalMux
    port map (
            O => \N__57349\,
            I => \N__57215\
        );

    \I__14257\ : Span12Mux_h
    port map (
            O => \N__57346\,
            I => \N__57215\
        );

    \I__14256\ : Span4Mux_h
    port map (
            O => \N__57335\,
            I => \N__57208\
        );

    \I__14255\ : Span4Mux_h
    port map (
            O => \N__57330\,
            I => \N__57208\
        );

    \I__14254\ : Span4Mux_h
    port map (
            O => \N__57323\,
            I => \N__57208\
        );

    \I__14253\ : LocalMux
    port map (
            O => \N__57320\,
            I => \N__57199\
        );

    \I__14252\ : LocalMux
    port map (
            O => \N__57317\,
            I => \N__57199\
        );

    \I__14251\ : Span4Mux_h
    port map (
            O => \N__57312\,
            I => \N__57199\
        );

    \I__14250\ : Span4Mux_v
    port map (
            O => \N__57303\,
            I => \N__57199\
        );

    \I__14249\ : LocalMux
    port map (
            O => \N__57300\,
            I => \N__57186\
        );

    \I__14248\ : LocalMux
    port map (
            O => \N__57293\,
            I => \N__57186\
        );

    \I__14247\ : Span4Mux_h
    port map (
            O => \N__57288\,
            I => \N__57186\
        );

    \I__14246\ : Span4Mux_h
    port map (
            O => \N__57281\,
            I => \N__57186\
        );

    \I__14245\ : Span4Mux_v
    port map (
            O => \N__57278\,
            I => \N__57186\
        );

    \I__14244\ : Span4Mux_v
    port map (
            O => \N__57263\,
            I => \N__57186\
        );

    \I__14243\ : InMux
    port map (
            O => \N__57262\,
            I => \N__57181\
        );

    \I__14242\ : InMux
    port map (
            O => \N__57261\,
            I => \N__57181\
        );

    \I__14241\ : Odrv4
    port map (
            O => \N__57258\,
            I => comm_cmd_0
        );

    \I__14240\ : Odrv4
    port map (
            O => \N__57251\,
            I => comm_cmd_0
        );

    \I__14239\ : LocalMux
    port map (
            O => \N__57246\,
            I => comm_cmd_0
        );

    \I__14238\ : LocalMux
    port map (
            O => \N__57241\,
            I => comm_cmd_0
        );

    \I__14237\ : LocalMux
    port map (
            O => \N__57232\,
            I => comm_cmd_0
        );

    \I__14236\ : Odrv12
    port map (
            O => \N__57225\,
            I => comm_cmd_0
        );

    \I__14235\ : Odrv12
    port map (
            O => \N__57222\,
            I => comm_cmd_0
        );

    \I__14234\ : Odrv12
    port map (
            O => \N__57215\,
            I => comm_cmd_0
        );

    \I__14233\ : Odrv4
    port map (
            O => \N__57208\,
            I => comm_cmd_0
        );

    \I__14232\ : Odrv4
    port map (
            O => \N__57199\,
            I => comm_cmd_0
        );

    \I__14231\ : Odrv4
    port map (
            O => \N__57186\,
            I => comm_cmd_0
        );

    \I__14230\ : LocalMux
    port map (
            O => \N__57181\,
            I => comm_cmd_0
        );

    \I__14229\ : InMux
    port map (
            O => \N__57156\,
            I => \N__57153\
        );

    \I__14228\ : LocalMux
    port map (
            O => \N__57153\,
            I => \N__57150\
        );

    \I__14227\ : Span12Mux_v
    port map (
            O => \N__57150\,
            I => \N__57147\
        );

    \I__14226\ : Odrv12
    port map (
            O => \N__57147\,
            I => n21529
        );

    \I__14225\ : CascadeMux
    port map (
            O => \N__57144\,
            I => \N__57140\
        );

    \I__14224\ : CascadeMux
    port map (
            O => \N__57143\,
            I => \N__57135\
        );

    \I__14223\ : InMux
    port map (
            O => \N__57140\,
            I => \N__57127\
        );

    \I__14222\ : InMux
    port map (
            O => \N__57139\,
            I => \N__57127\
        );

    \I__14221\ : InMux
    port map (
            O => \N__57138\,
            I => \N__57119\
        );

    \I__14220\ : InMux
    port map (
            O => \N__57135\,
            I => \N__57115\
        );

    \I__14219\ : InMux
    port map (
            O => \N__57134\,
            I => \N__57110\
        );

    \I__14218\ : InMux
    port map (
            O => \N__57133\,
            I => \N__57110\
        );

    \I__14217\ : CascadeMux
    port map (
            O => \N__57132\,
            I => \N__57105\
        );

    \I__14216\ : LocalMux
    port map (
            O => \N__57127\,
            I => \N__57102\
        );

    \I__14215\ : InMux
    port map (
            O => \N__57126\,
            I => \N__57099\
        );

    \I__14214\ : InMux
    port map (
            O => \N__57125\,
            I => \N__57082\
        );

    \I__14213\ : InMux
    port map (
            O => \N__57124\,
            I => \N__57082\
        );

    \I__14212\ : InMux
    port map (
            O => \N__57123\,
            I => \N__57079\
        );

    \I__14211\ : InMux
    port map (
            O => \N__57122\,
            I => \N__57076\
        );

    \I__14210\ : LocalMux
    port map (
            O => \N__57119\,
            I => \N__57073\
        );

    \I__14209\ : SRMux
    port map (
            O => \N__57118\,
            I => \N__57070\
        );

    \I__14208\ : LocalMux
    port map (
            O => \N__57115\,
            I => \N__57056\
        );

    \I__14207\ : LocalMux
    port map (
            O => \N__57110\,
            I => \N__57053\
        );

    \I__14206\ : CascadeMux
    port map (
            O => \N__57109\,
            I => \N__57050\
        );

    \I__14205\ : CascadeMux
    port map (
            O => \N__57108\,
            I => \N__57046\
        );

    \I__14204\ : InMux
    port map (
            O => \N__57105\,
            I => \N__57043\
        );

    \I__14203\ : Span4Mux_v
    port map (
            O => \N__57102\,
            I => \N__57038\
        );

    \I__14202\ : LocalMux
    port map (
            O => \N__57099\,
            I => \N__57038\
        );

    \I__14201\ : InMux
    port map (
            O => \N__57098\,
            I => \N__57035\
        );

    \I__14200\ : InMux
    port map (
            O => \N__57097\,
            I => \N__57032\
        );

    \I__14199\ : InMux
    port map (
            O => \N__57096\,
            I => \N__57029\
        );

    \I__14198\ : CascadeMux
    port map (
            O => \N__57095\,
            I => \N__57025\
        );

    \I__14197\ : InMux
    port map (
            O => \N__57094\,
            I => \N__57016\
        );

    \I__14196\ : InMux
    port map (
            O => \N__57093\,
            I => \N__57016\
        );

    \I__14195\ : InMux
    port map (
            O => \N__57092\,
            I => \N__57008\
        );

    \I__14194\ : InMux
    port map (
            O => \N__57091\,
            I => \N__57008\
        );

    \I__14193\ : InMux
    port map (
            O => \N__57090\,
            I => \N__57005\
        );

    \I__14192\ : InMux
    port map (
            O => \N__57089\,
            I => \N__57001\
        );

    \I__14191\ : CascadeMux
    port map (
            O => \N__57088\,
            I => \N__56996\
        );

    \I__14190\ : CascadeMux
    port map (
            O => \N__57087\,
            I => \N__56993\
        );

    \I__14189\ : LocalMux
    port map (
            O => \N__57082\,
            I => \N__56983\
        );

    \I__14188\ : LocalMux
    port map (
            O => \N__57079\,
            I => \N__56983\
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__57076\,
            I => \N__56983\
        );

    \I__14186\ : Span4Mux_h
    port map (
            O => \N__57073\,
            I => \N__56983\
        );

    \I__14185\ : LocalMux
    port map (
            O => \N__57070\,
            I => \N__56980\
        );

    \I__14184\ : InMux
    port map (
            O => \N__57069\,
            I => \N__56973\
        );

    \I__14183\ : InMux
    port map (
            O => \N__57068\,
            I => \N__56973\
        );

    \I__14182\ : InMux
    port map (
            O => \N__57067\,
            I => \N__56973\
        );

    \I__14181\ : InMux
    port map (
            O => \N__57066\,
            I => \N__56968\
        );

    \I__14180\ : InMux
    port map (
            O => \N__57065\,
            I => \N__56968\
        );

    \I__14179\ : InMux
    port map (
            O => \N__57064\,
            I => \N__56959\
        );

    \I__14178\ : InMux
    port map (
            O => \N__57063\,
            I => \N__56959\
        );

    \I__14177\ : InMux
    port map (
            O => \N__57062\,
            I => \N__56959\
        );

    \I__14176\ : InMux
    port map (
            O => \N__57061\,
            I => \N__56959\
        );

    \I__14175\ : InMux
    port map (
            O => \N__57060\,
            I => \N__56948\
        );

    \I__14174\ : InMux
    port map (
            O => \N__57059\,
            I => \N__56948\
        );

    \I__14173\ : Span4Mux_h
    port map (
            O => \N__57056\,
            I => \N__56940\
        );

    \I__14172\ : Span4Mux_h
    port map (
            O => \N__57053\,
            I => \N__56940\
        );

    \I__14171\ : InMux
    port map (
            O => \N__57050\,
            I => \N__56937\
        );

    \I__14170\ : InMux
    port map (
            O => \N__57049\,
            I => \N__56920\
        );

    \I__14169\ : InMux
    port map (
            O => \N__57046\,
            I => \N__56917\
        );

    \I__14168\ : LocalMux
    port map (
            O => \N__57043\,
            I => \N__56914\
        );

    \I__14167\ : Span4Mux_h
    port map (
            O => \N__57038\,
            I => \N__56905\
        );

    \I__14166\ : LocalMux
    port map (
            O => \N__57035\,
            I => \N__56905\
        );

    \I__14165\ : LocalMux
    port map (
            O => \N__57032\,
            I => \N__56905\
        );

    \I__14164\ : LocalMux
    port map (
            O => \N__57029\,
            I => \N__56905\
        );

    \I__14163\ : CascadeMux
    port map (
            O => \N__57028\,
            I => \N__56902\
        );

    \I__14162\ : InMux
    port map (
            O => \N__57025\,
            I => \N__56888\
        );

    \I__14161\ : InMux
    port map (
            O => \N__57024\,
            I => \N__56888\
        );

    \I__14160\ : InMux
    port map (
            O => \N__57023\,
            I => \N__56888\
        );

    \I__14159\ : InMux
    port map (
            O => \N__57022\,
            I => \N__56888\
        );

    \I__14158\ : InMux
    port map (
            O => \N__57021\,
            I => \N__56888\
        );

    \I__14157\ : LocalMux
    port map (
            O => \N__57016\,
            I => \N__56885\
        );

    \I__14156\ : InMux
    port map (
            O => \N__57015\,
            I => \N__56878\
        );

    \I__14155\ : InMux
    port map (
            O => \N__57014\,
            I => \N__56878\
        );

    \I__14154\ : InMux
    port map (
            O => \N__57013\,
            I => \N__56878\
        );

    \I__14153\ : LocalMux
    port map (
            O => \N__57008\,
            I => \N__56875\
        );

    \I__14152\ : LocalMux
    port map (
            O => \N__57005\,
            I => \N__56872\
        );

    \I__14151\ : CascadeMux
    port map (
            O => \N__57004\,
            I => \N__56869\
        );

    \I__14150\ : LocalMux
    port map (
            O => \N__57001\,
            I => \N__56860\
        );

    \I__14149\ : InMux
    port map (
            O => \N__57000\,
            I => \N__56857\
        );

    \I__14148\ : InMux
    port map (
            O => \N__56999\,
            I => \N__56854\
        );

    \I__14147\ : InMux
    port map (
            O => \N__56996\,
            I => \N__56845\
        );

    \I__14146\ : InMux
    port map (
            O => \N__56993\,
            I => \N__56845\
        );

    \I__14145\ : InMux
    port map (
            O => \N__56992\,
            I => \N__56845\
        );

    \I__14144\ : Span4Mux_v
    port map (
            O => \N__56983\,
            I => \N__56842\
        );

    \I__14143\ : Span4Mux_v
    port map (
            O => \N__56980\,
            I => \N__56835\
        );

    \I__14142\ : LocalMux
    port map (
            O => \N__56973\,
            I => \N__56835\
        );

    \I__14141\ : LocalMux
    port map (
            O => \N__56968\,
            I => \N__56835\
        );

    \I__14140\ : LocalMux
    port map (
            O => \N__56959\,
            I => \N__56832\
        );

    \I__14139\ : InMux
    port map (
            O => \N__56958\,
            I => \N__56827\
        );

    \I__14138\ : InMux
    port map (
            O => \N__56957\,
            I => \N__56811\
        );

    \I__14137\ : InMux
    port map (
            O => \N__56956\,
            I => \N__56811\
        );

    \I__14136\ : InMux
    port map (
            O => \N__56955\,
            I => \N__56811\
        );

    \I__14135\ : InMux
    port map (
            O => \N__56954\,
            I => \N__56811\
        );

    \I__14134\ : InMux
    port map (
            O => \N__56953\,
            I => \N__56811\
        );

    \I__14133\ : LocalMux
    port map (
            O => \N__56948\,
            I => \N__56808\
        );

    \I__14132\ : InMux
    port map (
            O => \N__56947\,
            I => \N__56801\
        );

    \I__14131\ : InMux
    port map (
            O => \N__56946\,
            I => \N__56801\
        );

    \I__14130\ : InMux
    port map (
            O => \N__56945\,
            I => \N__56801\
        );

    \I__14129\ : Span4Mux_v
    port map (
            O => \N__56940\,
            I => \N__56796\
        );

    \I__14128\ : LocalMux
    port map (
            O => \N__56937\,
            I => \N__56796\
        );

    \I__14127\ : InMux
    port map (
            O => \N__56936\,
            I => \N__56787\
        );

    \I__14126\ : InMux
    port map (
            O => \N__56935\,
            I => \N__56787\
        );

    \I__14125\ : InMux
    port map (
            O => \N__56934\,
            I => \N__56787\
        );

    \I__14124\ : InMux
    port map (
            O => \N__56933\,
            I => \N__56787\
        );

    \I__14123\ : InMux
    port map (
            O => \N__56932\,
            I => \N__56778\
        );

    \I__14122\ : InMux
    port map (
            O => \N__56931\,
            I => \N__56778\
        );

    \I__14121\ : InMux
    port map (
            O => \N__56930\,
            I => \N__56778\
        );

    \I__14120\ : InMux
    port map (
            O => \N__56929\,
            I => \N__56778\
        );

    \I__14119\ : InMux
    port map (
            O => \N__56928\,
            I => \N__56773\
        );

    \I__14118\ : InMux
    port map (
            O => \N__56927\,
            I => \N__56773\
        );

    \I__14117\ : InMux
    port map (
            O => \N__56926\,
            I => \N__56768\
        );

    \I__14116\ : InMux
    port map (
            O => \N__56925\,
            I => \N__56768\
        );

    \I__14115\ : InMux
    port map (
            O => \N__56924\,
            I => \N__56763\
        );

    \I__14114\ : InMux
    port map (
            O => \N__56923\,
            I => \N__56763\
        );

    \I__14113\ : LocalMux
    port map (
            O => \N__56920\,
            I => \N__56760\
        );

    \I__14112\ : LocalMux
    port map (
            O => \N__56917\,
            I => \N__56757\
        );

    \I__14111\ : Span4Mux_h
    port map (
            O => \N__56914\,
            I => \N__56752\
        );

    \I__14110\ : Span4Mux_v
    port map (
            O => \N__56905\,
            I => \N__56752\
        );

    \I__14109\ : InMux
    port map (
            O => \N__56902\,
            I => \N__56743\
        );

    \I__14108\ : InMux
    port map (
            O => \N__56901\,
            I => \N__56743\
        );

    \I__14107\ : InMux
    port map (
            O => \N__56900\,
            I => \N__56743\
        );

    \I__14106\ : InMux
    port map (
            O => \N__56899\,
            I => \N__56743\
        );

    \I__14105\ : LocalMux
    port map (
            O => \N__56888\,
            I => \N__56732\
        );

    \I__14104\ : Span4Mux_h
    port map (
            O => \N__56885\,
            I => \N__56732\
        );

    \I__14103\ : LocalMux
    port map (
            O => \N__56878\,
            I => \N__56732\
        );

    \I__14102\ : Span4Mux_h
    port map (
            O => \N__56875\,
            I => \N__56732\
        );

    \I__14101\ : Span4Mux_v
    port map (
            O => \N__56872\,
            I => \N__56732\
        );

    \I__14100\ : InMux
    port map (
            O => \N__56869\,
            I => \N__56727\
        );

    \I__14099\ : InMux
    port map (
            O => \N__56868\,
            I => \N__56727\
        );

    \I__14098\ : InMux
    port map (
            O => \N__56867\,
            I => \N__56724\
        );

    \I__14097\ : InMux
    port map (
            O => \N__56866\,
            I => \N__56715\
        );

    \I__14096\ : InMux
    port map (
            O => \N__56865\,
            I => \N__56715\
        );

    \I__14095\ : InMux
    port map (
            O => \N__56864\,
            I => \N__56715\
        );

    \I__14094\ : InMux
    port map (
            O => \N__56863\,
            I => \N__56715\
        );

    \I__14093\ : Sp12to4
    port map (
            O => \N__56860\,
            I => \N__56708\
        );

    \I__14092\ : LocalMux
    port map (
            O => \N__56857\,
            I => \N__56708\
        );

    \I__14091\ : LocalMux
    port map (
            O => \N__56854\,
            I => \N__56708\
        );

    \I__14090\ : InMux
    port map (
            O => \N__56853\,
            I => \N__56703\
        );

    \I__14089\ : InMux
    port map (
            O => \N__56852\,
            I => \N__56703\
        );

    \I__14088\ : LocalMux
    port map (
            O => \N__56845\,
            I => \N__56694\
        );

    \I__14087\ : Span4Mux_v
    port map (
            O => \N__56842\,
            I => \N__56694\
        );

    \I__14086\ : Span4Mux_h
    port map (
            O => \N__56835\,
            I => \N__56694\
        );

    \I__14085\ : Span4Mux_h
    port map (
            O => \N__56832\,
            I => \N__56694\
        );

    \I__14084\ : InMux
    port map (
            O => \N__56831\,
            I => \N__56689\
        );

    \I__14083\ : InMux
    port map (
            O => \N__56830\,
            I => \N__56686\
        );

    \I__14082\ : LocalMux
    port map (
            O => \N__56827\,
            I => \N__56683\
        );

    \I__14081\ : InMux
    port map (
            O => \N__56826\,
            I => \N__56676\
        );

    \I__14080\ : InMux
    port map (
            O => \N__56825\,
            I => \N__56676\
        );

    \I__14079\ : InMux
    port map (
            O => \N__56824\,
            I => \N__56676\
        );

    \I__14078\ : InMux
    port map (
            O => \N__56823\,
            I => \N__56671\
        );

    \I__14077\ : InMux
    port map (
            O => \N__56822\,
            I => \N__56671\
        );

    \I__14076\ : LocalMux
    port map (
            O => \N__56811\,
            I => \N__56668\
        );

    \I__14075\ : Sp12to4
    port map (
            O => \N__56808\,
            I => \N__56651\
        );

    \I__14074\ : LocalMux
    port map (
            O => \N__56801\,
            I => \N__56651\
        );

    \I__14073\ : Sp12to4
    port map (
            O => \N__56796\,
            I => \N__56651\
        );

    \I__14072\ : LocalMux
    port map (
            O => \N__56787\,
            I => \N__56651\
        );

    \I__14071\ : LocalMux
    port map (
            O => \N__56778\,
            I => \N__56651\
        );

    \I__14070\ : LocalMux
    port map (
            O => \N__56773\,
            I => \N__56651\
        );

    \I__14069\ : LocalMux
    port map (
            O => \N__56768\,
            I => \N__56651\
        );

    \I__14068\ : LocalMux
    port map (
            O => \N__56763\,
            I => \N__56651\
        );

    \I__14067\ : Span4Mux_h
    port map (
            O => \N__56760\,
            I => \N__56640\
        );

    \I__14066\ : Span4Mux_v
    port map (
            O => \N__56757\,
            I => \N__56640\
        );

    \I__14065\ : Span4Mux_h
    port map (
            O => \N__56752\,
            I => \N__56640\
        );

    \I__14064\ : LocalMux
    port map (
            O => \N__56743\,
            I => \N__56640\
        );

    \I__14063\ : Span4Mux_v
    port map (
            O => \N__56732\,
            I => \N__56640\
        );

    \I__14062\ : LocalMux
    port map (
            O => \N__56727\,
            I => \N__56629\
        );

    \I__14061\ : LocalMux
    port map (
            O => \N__56724\,
            I => \N__56629\
        );

    \I__14060\ : LocalMux
    port map (
            O => \N__56715\,
            I => \N__56629\
        );

    \I__14059\ : Span12Mux_v
    port map (
            O => \N__56708\,
            I => \N__56629\
        );

    \I__14058\ : LocalMux
    port map (
            O => \N__56703\,
            I => \N__56629\
        );

    \I__14057\ : Span4Mux_h
    port map (
            O => \N__56694\,
            I => \N__56626\
        );

    \I__14056\ : InMux
    port map (
            O => \N__56693\,
            I => \N__56621\
        );

    \I__14055\ : InMux
    port map (
            O => \N__56692\,
            I => \N__56621\
        );

    \I__14054\ : LocalMux
    port map (
            O => \N__56689\,
            I => comm_state_3
        );

    \I__14053\ : LocalMux
    port map (
            O => \N__56686\,
            I => comm_state_3
        );

    \I__14052\ : Odrv4
    port map (
            O => \N__56683\,
            I => comm_state_3
        );

    \I__14051\ : LocalMux
    port map (
            O => \N__56676\,
            I => comm_state_3
        );

    \I__14050\ : LocalMux
    port map (
            O => \N__56671\,
            I => comm_state_3
        );

    \I__14049\ : Odrv4
    port map (
            O => \N__56668\,
            I => comm_state_3
        );

    \I__14048\ : Odrv12
    port map (
            O => \N__56651\,
            I => comm_state_3
        );

    \I__14047\ : Odrv4
    port map (
            O => \N__56640\,
            I => comm_state_3
        );

    \I__14046\ : Odrv12
    port map (
            O => \N__56629\,
            I => comm_state_3
        );

    \I__14045\ : Odrv4
    port map (
            O => \N__56626\,
            I => comm_state_3
        );

    \I__14044\ : LocalMux
    port map (
            O => \N__56621\,
            I => comm_state_3
        );

    \I__14043\ : CascadeMux
    port map (
            O => \N__56598\,
            I => \N__56595\
        );

    \I__14042\ : InMux
    port map (
            O => \N__56595\,
            I => \N__56591\
        );

    \I__14041\ : InMux
    port map (
            O => \N__56594\,
            I => \N__56588\
        );

    \I__14040\ : LocalMux
    port map (
            O => \N__56591\,
            I => \N__56585\
        );

    \I__14039\ : LocalMux
    port map (
            O => \N__56588\,
            I => \N__56582\
        );

    \I__14038\ : Span4Mux_v
    port map (
            O => \N__56585\,
            I => \N__56579\
        );

    \I__14037\ : Span4Mux_v
    port map (
            O => \N__56582\,
            I => \N__56576\
        );

    \I__14036\ : Span4Mux_h
    port map (
            O => \N__56579\,
            I => \N__56571\
        );

    \I__14035\ : Span4Mux_h
    port map (
            O => \N__56576\,
            I => \N__56571\
        );

    \I__14034\ : Odrv4
    port map (
            O => \N__56571\,
            I => n17489
        );

    \I__14033\ : CascadeMux
    port map (
            O => \N__56568\,
            I => \N__56564\
        );

    \I__14032\ : CascadeMux
    port map (
            O => \N__56567\,
            I => \N__56541\
        );

    \I__14031\ : InMux
    port map (
            O => \N__56564\,
            I => \N__56532\
        );

    \I__14030\ : InMux
    port map (
            O => \N__56563\,
            I => \N__56532\
        );

    \I__14029\ : InMux
    port map (
            O => \N__56562\,
            I => \N__56532\
        );

    \I__14028\ : InMux
    port map (
            O => \N__56561\,
            I => \N__56527\
        );

    \I__14027\ : InMux
    port map (
            O => \N__56560\,
            I => \N__56527\
        );

    \I__14026\ : InMux
    port map (
            O => \N__56559\,
            I => \N__56520\
        );

    \I__14025\ : InMux
    port map (
            O => \N__56558\,
            I => \N__56520\
        );

    \I__14024\ : InMux
    port map (
            O => \N__56557\,
            I => \N__56520\
        );

    \I__14023\ : CascadeMux
    port map (
            O => \N__56556\,
            I => \N__56513\
        );

    \I__14022\ : InMux
    port map (
            O => \N__56555\,
            I => \N__56509\
        );

    \I__14021\ : InMux
    port map (
            O => \N__56554\,
            I => \N__56506\
        );

    \I__14020\ : CascadeMux
    port map (
            O => \N__56553\,
            I => \N__56501\
        );

    \I__14019\ : InMux
    port map (
            O => \N__56552\,
            I => \N__56494\
        );

    \I__14018\ : InMux
    port map (
            O => \N__56551\,
            I => \N__56489\
        );

    \I__14017\ : InMux
    port map (
            O => \N__56550\,
            I => \N__56489\
        );

    \I__14016\ : CascadeMux
    port map (
            O => \N__56549\,
            I => \N__56485\
        );

    \I__14015\ : CascadeMux
    port map (
            O => \N__56548\,
            I => \N__56468\
        );

    \I__14014\ : InMux
    port map (
            O => \N__56547\,
            I => \N__56459\
        );

    \I__14013\ : InMux
    port map (
            O => \N__56546\,
            I => \N__56459\
        );

    \I__14012\ : InMux
    port map (
            O => \N__56545\,
            I => \N__56459\
        );

    \I__14011\ : InMux
    port map (
            O => \N__56544\,
            I => \N__56456\
        );

    \I__14010\ : InMux
    port map (
            O => \N__56541\,
            I => \N__56453\
        );

    \I__14009\ : CascadeMux
    port map (
            O => \N__56540\,
            I => \N__56447\
        );

    \I__14008\ : CascadeMux
    port map (
            O => \N__56539\,
            I => \N__56442\
        );

    \I__14007\ : LocalMux
    port map (
            O => \N__56532\,
            I => \N__56433\
        );

    \I__14006\ : LocalMux
    port map (
            O => \N__56527\,
            I => \N__56433\
        );

    \I__14005\ : LocalMux
    port map (
            O => \N__56520\,
            I => \N__56433\
        );

    \I__14004\ : InMux
    port map (
            O => \N__56519\,
            I => \N__56430\
        );

    \I__14003\ : CascadeMux
    port map (
            O => \N__56518\,
            I => \N__56427\
        );

    \I__14002\ : CascadeMux
    port map (
            O => \N__56517\,
            I => \N__56424\
        );

    \I__14001\ : CascadeMux
    port map (
            O => \N__56516\,
            I => \N__56421\
        );

    \I__14000\ : InMux
    port map (
            O => \N__56513\,
            I => \N__56414\
        );

    \I__13999\ : InMux
    port map (
            O => \N__56512\,
            I => \N__56414\
        );

    \I__13998\ : LocalMux
    port map (
            O => \N__56509\,
            I => \N__56409\
        );

    \I__13997\ : LocalMux
    port map (
            O => \N__56506\,
            I => \N__56409\
        );

    \I__13996\ : InMux
    port map (
            O => \N__56505\,
            I => \N__56406\
        );

    \I__13995\ : InMux
    port map (
            O => \N__56504\,
            I => \N__56401\
        );

    \I__13994\ : InMux
    port map (
            O => \N__56501\,
            I => \N__56401\
        );

    \I__13993\ : InMux
    port map (
            O => \N__56500\,
            I => \N__56395\
        );

    \I__13992\ : InMux
    port map (
            O => \N__56499\,
            I => \N__56395\
        );

    \I__13991\ : InMux
    port map (
            O => \N__56498\,
            I => \N__56390\
        );

    \I__13990\ : InMux
    port map (
            O => \N__56497\,
            I => \N__56390\
        );

    \I__13989\ : LocalMux
    port map (
            O => \N__56494\,
            I => \N__56387\
        );

    \I__13988\ : LocalMux
    port map (
            O => \N__56489\,
            I => \N__56384\
        );

    \I__13987\ : InMux
    port map (
            O => \N__56488\,
            I => \N__56379\
        );

    \I__13986\ : InMux
    port map (
            O => \N__56485\,
            I => \N__56379\
        );

    \I__13985\ : InMux
    port map (
            O => \N__56484\,
            I => \N__56364\
        );

    \I__13984\ : InMux
    port map (
            O => \N__56483\,
            I => \N__56364\
        );

    \I__13983\ : InMux
    port map (
            O => \N__56482\,
            I => \N__56364\
        );

    \I__13982\ : InMux
    port map (
            O => \N__56481\,
            I => \N__56364\
        );

    \I__13981\ : InMux
    port map (
            O => \N__56480\,
            I => \N__56364\
        );

    \I__13980\ : InMux
    port map (
            O => \N__56479\,
            I => \N__56364\
        );

    \I__13979\ : InMux
    port map (
            O => \N__56478\,
            I => \N__56364\
        );

    \I__13978\ : CascadeMux
    port map (
            O => \N__56477\,
            I => \N__56361\
        );

    \I__13977\ : CascadeMux
    port map (
            O => \N__56476\,
            I => \N__56358\
        );

    \I__13976\ : InMux
    port map (
            O => \N__56475\,
            I => \N__56351\
        );

    \I__13975\ : InMux
    port map (
            O => \N__56474\,
            I => \N__56351\
        );

    \I__13974\ : CascadeMux
    port map (
            O => \N__56473\,
            I => \N__56348\
        );

    \I__13973\ : CascadeMux
    port map (
            O => \N__56472\,
            I => \N__56345\
        );

    \I__13972\ : InMux
    port map (
            O => \N__56471\,
            I => \N__56334\
        );

    \I__13971\ : InMux
    port map (
            O => \N__56468\,
            I => \N__56334\
        );

    \I__13970\ : InMux
    port map (
            O => \N__56467\,
            I => \N__56334\
        );

    \I__13969\ : InMux
    port map (
            O => \N__56466\,
            I => \N__56334\
        );

    \I__13968\ : LocalMux
    port map (
            O => \N__56459\,
            I => \N__56331\
        );

    \I__13967\ : LocalMux
    port map (
            O => \N__56456\,
            I => \N__56328\
        );

    \I__13966\ : LocalMux
    port map (
            O => \N__56453\,
            I => \N__56325\
        );

    \I__13965\ : InMux
    port map (
            O => \N__56452\,
            I => \N__56322\
        );

    \I__13964\ : InMux
    port map (
            O => \N__56451\,
            I => \N__56317\
        );

    \I__13963\ : InMux
    port map (
            O => \N__56450\,
            I => \N__56312\
        );

    \I__13962\ : InMux
    port map (
            O => \N__56447\,
            I => \N__56305\
        );

    \I__13961\ : InMux
    port map (
            O => \N__56446\,
            I => \N__56305\
        );

    \I__13960\ : InMux
    port map (
            O => \N__56445\,
            I => \N__56305\
        );

    \I__13959\ : InMux
    port map (
            O => \N__56442\,
            I => \N__56298\
        );

    \I__13958\ : InMux
    port map (
            O => \N__56441\,
            I => \N__56298\
        );

    \I__13957\ : InMux
    port map (
            O => \N__56440\,
            I => \N__56298\
        );

    \I__13956\ : Span4Mux_v
    port map (
            O => \N__56433\,
            I => \N__56293\
        );

    \I__13955\ : LocalMux
    port map (
            O => \N__56430\,
            I => \N__56293\
        );

    \I__13954\ : InMux
    port map (
            O => \N__56427\,
            I => \N__56288\
        );

    \I__13953\ : InMux
    port map (
            O => \N__56424\,
            I => \N__56281\
        );

    \I__13952\ : InMux
    port map (
            O => \N__56421\,
            I => \N__56281\
        );

    \I__13951\ : InMux
    port map (
            O => \N__56420\,
            I => \N__56281\
        );

    \I__13950\ : InMux
    port map (
            O => \N__56419\,
            I => \N__56278\
        );

    \I__13949\ : LocalMux
    port map (
            O => \N__56414\,
            I => \N__56275\
        );

    \I__13948\ : Span4Mux_v
    port map (
            O => \N__56409\,
            I => \N__56272\
        );

    \I__13947\ : LocalMux
    port map (
            O => \N__56406\,
            I => \N__56267\
        );

    \I__13946\ : LocalMux
    port map (
            O => \N__56401\,
            I => \N__56267\
        );

    \I__13945\ : InMux
    port map (
            O => \N__56400\,
            I => \N__56264\
        );

    \I__13944\ : LocalMux
    port map (
            O => \N__56395\,
            I => \N__56253\
        );

    \I__13943\ : LocalMux
    port map (
            O => \N__56390\,
            I => \N__56253\
        );

    \I__13942\ : Span4Mux_h
    port map (
            O => \N__56387\,
            I => \N__56253\
        );

    \I__13941\ : Span4Mux_h
    port map (
            O => \N__56384\,
            I => \N__56253\
        );

    \I__13940\ : LocalMux
    port map (
            O => \N__56379\,
            I => \N__56253\
        );

    \I__13939\ : LocalMux
    port map (
            O => \N__56364\,
            I => \N__56250\
        );

    \I__13938\ : InMux
    port map (
            O => \N__56361\,
            I => \N__56247\
        );

    \I__13937\ : InMux
    port map (
            O => \N__56358\,
            I => \N__56240\
        );

    \I__13936\ : InMux
    port map (
            O => \N__56357\,
            I => \N__56240\
        );

    \I__13935\ : InMux
    port map (
            O => \N__56356\,
            I => \N__56240\
        );

    \I__13934\ : LocalMux
    port map (
            O => \N__56351\,
            I => \N__56237\
        );

    \I__13933\ : InMux
    port map (
            O => \N__56348\,
            I => \N__56232\
        );

    \I__13932\ : InMux
    port map (
            O => \N__56345\,
            I => \N__56232\
        );

    \I__13931\ : CascadeMux
    port map (
            O => \N__56344\,
            I => \N__56229\
        );

    \I__13930\ : CascadeMux
    port map (
            O => \N__56343\,
            I => \N__56224\
        );

    \I__13929\ : LocalMux
    port map (
            O => \N__56334\,
            I => \N__56215\
        );

    \I__13928\ : Span4Mux_v
    port map (
            O => \N__56331\,
            I => \N__56215\
        );

    \I__13927\ : Span4Mux_h
    port map (
            O => \N__56328\,
            I => \N__56212\
        );

    \I__13926\ : Span4Mux_h
    port map (
            O => \N__56325\,
            I => \N__56207\
        );

    \I__13925\ : LocalMux
    port map (
            O => \N__56322\,
            I => \N__56207\
        );

    \I__13924\ : CascadeMux
    port map (
            O => \N__56321\,
            I => \N__56204\
        );

    \I__13923\ : CascadeMux
    port map (
            O => \N__56320\,
            I => \N__56199\
        );

    \I__13922\ : LocalMux
    port map (
            O => \N__56317\,
            I => \N__56196\
        );

    \I__13921\ : InMux
    port map (
            O => \N__56316\,
            I => \N__56191\
        );

    \I__13920\ : InMux
    port map (
            O => \N__56315\,
            I => \N__56191\
        );

    \I__13919\ : LocalMux
    port map (
            O => \N__56312\,
            I => \N__56188\
        );

    \I__13918\ : LocalMux
    port map (
            O => \N__56305\,
            I => \N__56181\
        );

    \I__13917\ : LocalMux
    port map (
            O => \N__56298\,
            I => \N__56181\
        );

    \I__13916\ : Span4Mux_h
    port map (
            O => \N__56293\,
            I => \N__56181\
        );

    \I__13915\ : CascadeMux
    port map (
            O => \N__56292\,
            I => \N__56176\
        );

    \I__13914\ : CascadeMux
    port map (
            O => \N__56291\,
            I => \N__56171\
        );

    \I__13913\ : LocalMux
    port map (
            O => \N__56288\,
            I => \N__56165\
        );

    \I__13912\ : LocalMux
    port map (
            O => \N__56281\,
            I => \N__56160\
        );

    \I__13911\ : LocalMux
    port map (
            O => \N__56278\,
            I => \N__56160\
        );

    \I__13910\ : Span4Mux_v
    port map (
            O => \N__56275\,
            I => \N__56157\
        );

    \I__13909\ : Span4Mux_h
    port map (
            O => \N__56272\,
            I => \N__56146\
        );

    \I__13908\ : Span4Mux_v
    port map (
            O => \N__56267\,
            I => \N__56146\
        );

    \I__13907\ : LocalMux
    port map (
            O => \N__56264\,
            I => \N__56146\
        );

    \I__13906\ : Span4Mux_v
    port map (
            O => \N__56253\,
            I => \N__56146\
        );

    \I__13905\ : Span4Mux_v
    port map (
            O => \N__56250\,
            I => \N__56146\
        );

    \I__13904\ : LocalMux
    port map (
            O => \N__56247\,
            I => \N__56143\
        );

    \I__13903\ : LocalMux
    port map (
            O => \N__56240\,
            I => \N__56136\
        );

    \I__13902\ : Span4Mux_v
    port map (
            O => \N__56237\,
            I => \N__56136\
        );

    \I__13901\ : LocalMux
    port map (
            O => \N__56232\,
            I => \N__56136\
        );

    \I__13900\ : InMux
    port map (
            O => \N__56229\,
            I => \N__56129\
        );

    \I__13899\ : InMux
    port map (
            O => \N__56228\,
            I => \N__56129\
        );

    \I__13898\ : InMux
    port map (
            O => \N__56227\,
            I => \N__56129\
        );

    \I__13897\ : InMux
    port map (
            O => \N__56224\,
            I => \N__56124\
        );

    \I__13896\ : InMux
    port map (
            O => \N__56223\,
            I => \N__56124\
        );

    \I__13895\ : InMux
    port map (
            O => \N__56222\,
            I => \N__56121\
        );

    \I__13894\ : InMux
    port map (
            O => \N__56221\,
            I => \N__56116\
        );

    \I__13893\ : InMux
    port map (
            O => \N__56220\,
            I => \N__56116\
        );

    \I__13892\ : Span4Mux_h
    port map (
            O => \N__56215\,
            I => \N__56109\
        );

    \I__13891\ : Span4Mux_v
    port map (
            O => \N__56212\,
            I => \N__56109\
        );

    \I__13890\ : Span4Mux_v
    port map (
            O => \N__56207\,
            I => \N__56109\
        );

    \I__13889\ : InMux
    port map (
            O => \N__56204\,
            I => \N__56100\
        );

    \I__13888\ : InMux
    port map (
            O => \N__56203\,
            I => \N__56100\
        );

    \I__13887\ : InMux
    port map (
            O => \N__56202\,
            I => \N__56100\
        );

    \I__13886\ : InMux
    port map (
            O => \N__56199\,
            I => \N__56100\
        );

    \I__13885\ : Span4Mux_h
    port map (
            O => \N__56196\,
            I => \N__56091\
        );

    \I__13884\ : LocalMux
    port map (
            O => \N__56191\,
            I => \N__56091\
        );

    \I__13883\ : Span4Mux_v
    port map (
            O => \N__56188\,
            I => \N__56091\
        );

    \I__13882\ : Span4Mux_h
    port map (
            O => \N__56181\,
            I => \N__56091\
        );

    \I__13881\ : InMux
    port map (
            O => \N__56180\,
            I => \N__56084\
        );

    \I__13880\ : InMux
    port map (
            O => \N__56179\,
            I => \N__56084\
        );

    \I__13879\ : InMux
    port map (
            O => \N__56176\,
            I => \N__56084\
        );

    \I__13878\ : InMux
    port map (
            O => \N__56175\,
            I => \N__56075\
        );

    \I__13877\ : InMux
    port map (
            O => \N__56174\,
            I => \N__56075\
        );

    \I__13876\ : InMux
    port map (
            O => \N__56171\,
            I => \N__56075\
        );

    \I__13875\ : InMux
    port map (
            O => \N__56170\,
            I => \N__56075\
        );

    \I__13874\ : InMux
    port map (
            O => \N__56169\,
            I => \N__56070\
        );

    \I__13873\ : InMux
    port map (
            O => \N__56168\,
            I => \N__56070\
        );

    \I__13872\ : Span4Mux_h
    port map (
            O => \N__56165\,
            I => \N__56065\
        );

    \I__13871\ : Span4Mux_h
    port map (
            O => \N__56160\,
            I => \N__56065\
        );

    \I__13870\ : Span4Mux_v
    port map (
            O => \N__56157\,
            I => \N__56054\
        );

    \I__13869\ : Span4Mux_h
    port map (
            O => \N__56146\,
            I => \N__56054\
        );

    \I__13868\ : Span4Mux_v
    port map (
            O => \N__56143\,
            I => \N__56054\
        );

    \I__13867\ : Span4Mux_v
    port map (
            O => \N__56136\,
            I => \N__56054\
        );

    \I__13866\ : LocalMux
    port map (
            O => \N__56129\,
            I => \N__56054\
        );

    \I__13865\ : LocalMux
    port map (
            O => \N__56124\,
            I => n9306
        );

    \I__13864\ : LocalMux
    port map (
            O => \N__56121\,
            I => n9306
        );

    \I__13863\ : LocalMux
    port map (
            O => \N__56116\,
            I => n9306
        );

    \I__13862\ : Odrv4
    port map (
            O => \N__56109\,
            I => n9306
        );

    \I__13861\ : LocalMux
    port map (
            O => \N__56100\,
            I => n9306
        );

    \I__13860\ : Odrv4
    port map (
            O => \N__56091\,
            I => n9306
        );

    \I__13859\ : LocalMux
    port map (
            O => \N__56084\,
            I => n9306
        );

    \I__13858\ : LocalMux
    port map (
            O => \N__56075\,
            I => n9306
        );

    \I__13857\ : LocalMux
    port map (
            O => \N__56070\,
            I => n9306
        );

    \I__13856\ : Odrv4
    port map (
            O => \N__56065\,
            I => n9306
        );

    \I__13855\ : Odrv4
    port map (
            O => \N__56054\,
            I => n9306
        );

    \I__13854\ : InMux
    port map (
            O => \N__56031\,
            I => \N__56027\
        );

    \I__13853\ : InMux
    port map (
            O => \N__56030\,
            I => \N__56024\
        );

    \I__13852\ : LocalMux
    port map (
            O => \N__56027\,
            I => \N__56021\
        );

    \I__13851\ : LocalMux
    port map (
            O => \N__56024\,
            I => \N__56018\
        );

    \I__13850\ : Span4Mux_v
    port map (
            O => \N__56021\,
            I => \N__56015\
        );

    \I__13849\ : Span4Mux_v
    port map (
            O => \N__56018\,
            I => \N__56010\
        );

    \I__13848\ : Span4Mux_h
    port map (
            O => \N__56015\,
            I => \N__56010\
        );

    \I__13847\ : Odrv4
    port map (
            O => \N__56010\,
            I => n17487
        );

    \I__13846\ : CascadeMux
    port map (
            O => \N__56007\,
            I => \N__56004\
        );

    \I__13845\ : CascadeBuf
    port map (
            O => \N__56004\,
            I => \N__56001\
        );

    \I__13844\ : CascadeMux
    port map (
            O => \N__56001\,
            I => \N__55998\
        );

    \I__13843\ : CascadeBuf
    port map (
            O => \N__55998\,
            I => \N__55995\
        );

    \I__13842\ : CascadeMux
    port map (
            O => \N__55995\,
            I => \N__55992\
        );

    \I__13841\ : CascadeBuf
    port map (
            O => \N__55992\,
            I => \N__55989\
        );

    \I__13840\ : CascadeMux
    port map (
            O => \N__55989\,
            I => \N__55986\
        );

    \I__13839\ : CascadeBuf
    port map (
            O => \N__55986\,
            I => \N__55983\
        );

    \I__13838\ : CascadeMux
    port map (
            O => \N__55983\,
            I => \N__55980\
        );

    \I__13837\ : CascadeBuf
    port map (
            O => \N__55980\,
            I => \N__55977\
        );

    \I__13836\ : CascadeMux
    port map (
            O => \N__55977\,
            I => \N__55974\
        );

    \I__13835\ : CascadeBuf
    port map (
            O => \N__55974\,
            I => \N__55971\
        );

    \I__13834\ : CascadeMux
    port map (
            O => \N__55971\,
            I => \N__55968\
        );

    \I__13833\ : CascadeBuf
    port map (
            O => \N__55968\,
            I => \N__55964\
        );

    \I__13832\ : CascadeMux
    port map (
            O => \N__55967\,
            I => \N__55961\
        );

    \I__13831\ : CascadeMux
    port map (
            O => \N__55964\,
            I => \N__55958\
        );

    \I__13830\ : CascadeBuf
    port map (
            O => \N__55961\,
            I => \N__55955\
        );

    \I__13829\ : CascadeBuf
    port map (
            O => \N__55958\,
            I => \N__55952\
        );

    \I__13828\ : CascadeMux
    port map (
            O => \N__55955\,
            I => \N__55949\
        );

    \I__13827\ : CascadeMux
    port map (
            O => \N__55952\,
            I => \N__55946\
        );

    \I__13826\ : InMux
    port map (
            O => \N__55949\,
            I => \N__55943\
        );

    \I__13825\ : CascadeBuf
    port map (
            O => \N__55946\,
            I => \N__55940\
        );

    \I__13824\ : LocalMux
    port map (
            O => \N__55943\,
            I => \N__55937\
        );

    \I__13823\ : CascadeMux
    port map (
            O => \N__55940\,
            I => \N__55934\
        );

    \I__13822\ : Span12Mux_h
    port map (
            O => \N__55937\,
            I => \N__55931\
        );

    \I__13821\ : InMux
    port map (
            O => \N__55934\,
            I => \N__55928\
        );

    \I__13820\ : Span12Mux_v
    port map (
            O => \N__55931\,
            I => \N__55925\
        );

    \I__13819\ : LocalMux
    port map (
            O => \N__55928\,
            I => \N__55922\
        );

    \I__13818\ : Odrv12
    port map (
            O => \N__55925\,
            I => \data_index_9_N_216_5\
        );

    \I__13817\ : Odrv4
    port map (
            O => \N__55922\,
            I => \data_index_9_N_216_5\
        );

    \I__13816\ : InMux
    port map (
            O => \N__55917\,
            I => \bfn_22_7_0_\
        );

    \I__13815\ : InMux
    port map (
            O => \N__55914\,
            I => \ADC_VDC.genclk.n19724\
        );

    \I__13814\ : InMux
    port map (
            O => \N__55911\,
            I => \ADC_VDC.genclk.n19725\
        );

    \I__13813\ : InMux
    port map (
            O => \N__55908\,
            I => \ADC_VDC.genclk.n19726\
        );

    \I__13812\ : InMux
    port map (
            O => \N__55905\,
            I => \ADC_VDC.genclk.n19727\
        );

    \I__13811\ : InMux
    port map (
            O => \N__55902\,
            I => \N__55897\
        );

    \I__13810\ : InMux
    port map (
            O => \N__55901\,
            I => \N__55894\
        );

    \I__13809\ : InMux
    port map (
            O => \N__55900\,
            I => \N__55891\
        );

    \I__13808\ : LocalMux
    port map (
            O => \N__55897\,
            I => \N__55888\
        );

    \I__13807\ : LocalMux
    port map (
            O => \N__55894\,
            I => \N__55885\
        );

    \I__13806\ : LocalMux
    port map (
            O => \N__55891\,
            I => \N__55882\
        );

    \I__13805\ : Odrv4
    port map (
            O => \N__55888\,
            I => \comm_spi.n14600\
        );

    \I__13804\ : Odrv4
    port map (
            O => \N__55885\,
            I => \comm_spi.n14600\
        );

    \I__13803\ : Odrv4
    port map (
            O => \N__55882\,
            I => \comm_spi.n14600\
        );

    \I__13802\ : InMux
    port map (
            O => \N__55875\,
            I => \N__55862\
        );

    \I__13801\ : InMux
    port map (
            O => \N__55874\,
            I => \N__55859\
        );

    \I__13800\ : CascadeMux
    port map (
            O => \N__55873\,
            I => \N__55854\
        );

    \I__13799\ : CascadeMux
    port map (
            O => \N__55872\,
            I => \N__55851\
        );

    \I__13798\ : CascadeMux
    port map (
            O => \N__55871\,
            I => \N__55844\
        );

    \I__13797\ : SRMux
    port map (
            O => \N__55870\,
            I => \N__55840\
        );

    \I__13796\ : SRMux
    port map (
            O => \N__55869\,
            I => \N__55837\
        );

    \I__13795\ : InMux
    port map (
            O => \N__55868\,
            I => \N__55834\
        );

    \I__13794\ : InMux
    port map (
            O => \N__55867\,
            I => \N__55828\
        );

    \I__13793\ : InMux
    port map (
            O => \N__55866\,
            I => \N__55824\
        );

    \I__13792\ : InMux
    port map (
            O => \N__55865\,
            I => \N__55821\
        );

    \I__13791\ : LocalMux
    port map (
            O => \N__55862\,
            I => \N__55811\
        );

    \I__13790\ : LocalMux
    port map (
            O => \N__55859\,
            I => \N__55811\
        );

    \I__13789\ : InMux
    port map (
            O => \N__55858\,
            I => \N__55795\
        );

    \I__13788\ : InMux
    port map (
            O => \N__55857\,
            I => \N__55795\
        );

    \I__13787\ : InMux
    port map (
            O => \N__55854\,
            I => \N__55795\
        );

    \I__13786\ : InMux
    port map (
            O => \N__55851\,
            I => \N__55795\
        );

    \I__13785\ : InMux
    port map (
            O => \N__55850\,
            I => \N__55795\
        );

    \I__13784\ : InMux
    port map (
            O => \N__55849\,
            I => \N__55795\
        );

    \I__13783\ : InMux
    port map (
            O => \N__55848\,
            I => \N__55795\
        );

    \I__13782\ : InMux
    port map (
            O => \N__55847\,
            I => \N__55792\
        );

    \I__13781\ : InMux
    port map (
            O => \N__55844\,
            I => \N__55787\
        );

    \I__13780\ : InMux
    port map (
            O => \N__55843\,
            I => \N__55787\
        );

    \I__13779\ : LocalMux
    port map (
            O => \N__55840\,
            I => \N__55782\
        );

    \I__13778\ : LocalMux
    port map (
            O => \N__55837\,
            I => \N__55782\
        );

    \I__13777\ : LocalMux
    port map (
            O => \N__55834\,
            I => \N__55779\
        );

    \I__13776\ : InMux
    port map (
            O => \N__55833\,
            I => \N__55772\
        );

    \I__13775\ : InMux
    port map (
            O => \N__55832\,
            I => \N__55772\
        );

    \I__13774\ : InMux
    port map (
            O => \N__55831\,
            I => \N__55769\
        );

    \I__13773\ : LocalMux
    port map (
            O => \N__55828\,
            I => \N__55766\
        );

    \I__13772\ : InMux
    port map (
            O => \N__55827\,
            I => \N__55760\
        );

    \I__13771\ : LocalMux
    port map (
            O => \N__55824\,
            I => \N__55752\
        );

    \I__13770\ : LocalMux
    port map (
            O => \N__55821\,
            I => \N__55752\
        );

    \I__13769\ : SRMux
    port map (
            O => \N__55820\,
            I => \N__55749\
        );

    \I__13768\ : InMux
    port map (
            O => \N__55819\,
            I => \N__55742\
        );

    \I__13767\ : InMux
    port map (
            O => \N__55818\,
            I => \N__55742\
        );

    \I__13766\ : InMux
    port map (
            O => \N__55817\,
            I => \N__55742\
        );

    \I__13765\ : InMux
    port map (
            O => \N__55816\,
            I => \N__55739\
        );

    \I__13764\ : Span4Mux_h
    port map (
            O => \N__55811\,
            I => \N__55736\
        );

    \I__13763\ : InMux
    port map (
            O => \N__55810\,
            I => \N__55733\
        );

    \I__13762\ : LocalMux
    port map (
            O => \N__55795\,
            I => \N__55730\
        );

    \I__13761\ : LocalMux
    port map (
            O => \N__55792\,
            I => \N__55725\
        );

    \I__13760\ : LocalMux
    port map (
            O => \N__55787\,
            I => \N__55725\
        );

    \I__13759\ : Span4Mux_h
    port map (
            O => \N__55782\,
            I => \N__55720\
        );

    \I__13758\ : Span4Mux_h
    port map (
            O => \N__55779\,
            I => \N__55720\
        );

    \I__13757\ : InMux
    port map (
            O => \N__55778\,
            I => \N__55717\
        );

    \I__13756\ : InMux
    port map (
            O => \N__55777\,
            I => \N__55714\
        );

    \I__13755\ : LocalMux
    port map (
            O => \N__55772\,
            I => \N__55709\
        );

    \I__13754\ : LocalMux
    port map (
            O => \N__55769\,
            I => \N__55709\
        );

    \I__13753\ : Span4Mux_v
    port map (
            O => \N__55766\,
            I => \N__55706\
        );

    \I__13752\ : InMux
    port map (
            O => \N__55765\,
            I => \N__55699\
        );

    \I__13751\ : InMux
    port map (
            O => \N__55764\,
            I => \N__55699\
        );

    \I__13750\ : InMux
    port map (
            O => \N__55763\,
            I => \N__55699\
        );

    \I__13749\ : LocalMux
    port map (
            O => \N__55760\,
            I => \N__55696\
        );

    \I__13748\ : InMux
    port map (
            O => \N__55759\,
            I => \N__55689\
        );

    \I__13747\ : InMux
    port map (
            O => \N__55758\,
            I => \N__55689\
        );

    \I__13746\ : InMux
    port map (
            O => \N__55757\,
            I => \N__55689\
        );

    \I__13745\ : Span4Mux_h
    port map (
            O => \N__55752\,
            I => \N__55680\
        );

    \I__13744\ : LocalMux
    port map (
            O => \N__55749\,
            I => \N__55680\
        );

    \I__13743\ : LocalMux
    port map (
            O => \N__55742\,
            I => \N__55680\
        );

    \I__13742\ : LocalMux
    port map (
            O => \N__55739\,
            I => \N__55680\
        );

    \I__13741\ : Span4Mux_v
    port map (
            O => \N__55736\,
            I => \N__55677\
        );

    \I__13740\ : LocalMux
    port map (
            O => \N__55733\,
            I => \N__55674\
        );

    \I__13739\ : Span4Mux_h
    port map (
            O => \N__55730\,
            I => \N__55667\
        );

    \I__13738\ : Span4Mux_h
    port map (
            O => \N__55725\,
            I => \N__55667\
        );

    \I__13737\ : Span4Mux_h
    port map (
            O => \N__55720\,
            I => \N__55667\
        );

    \I__13736\ : LocalMux
    port map (
            O => \N__55717\,
            I => \N__55656\
        );

    \I__13735\ : LocalMux
    port map (
            O => \N__55714\,
            I => \N__55656\
        );

    \I__13734\ : Span12Mux_v
    port map (
            O => \N__55709\,
            I => \N__55656\
        );

    \I__13733\ : Sp12to4
    port map (
            O => \N__55706\,
            I => \N__55656\
        );

    \I__13732\ : LocalMux
    port map (
            O => \N__55699\,
            I => \N__55656\
        );

    \I__13731\ : Span4Mux_v
    port map (
            O => \N__55696\,
            I => \N__55649\
        );

    \I__13730\ : LocalMux
    port map (
            O => \N__55689\,
            I => \N__55649\
        );

    \I__13729\ : Span4Mux_v
    port map (
            O => \N__55680\,
            I => \N__55649\
        );

    \I__13728\ : Odrv4
    port map (
            O => \N__55677\,
            I => comm_clear
        );

    \I__13727\ : Odrv4
    port map (
            O => \N__55674\,
            I => comm_clear
        );

    \I__13726\ : Odrv4
    port map (
            O => \N__55667\,
            I => comm_clear
        );

    \I__13725\ : Odrv12
    port map (
            O => \N__55656\,
            I => comm_clear
        );

    \I__13724\ : Odrv4
    port map (
            O => \N__55649\,
            I => comm_clear
        );

    \I__13723\ : InMux
    port map (
            O => \N__55638\,
            I => \N__55633\
        );

    \I__13722\ : InMux
    port map (
            O => \N__55637\,
            I => \N__55630\
        );

    \I__13721\ : InMux
    port map (
            O => \N__55636\,
            I => \N__55627\
        );

    \I__13720\ : LocalMux
    port map (
            O => \N__55633\,
            I => \N__55624\
        );

    \I__13719\ : LocalMux
    port map (
            O => \N__55630\,
            I => \N__55621\
        );

    \I__13718\ : LocalMux
    port map (
            O => \N__55627\,
            I => \N__55618\
        );

    \I__13717\ : Span4Mux_v
    port map (
            O => \N__55624\,
            I => \N__55615\
        );

    \I__13716\ : Span4Mux_h
    port map (
            O => \N__55621\,
            I => \N__55611\
        );

    \I__13715\ : Span4Mux_h
    port map (
            O => \N__55618\,
            I => \N__55608\
        );

    \I__13714\ : Span4Mux_h
    port map (
            O => \N__55615\,
            I => \N__55605\
        );

    \I__13713\ : InMux
    port map (
            O => \N__55614\,
            I => \N__55602\
        );

    \I__13712\ : Span4Mux_h
    port map (
            O => \N__55611\,
            I => \N__55598\
        );

    \I__13711\ : Span4Mux_v
    port map (
            O => \N__55608\,
            I => \N__55595\
        );

    \I__13710\ : Sp12to4
    port map (
            O => \N__55605\,
            I => \N__55590\
        );

    \I__13709\ : LocalMux
    port map (
            O => \N__55602\,
            I => \N__55590\
        );

    \I__13708\ : InMux
    port map (
            O => \N__55601\,
            I => \N__55587\
        );

    \I__13707\ : Sp12to4
    port map (
            O => \N__55598\,
            I => \N__55578\
        );

    \I__13706\ : Sp12to4
    port map (
            O => \N__55595\,
            I => \N__55578\
        );

    \I__13705\ : Span12Mux_s10_h
    port map (
            O => \N__55590\,
            I => \N__55578\
        );

    \I__13704\ : LocalMux
    port map (
            O => \N__55587\,
            I => \N__55578\
        );

    \I__13703\ : Span12Mux_v
    port map (
            O => \N__55578\,
            I => \N__55575\
        );

    \I__13702\ : Odrv12
    port map (
            O => \N__55575\,
            I => \ICE_SPI_MOSI\
        );

    \I__13701\ : SRMux
    port map (
            O => \N__55572\,
            I => \N__55569\
        );

    \I__13700\ : LocalMux
    port map (
            O => \N__55569\,
            I => \N__55566\
        );

    \I__13699\ : Span4Mux_h
    port map (
            O => \N__55566\,
            I => \N__55563\
        );

    \I__13698\ : Odrv4
    port map (
            O => \N__55563\,
            I => \comm_spi.imosi_N_752\
        );

    \I__13697\ : InMux
    port map (
            O => \N__55560\,
            I => \N__55557\
        );

    \I__13696\ : LocalMux
    port map (
            O => \N__55557\,
            I => \N__55553\
        );

    \I__13695\ : CascadeMux
    port map (
            O => \N__55556\,
            I => \N__55538\
        );

    \I__13694\ : Span4Mux_h
    port map (
            O => \N__55553\,
            I => \N__55535\
        );

    \I__13693\ : InMux
    port map (
            O => \N__55552\,
            I => \N__55526\
        );

    \I__13692\ : InMux
    port map (
            O => \N__55551\,
            I => \N__55526\
        );

    \I__13691\ : InMux
    port map (
            O => \N__55550\,
            I => \N__55526\
        );

    \I__13690\ : InMux
    port map (
            O => \N__55549\,
            I => \N__55526\
        );

    \I__13689\ : InMux
    port map (
            O => \N__55548\,
            I => \N__55519\
        );

    \I__13688\ : InMux
    port map (
            O => \N__55547\,
            I => \N__55507\
        );

    \I__13687\ : InMux
    port map (
            O => \N__55546\,
            I => \N__55504\
        );

    \I__13686\ : InMux
    port map (
            O => \N__55545\,
            I => \N__55501\
        );

    \I__13685\ : InMux
    port map (
            O => \N__55544\,
            I => \N__55492\
        );

    \I__13684\ : InMux
    port map (
            O => \N__55543\,
            I => \N__55492\
        );

    \I__13683\ : InMux
    port map (
            O => \N__55542\,
            I => \N__55492\
        );

    \I__13682\ : InMux
    port map (
            O => \N__55541\,
            I => \N__55489\
        );

    \I__13681\ : InMux
    port map (
            O => \N__55538\,
            I => \N__55486\
        );

    \I__13680\ : Span4Mux_h
    port map (
            O => \N__55535\,
            I => \N__55481\
        );

    \I__13679\ : LocalMux
    port map (
            O => \N__55526\,
            I => \N__55481\
        );

    \I__13678\ : InMux
    port map (
            O => \N__55525\,
            I => \N__55473\
        );

    \I__13677\ : InMux
    port map (
            O => \N__55524\,
            I => \N__55473\
        );

    \I__13676\ : InMux
    port map (
            O => \N__55523\,
            I => \N__55473\
        );

    \I__13675\ : InMux
    port map (
            O => \N__55522\,
            I => \N__55470\
        );

    \I__13674\ : LocalMux
    port map (
            O => \N__55519\,
            I => \N__55467\
        );

    \I__13673\ : InMux
    port map (
            O => \N__55518\,
            I => \N__55464\
        );

    \I__13672\ : InMux
    port map (
            O => \N__55517\,
            I => \N__55459\
        );

    \I__13671\ : InMux
    port map (
            O => \N__55516\,
            I => \N__55459\
        );

    \I__13670\ : InMux
    port map (
            O => \N__55515\,
            I => \N__55452\
        );

    \I__13669\ : InMux
    port map (
            O => \N__55514\,
            I => \N__55452\
        );

    \I__13668\ : InMux
    port map (
            O => \N__55513\,
            I => \N__55452\
        );

    \I__13667\ : CascadeMux
    port map (
            O => \N__55512\,
            I => \N__55448\
        );

    \I__13666\ : CascadeMux
    port map (
            O => \N__55511\,
            I => \N__55444\
        );

    \I__13665\ : CascadeMux
    port map (
            O => \N__55510\,
            I => \N__55441\
        );

    \I__13664\ : LocalMux
    port map (
            O => \N__55507\,
            I => \N__55434\
        );

    \I__13663\ : LocalMux
    port map (
            O => \N__55504\,
            I => \N__55434\
        );

    \I__13662\ : LocalMux
    port map (
            O => \N__55501\,
            I => \N__55434\
        );

    \I__13661\ : InMux
    port map (
            O => \N__55500\,
            I => \N__55431\
        );

    \I__13660\ : InMux
    port map (
            O => \N__55499\,
            I => \N__55426\
        );

    \I__13659\ : LocalMux
    port map (
            O => \N__55492\,
            I => \N__55423\
        );

    \I__13658\ : LocalMux
    port map (
            O => \N__55489\,
            I => \N__55418\
        );

    \I__13657\ : LocalMux
    port map (
            O => \N__55486\,
            I => \N__55415\
        );

    \I__13656\ : Span4Mux_v
    port map (
            O => \N__55481\,
            I => \N__55412\
        );

    \I__13655\ : InMux
    port map (
            O => \N__55480\,
            I => \N__55409\
        );

    \I__13654\ : LocalMux
    port map (
            O => \N__55473\,
            I => \N__55397\
        );

    \I__13653\ : LocalMux
    port map (
            O => \N__55470\,
            I => \N__55397\
        );

    \I__13652\ : Span4Mux_v
    port map (
            O => \N__55467\,
            I => \N__55397\
        );

    \I__13651\ : LocalMux
    port map (
            O => \N__55464\,
            I => \N__55394\
        );

    \I__13650\ : LocalMux
    port map (
            O => \N__55459\,
            I => \N__55391\
        );

    \I__13649\ : LocalMux
    port map (
            O => \N__55452\,
            I => \N__55388\
        );

    \I__13648\ : InMux
    port map (
            O => \N__55451\,
            I => \N__55385\
        );

    \I__13647\ : InMux
    port map (
            O => \N__55448\,
            I => \N__55380\
        );

    \I__13646\ : InMux
    port map (
            O => \N__55447\,
            I => \N__55380\
        );

    \I__13645\ : InMux
    port map (
            O => \N__55444\,
            I => \N__55375\
        );

    \I__13644\ : InMux
    port map (
            O => \N__55441\,
            I => \N__55375\
        );

    \I__13643\ : Span4Mux_v
    port map (
            O => \N__55434\,
            I => \N__55370\
        );

    \I__13642\ : LocalMux
    port map (
            O => \N__55431\,
            I => \N__55370\
        );

    \I__13641\ : InMux
    port map (
            O => \N__55430\,
            I => \N__55365\
        );

    \I__13640\ : InMux
    port map (
            O => \N__55429\,
            I => \N__55365\
        );

    \I__13639\ : LocalMux
    port map (
            O => \N__55426\,
            I => \N__55360\
        );

    \I__13638\ : Span4Mux_h
    port map (
            O => \N__55423\,
            I => \N__55360\
        );

    \I__13637\ : InMux
    port map (
            O => \N__55422\,
            I => \N__55357\
        );

    \I__13636\ : InMux
    port map (
            O => \N__55421\,
            I => \N__55354\
        );

    \I__13635\ : Span4Mux_v
    port map (
            O => \N__55418\,
            I => \N__55339\
        );

    \I__13634\ : Span4Mux_h
    port map (
            O => \N__55415\,
            I => \N__55339\
        );

    \I__13633\ : Span4Mux_h
    port map (
            O => \N__55412\,
            I => \N__55339\
        );

    \I__13632\ : LocalMux
    port map (
            O => \N__55409\,
            I => \N__55339\
        );

    \I__13631\ : InMux
    port map (
            O => \N__55408\,
            I => \N__55336\
        );

    \I__13630\ : InMux
    port map (
            O => \N__55407\,
            I => \N__55331\
        );

    \I__13629\ : InMux
    port map (
            O => \N__55406\,
            I => \N__55331\
        );

    \I__13628\ : InMux
    port map (
            O => \N__55405\,
            I => \N__55326\
        );

    \I__13627\ : InMux
    port map (
            O => \N__55404\,
            I => \N__55326\
        );

    \I__13626\ : Span4Mux_v
    port map (
            O => \N__55397\,
            I => \N__55317\
        );

    \I__13625\ : Span4Mux_v
    port map (
            O => \N__55394\,
            I => \N__55317\
        );

    \I__13624\ : Span4Mux_h
    port map (
            O => \N__55391\,
            I => \N__55317\
        );

    \I__13623\ : Span4Mux_v
    port map (
            O => \N__55388\,
            I => \N__55317\
        );

    \I__13622\ : LocalMux
    port map (
            O => \N__55385\,
            I => \N__55314\
        );

    \I__13621\ : LocalMux
    port map (
            O => \N__55380\,
            I => \N__55309\
        );

    \I__13620\ : LocalMux
    port map (
            O => \N__55375\,
            I => \N__55309\
        );

    \I__13619\ : Span4Mux_h
    port map (
            O => \N__55370\,
            I => \N__55302\
        );

    \I__13618\ : LocalMux
    port map (
            O => \N__55365\,
            I => \N__55302\
        );

    \I__13617\ : Span4Mux_v
    port map (
            O => \N__55360\,
            I => \N__55302\
        );

    \I__13616\ : LocalMux
    port map (
            O => \N__55357\,
            I => \N__55299\
        );

    \I__13615\ : LocalMux
    port map (
            O => \N__55354\,
            I => \N__55296\
        );

    \I__13614\ : InMux
    port map (
            O => \N__55353\,
            I => \N__55287\
        );

    \I__13613\ : InMux
    port map (
            O => \N__55352\,
            I => \N__55287\
        );

    \I__13612\ : InMux
    port map (
            O => \N__55351\,
            I => \N__55287\
        );

    \I__13611\ : InMux
    port map (
            O => \N__55350\,
            I => \N__55287\
        );

    \I__13610\ : InMux
    port map (
            O => \N__55349\,
            I => \N__55282\
        );

    \I__13609\ : InMux
    port map (
            O => \N__55348\,
            I => \N__55282\
        );

    \I__13608\ : Span4Mux_v
    port map (
            O => \N__55339\,
            I => \N__55277\
        );

    \I__13607\ : LocalMux
    port map (
            O => \N__55336\,
            I => \N__55277\
        );

    \I__13606\ : LocalMux
    port map (
            O => \N__55331\,
            I => \N__55270\
        );

    \I__13605\ : LocalMux
    port map (
            O => \N__55326\,
            I => \N__55270\
        );

    \I__13604\ : Sp12to4
    port map (
            O => \N__55317\,
            I => \N__55270\
        );

    \I__13603\ : Span4Mux_h
    port map (
            O => \N__55314\,
            I => \N__55263\
        );

    \I__13602\ : Span4Mux_v
    port map (
            O => \N__55309\,
            I => \N__55263\
        );

    \I__13601\ : Span4Mux_v
    port map (
            O => \N__55302\,
            I => \N__55263\
        );

    \I__13600\ : Odrv4
    port map (
            O => \N__55299\,
            I => comm_state_2
        );

    \I__13599\ : Odrv12
    port map (
            O => \N__55296\,
            I => comm_state_2
        );

    \I__13598\ : LocalMux
    port map (
            O => \N__55287\,
            I => comm_state_2
        );

    \I__13597\ : LocalMux
    port map (
            O => \N__55282\,
            I => comm_state_2
        );

    \I__13596\ : Odrv4
    port map (
            O => \N__55277\,
            I => comm_state_2
        );

    \I__13595\ : Odrv12
    port map (
            O => \N__55270\,
            I => comm_state_2
        );

    \I__13594\ : Odrv4
    port map (
            O => \N__55263\,
            I => comm_state_2
        );

    \I__13593\ : CascadeMux
    port map (
            O => \N__55248\,
            I => \N__55245\
        );

    \I__13592\ : InMux
    port map (
            O => \N__55245\,
            I => \N__55242\
        );

    \I__13591\ : LocalMux
    port map (
            O => \N__55242\,
            I => comm_length_0
        );

    \I__13590\ : CascadeMux
    port map (
            O => \N__55239\,
            I => \N__55236\
        );

    \I__13589\ : InMux
    port map (
            O => \N__55236\,
            I => \N__55225\
        );

    \I__13588\ : InMux
    port map (
            O => \N__55235\,
            I => \N__55225\
        );

    \I__13587\ : InMux
    port map (
            O => \N__55234\,
            I => \N__55220\
        );

    \I__13586\ : InMux
    port map (
            O => \N__55233\,
            I => \N__55220\
        );

    \I__13585\ : InMux
    port map (
            O => \N__55232\,
            I => \N__55205\
        );

    \I__13584\ : InMux
    port map (
            O => \N__55231\,
            I => \N__55200\
        );

    \I__13583\ : InMux
    port map (
            O => \N__55230\,
            I => \N__55200\
        );

    \I__13582\ : LocalMux
    port map (
            O => \N__55225\,
            I => \N__55195\
        );

    \I__13581\ : LocalMux
    port map (
            O => \N__55220\,
            I => \N__55195\
        );

    \I__13580\ : InMux
    port map (
            O => \N__55219\,
            I => \N__55190\
        );

    \I__13579\ : InMux
    port map (
            O => \N__55218\,
            I => \N__55190\
        );

    \I__13578\ : InMux
    port map (
            O => \N__55217\,
            I => \N__55184\
        );

    \I__13577\ : InMux
    port map (
            O => \N__55216\,
            I => \N__55177\
        );

    \I__13576\ : InMux
    port map (
            O => \N__55215\,
            I => \N__55177\
        );

    \I__13575\ : InMux
    port map (
            O => \N__55214\,
            I => \N__55177\
        );

    \I__13574\ : CascadeMux
    port map (
            O => \N__55213\,
            I => \N__55166\
        );

    \I__13573\ : CascadeMux
    port map (
            O => \N__55212\,
            I => \N__55142\
        );

    \I__13572\ : CascadeMux
    port map (
            O => \N__55211\,
            I => \N__55137\
        );

    \I__13571\ : CascadeMux
    port map (
            O => \N__55210\,
            I => \N__55133\
        );

    \I__13570\ : CascadeMux
    port map (
            O => \N__55209\,
            I => \N__55129\
        );

    \I__13569\ : InMux
    port map (
            O => \N__55208\,
            I => \N__55126\
        );

    \I__13568\ : LocalMux
    port map (
            O => \N__55205\,
            I => \N__55116\
        );

    \I__13567\ : LocalMux
    port map (
            O => \N__55200\,
            I => \N__55116\
        );

    \I__13566\ : Span4Mux_v
    port map (
            O => \N__55195\,
            I => \N__55116\
        );

    \I__13565\ : LocalMux
    port map (
            O => \N__55190\,
            I => \N__55116\
        );

    \I__13564\ : InMux
    port map (
            O => \N__55189\,
            I => \N__55109\
        );

    \I__13563\ : InMux
    port map (
            O => \N__55188\,
            I => \N__55109\
        );

    \I__13562\ : InMux
    port map (
            O => \N__55187\,
            I => \N__55109\
        );

    \I__13561\ : LocalMux
    port map (
            O => \N__55184\,
            I => \N__55104\
        );

    \I__13560\ : LocalMux
    port map (
            O => \N__55177\,
            I => \N__55104\
        );

    \I__13559\ : InMux
    port map (
            O => \N__55176\,
            I => \N__55101\
        );

    \I__13558\ : InMux
    port map (
            O => \N__55175\,
            I => \N__55098\
        );

    \I__13557\ : InMux
    port map (
            O => \N__55174\,
            I => \N__55095\
        );

    \I__13556\ : InMux
    port map (
            O => \N__55173\,
            I => \N__55092\
        );

    \I__13555\ : InMux
    port map (
            O => \N__55172\,
            I => \N__55085\
        );

    \I__13554\ : InMux
    port map (
            O => \N__55171\,
            I => \N__55085\
        );

    \I__13553\ : InMux
    port map (
            O => \N__55170\,
            I => \N__55085\
        );

    \I__13552\ : InMux
    port map (
            O => \N__55169\,
            I => \N__55082\
        );

    \I__13551\ : InMux
    port map (
            O => \N__55166\,
            I => \N__55071\
        );

    \I__13550\ : InMux
    port map (
            O => \N__55165\,
            I => \N__55071\
        );

    \I__13549\ : InMux
    port map (
            O => \N__55164\,
            I => \N__55071\
        );

    \I__13548\ : InMux
    port map (
            O => \N__55163\,
            I => \N__55071\
        );

    \I__13547\ : InMux
    port map (
            O => \N__55162\,
            I => \N__55071\
        );

    \I__13546\ : InMux
    port map (
            O => \N__55161\,
            I => \N__55066\
        );

    \I__13545\ : InMux
    port map (
            O => \N__55160\,
            I => \N__55066\
        );

    \I__13544\ : InMux
    port map (
            O => \N__55159\,
            I => \N__55063\
        );

    \I__13543\ : InMux
    port map (
            O => \N__55158\,
            I => \N__55060\
        );

    \I__13542\ : InMux
    port map (
            O => \N__55157\,
            I => \N__55053\
        );

    \I__13541\ : InMux
    port map (
            O => \N__55156\,
            I => \N__55050\
        );

    \I__13540\ : InMux
    port map (
            O => \N__55155\,
            I => \N__55047\
        );

    \I__13539\ : InMux
    port map (
            O => \N__55154\,
            I => \N__55042\
        );

    \I__13538\ : InMux
    port map (
            O => \N__55153\,
            I => \N__55042\
        );

    \I__13537\ : InMux
    port map (
            O => \N__55152\,
            I => \N__55037\
        );

    \I__13536\ : InMux
    port map (
            O => \N__55151\,
            I => \N__55037\
        );

    \I__13535\ : InMux
    port map (
            O => \N__55150\,
            I => \N__55029\
        );

    \I__13534\ : InMux
    port map (
            O => \N__55149\,
            I => \N__55029\
        );

    \I__13533\ : InMux
    port map (
            O => \N__55148\,
            I => \N__55026\
        );

    \I__13532\ : CascadeMux
    port map (
            O => \N__55147\,
            I => \N__55023\
        );

    \I__13531\ : CascadeMux
    port map (
            O => \N__55146\,
            I => \N__55019\
        );

    \I__13530\ : InMux
    port map (
            O => \N__55145\,
            I => \N__55012\
        );

    \I__13529\ : InMux
    port map (
            O => \N__55142\,
            I => \N__55012\
        );

    \I__13528\ : InMux
    port map (
            O => \N__55141\,
            I => \N__55012\
        );

    \I__13527\ : InMux
    port map (
            O => \N__55140\,
            I => \N__55009\
        );

    \I__13526\ : InMux
    port map (
            O => \N__55137\,
            I => \N__55006\
        );

    \I__13525\ : InMux
    port map (
            O => \N__55136\,
            I => \N__55003\
        );

    \I__13524\ : InMux
    port map (
            O => \N__55133\,
            I => \N__54996\
        );

    \I__13523\ : InMux
    port map (
            O => \N__55132\,
            I => \N__54996\
        );

    \I__13522\ : InMux
    port map (
            O => \N__55129\,
            I => \N__54996\
        );

    \I__13521\ : LocalMux
    port map (
            O => \N__55126\,
            I => \N__54993\
        );

    \I__13520\ : InMux
    port map (
            O => \N__55125\,
            I => \N__54990\
        );

    \I__13519\ : Span4Mux_v
    port map (
            O => \N__55116\,
            I => \N__54985\
        );

    \I__13518\ : LocalMux
    port map (
            O => \N__55109\,
            I => \N__54985\
        );

    \I__13517\ : Span4Mux_v
    port map (
            O => \N__55104\,
            I => \N__54980\
        );

    \I__13516\ : LocalMux
    port map (
            O => \N__55101\,
            I => \N__54980\
        );

    \I__13515\ : LocalMux
    port map (
            O => \N__55098\,
            I => \N__54975\
        );

    \I__13514\ : LocalMux
    port map (
            O => \N__55095\,
            I => \N__54968\
        );

    \I__13513\ : LocalMux
    port map (
            O => \N__55092\,
            I => \N__54968\
        );

    \I__13512\ : LocalMux
    port map (
            O => \N__55085\,
            I => \N__54968\
        );

    \I__13511\ : LocalMux
    port map (
            O => \N__55082\,
            I => \N__54965\
        );

    \I__13510\ : LocalMux
    port map (
            O => \N__55071\,
            I => \N__54962\
        );

    \I__13509\ : LocalMux
    port map (
            O => \N__55066\,
            I => \N__54959\
        );

    \I__13508\ : LocalMux
    port map (
            O => \N__55063\,
            I => \N__54956\
        );

    \I__13507\ : LocalMux
    port map (
            O => \N__55060\,
            I => \N__54953\
        );

    \I__13506\ : InMux
    port map (
            O => \N__55059\,
            I => \N__54950\
        );

    \I__13505\ : InMux
    port map (
            O => \N__55058\,
            I => \N__54947\
        );

    \I__13504\ : InMux
    port map (
            O => \N__55057\,
            I => \N__54944\
        );

    \I__13503\ : InMux
    port map (
            O => \N__55056\,
            I => \N__54941\
        );

    \I__13502\ : LocalMux
    port map (
            O => \N__55053\,
            I => \N__54930\
        );

    \I__13501\ : LocalMux
    port map (
            O => \N__55050\,
            I => \N__54930\
        );

    \I__13500\ : LocalMux
    port map (
            O => \N__55047\,
            I => \N__54930\
        );

    \I__13499\ : LocalMux
    port map (
            O => \N__55042\,
            I => \N__54930\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__55037\,
            I => \N__54930\
        );

    \I__13497\ : InMux
    port map (
            O => \N__55036\,
            I => \N__54925\
        );

    \I__13496\ : InMux
    port map (
            O => \N__55035\,
            I => \N__54925\
        );

    \I__13495\ : InMux
    port map (
            O => \N__55034\,
            I => \N__54922\
        );

    \I__13494\ : LocalMux
    port map (
            O => \N__55029\,
            I => \N__54917\
        );

    \I__13493\ : LocalMux
    port map (
            O => \N__55026\,
            I => \N__54917\
        );

    \I__13492\ : InMux
    port map (
            O => \N__55023\,
            I => \N__54914\
        );

    \I__13491\ : InMux
    port map (
            O => \N__55022\,
            I => \N__54910\
        );

    \I__13490\ : InMux
    port map (
            O => \N__55019\,
            I => \N__54907\
        );

    \I__13489\ : LocalMux
    port map (
            O => \N__55012\,
            I => \N__54904\
        );

    \I__13488\ : LocalMux
    port map (
            O => \N__55009\,
            I => \N__54895\
        );

    \I__13487\ : LocalMux
    port map (
            O => \N__55006\,
            I => \N__54895\
        );

    \I__13486\ : LocalMux
    port map (
            O => \N__55003\,
            I => \N__54895\
        );

    \I__13485\ : LocalMux
    port map (
            O => \N__54996\,
            I => \N__54895\
        );

    \I__13484\ : Span4Mux_v
    port map (
            O => \N__54993\,
            I => \N__54892\
        );

    \I__13483\ : LocalMux
    port map (
            O => \N__54990\,
            I => \N__54885\
        );

    \I__13482\ : Span4Mux_h
    port map (
            O => \N__54985\,
            I => \N__54885\
        );

    \I__13481\ : Span4Mux_v
    port map (
            O => \N__54980\,
            I => \N__54885\
        );

    \I__13480\ : InMux
    port map (
            O => \N__54979\,
            I => \N__54879\
        );

    \I__13479\ : InMux
    port map (
            O => \N__54978\,
            I => \N__54879\
        );

    \I__13478\ : Span4Mux_v
    port map (
            O => \N__54975\,
            I => \N__54874\
        );

    \I__13477\ : Span4Mux_v
    port map (
            O => \N__54968\,
            I => \N__54874\
        );

    \I__13476\ : Span4Mux_v
    port map (
            O => \N__54965\,
            I => \N__54869\
        );

    \I__13475\ : Span4Mux_v
    port map (
            O => \N__54962\,
            I => \N__54869\
        );

    \I__13474\ : Span4Mux_v
    port map (
            O => \N__54959\,
            I => \N__54865\
        );

    \I__13473\ : Span4Mux_v
    port map (
            O => \N__54956\,
            I => \N__54860\
        );

    \I__13472\ : Span4Mux_v
    port map (
            O => \N__54953\,
            I => \N__54860\
        );

    \I__13471\ : LocalMux
    port map (
            O => \N__54950\,
            I => \N__54857\
        );

    \I__13470\ : LocalMux
    port map (
            O => \N__54947\,
            I => \N__54852\
        );

    \I__13469\ : LocalMux
    port map (
            O => \N__54944\,
            I => \N__54852\
        );

    \I__13468\ : LocalMux
    port map (
            O => \N__54941\,
            I => \N__54849\
        );

    \I__13467\ : Span4Mux_v
    port map (
            O => \N__54930\,
            I => \N__54838\
        );

    \I__13466\ : LocalMux
    port map (
            O => \N__54925\,
            I => \N__54838\
        );

    \I__13465\ : LocalMux
    port map (
            O => \N__54922\,
            I => \N__54838\
        );

    \I__13464\ : Span4Mux_h
    port map (
            O => \N__54917\,
            I => \N__54838\
        );

    \I__13463\ : LocalMux
    port map (
            O => \N__54914\,
            I => \N__54838\
        );

    \I__13462\ : InMux
    port map (
            O => \N__54913\,
            I => \N__54832\
        );

    \I__13461\ : LocalMux
    port map (
            O => \N__54910\,
            I => \N__54827\
        );

    \I__13460\ : LocalMux
    port map (
            O => \N__54907\,
            I => \N__54827\
        );

    \I__13459\ : Span4Mux_h
    port map (
            O => \N__54904\,
            I => \N__54818\
        );

    \I__13458\ : Span4Mux_v
    port map (
            O => \N__54895\,
            I => \N__54818\
        );

    \I__13457\ : Span4Mux_v
    port map (
            O => \N__54892\,
            I => \N__54818\
        );

    \I__13456\ : Span4Mux_v
    port map (
            O => \N__54885\,
            I => \N__54818\
        );

    \I__13455\ : InMux
    port map (
            O => \N__54884\,
            I => \N__54815\
        );

    \I__13454\ : LocalMux
    port map (
            O => \N__54879\,
            I => \N__54808\
        );

    \I__13453\ : Span4Mux_h
    port map (
            O => \N__54874\,
            I => \N__54808\
        );

    \I__13452\ : Span4Mux_h
    port map (
            O => \N__54869\,
            I => \N__54808\
        );

    \I__13451\ : InMux
    port map (
            O => \N__54868\,
            I => \N__54805\
        );

    \I__13450\ : Span4Mux_h
    port map (
            O => \N__54865\,
            I => \N__54800\
        );

    \I__13449\ : Span4Mux_h
    port map (
            O => \N__54860\,
            I => \N__54800\
        );

    \I__13448\ : Span4Mux_h
    port map (
            O => \N__54857\,
            I => \N__54791\
        );

    \I__13447\ : Span4Mux_h
    port map (
            O => \N__54852\,
            I => \N__54791\
        );

    \I__13446\ : Span4Mux_v
    port map (
            O => \N__54849\,
            I => \N__54791\
        );

    \I__13445\ : Span4Mux_h
    port map (
            O => \N__54838\,
            I => \N__54791\
        );

    \I__13444\ : InMux
    port map (
            O => \N__54837\,
            I => \N__54784\
        );

    \I__13443\ : InMux
    port map (
            O => \N__54836\,
            I => \N__54784\
        );

    \I__13442\ : InMux
    port map (
            O => \N__54835\,
            I => \N__54784\
        );

    \I__13441\ : LocalMux
    port map (
            O => \N__54832\,
            I => comm_cmd_1
        );

    \I__13440\ : Odrv12
    port map (
            O => \N__54827\,
            I => comm_cmd_1
        );

    \I__13439\ : Odrv4
    port map (
            O => \N__54818\,
            I => comm_cmd_1
        );

    \I__13438\ : LocalMux
    port map (
            O => \N__54815\,
            I => comm_cmd_1
        );

    \I__13437\ : Odrv4
    port map (
            O => \N__54808\,
            I => comm_cmd_1
        );

    \I__13436\ : LocalMux
    port map (
            O => \N__54805\,
            I => comm_cmd_1
        );

    \I__13435\ : Odrv4
    port map (
            O => \N__54800\,
            I => comm_cmd_1
        );

    \I__13434\ : Odrv4
    port map (
            O => \N__54791\,
            I => comm_cmd_1
        );

    \I__13433\ : LocalMux
    port map (
            O => \N__54784\,
            I => comm_cmd_1
        );

    \I__13432\ : InMux
    port map (
            O => \N__54765\,
            I => \N__54750\
        );

    \I__13431\ : InMux
    port map (
            O => \N__54764\,
            I => \N__54741\
        );

    \I__13430\ : InMux
    port map (
            O => \N__54763\,
            I => \N__54738\
        );

    \I__13429\ : InMux
    port map (
            O => \N__54762\,
            I => \N__54733\
        );

    \I__13428\ : InMux
    port map (
            O => \N__54761\,
            I => \N__54733\
        );

    \I__13427\ : InMux
    port map (
            O => \N__54760\,
            I => \N__54728\
        );

    \I__13426\ : InMux
    port map (
            O => \N__54759\,
            I => \N__54728\
        );

    \I__13425\ : InMux
    port map (
            O => \N__54758\,
            I => \N__54723\
        );

    \I__13424\ : InMux
    port map (
            O => \N__54757\,
            I => \N__54723\
        );

    \I__13423\ : InMux
    port map (
            O => \N__54756\,
            I => \N__54720\
        );

    \I__13422\ : InMux
    port map (
            O => \N__54755\,
            I => \N__54716\
        );

    \I__13421\ : InMux
    port map (
            O => \N__54754\,
            I => \N__54713\
        );

    \I__13420\ : InMux
    port map (
            O => \N__54753\,
            I => \N__54708\
        );

    \I__13419\ : LocalMux
    port map (
            O => \N__54750\,
            I => \N__54703\
        );

    \I__13418\ : InMux
    port map (
            O => \N__54749\,
            I => \N__54698\
        );

    \I__13417\ : InMux
    port map (
            O => \N__54748\,
            I => \N__54698\
        );

    \I__13416\ : InMux
    port map (
            O => \N__54747\,
            I => \N__54688\
        );

    \I__13415\ : InMux
    port map (
            O => \N__54746\,
            I => \N__54683\
        );

    \I__13414\ : InMux
    port map (
            O => \N__54745\,
            I => \N__54680\
        );

    \I__13413\ : InMux
    port map (
            O => \N__54744\,
            I => \N__54677\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__54741\,
            I => \N__54672\
        );

    \I__13411\ : LocalMux
    port map (
            O => \N__54738\,
            I => \N__54672\
        );

    \I__13410\ : LocalMux
    port map (
            O => \N__54733\,
            I => \N__54665\
        );

    \I__13409\ : LocalMux
    port map (
            O => \N__54728\,
            I => \N__54665\
        );

    \I__13408\ : LocalMux
    port map (
            O => \N__54723\,
            I => \N__54665\
        );

    \I__13407\ : LocalMux
    port map (
            O => \N__54720\,
            I => \N__54662\
        );

    \I__13406\ : InMux
    port map (
            O => \N__54719\,
            I => \N__54659\
        );

    \I__13405\ : LocalMux
    port map (
            O => \N__54716\,
            I => \N__54654\
        );

    \I__13404\ : LocalMux
    port map (
            O => \N__54713\,
            I => \N__54654\
        );

    \I__13403\ : InMux
    port map (
            O => \N__54712\,
            I => \N__54648\
        );

    \I__13402\ : InMux
    port map (
            O => \N__54711\,
            I => \N__54648\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__54708\,
            I => \N__54645\
        );

    \I__13400\ : InMux
    port map (
            O => \N__54707\,
            I => \N__54641\
        );

    \I__13399\ : InMux
    port map (
            O => \N__54706\,
            I => \N__54638\
        );

    \I__13398\ : Span4Mux_h
    port map (
            O => \N__54703\,
            I => \N__54635\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__54698\,
            I => \N__54632\
        );

    \I__13396\ : InMux
    port map (
            O => \N__54697\,
            I => \N__54628\
        );

    \I__13395\ : InMux
    port map (
            O => \N__54696\,
            I => \N__54625\
        );

    \I__13394\ : InMux
    port map (
            O => \N__54695\,
            I => \N__54622\
        );

    \I__13393\ : InMux
    port map (
            O => \N__54694\,
            I => \N__54619\
        );

    \I__13392\ : InMux
    port map (
            O => \N__54693\,
            I => \N__54614\
        );

    \I__13391\ : InMux
    port map (
            O => \N__54692\,
            I => \N__54614\
        );

    \I__13390\ : InMux
    port map (
            O => \N__54691\,
            I => \N__54611\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__54688\,
            I => \N__54608\
        );

    \I__13388\ : InMux
    port map (
            O => \N__54687\,
            I => \N__54603\
        );

    \I__13387\ : InMux
    port map (
            O => \N__54686\,
            I => \N__54603\
        );

    \I__13386\ : LocalMux
    port map (
            O => \N__54683\,
            I => \N__54598\
        );

    \I__13385\ : LocalMux
    port map (
            O => \N__54680\,
            I => \N__54595\
        );

    \I__13384\ : LocalMux
    port map (
            O => \N__54677\,
            I => \N__54588\
        );

    \I__13383\ : Span4Mux_v
    port map (
            O => \N__54672\,
            I => \N__54588\
        );

    \I__13382\ : Span4Mux_v
    port map (
            O => \N__54665\,
            I => \N__54588\
        );

    \I__13381\ : Span4Mux_v
    port map (
            O => \N__54662\,
            I => \N__54585\
        );

    \I__13380\ : LocalMux
    port map (
            O => \N__54659\,
            I => \N__54582\
        );

    \I__13379\ : Span4Mux_h
    port map (
            O => \N__54654\,
            I => \N__54579\
        );

    \I__13378\ : InMux
    port map (
            O => \N__54653\,
            I => \N__54576\
        );

    \I__13377\ : LocalMux
    port map (
            O => \N__54648\,
            I => \N__54573\
        );

    \I__13376\ : Sp12to4
    port map (
            O => \N__54645\,
            I => \N__54570\
        );

    \I__13375\ : InMux
    port map (
            O => \N__54644\,
            I => \N__54566\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__54641\,
            I => \N__54563\
        );

    \I__13373\ : LocalMux
    port map (
            O => \N__54638\,
            I => \N__54558\
        );

    \I__13372\ : Span4Mux_v
    port map (
            O => \N__54635\,
            I => \N__54558\
        );

    \I__13371\ : Span4Mux_h
    port map (
            O => \N__54632\,
            I => \N__54555\
        );

    \I__13370\ : InMux
    port map (
            O => \N__54631\,
            I => \N__54551\
        );

    \I__13369\ : LocalMux
    port map (
            O => \N__54628\,
            I => \N__54546\
        );

    \I__13368\ : LocalMux
    port map (
            O => \N__54625\,
            I => \N__54546\
        );

    \I__13367\ : LocalMux
    port map (
            O => \N__54622\,
            I => \N__54539\
        );

    \I__13366\ : LocalMux
    port map (
            O => \N__54619\,
            I => \N__54539\
        );

    \I__13365\ : LocalMux
    port map (
            O => \N__54614\,
            I => \N__54539\
        );

    \I__13364\ : LocalMux
    port map (
            O => \N__54611\,
            I => \N__54532\
        );

    \I__13363\ : Span4Mux_h
    port map (
            O => \N__54608\,
            I => \N__54532\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__54603\,
            I => \N__54532\
        );

    \I__13361\ : InMux
    port map (
            O => \N__54602\,
            I => \N__54529\
        );

    \I__13360\ : InMux
    port map (
            O => \N__54601\,
            I => \N__54526\
        );

    \I__13359\ : Span4Mux_h
    port map (
            O => \N__54598\,
            I => \N__54517\
        );

    \I__13358\ : Span4Mux_v
    port map (
            O => \N__54595\,
            I => \N__54517\
        );

    \I__13357\ : Span4Mux_h
    port map (
            O => \N__54588\,
            I => \N__54517\
        );

    \I__13356\ : Span4Mux_v
    port map (
            O => \N__54585\,
            I => \N__54517\
        );

    \I__13355\ : Span4Mux_h
    port map (
            O => \N__54582\,
            I => \N__54512\
        );

    \I__13354\ : Span4Mux_v
    port map (
            O => \N__54579\,
            I => \N__54512\
        );

    \I__13353\ : LocalMux
    port map (
            O => \N__54576\,
            I => \N__54505\
        );

    \I__13352\ : Span12Mux_v
    port map (
            O => \N__54573\,
            I => \N__54505\
        );

    \I__13351\ : Span12Mux_v
    port map (
            O => \N__54570\,
            I => \N__54505\
        );

    \I__13350\ : InMux
    port map (
            O => \N__54569\,
            I => \N__54502\
        );

    \I__13349\ : LocalMux
    port map (
            O => \N__54566\,
            I => \N__54493\
        );

    \I__13348\ : Span4Mux_v
    port map (
            O => \N__54563\,
            I => \N__54493\
        );

    \I__13347\ : Span4Mux_h
    port map (
            O => \N__54558\,
            I => \N__54493\
        );

    \I__13346\ : Span4Mux_h
    port map (
            O => \N__54555\,
            I => \N__54493\
        );

    \I__13345\ : InMux
    port map (
            O => \N__54554\,
            I => \N__54490\
        );

    \I__13344\ : LocalMux
    port map (
            O => \N__54551\,
            I => \N__54481\
        );

    \I__13343\ : Span4Mux_v
    port map (
            O => \N__54546\,
            I => \N__54481\
        );

    \I__13342\ : Span4Mux_v
    port map (
            O => \N__54539\,
            I => \N__54481\
        );

    \I__13341\ : Span4Mux_v
    port map (
            O => \N__54532\,
            I => \N__54481\
        );

    \I__13340\ : LocalMux
    port map (
            O => \N__54529\,
            I => \N__54478\
        );

    \I__13339\ : LocalMux
    port map (
            O => \N__54526\,
            I => comm_cmd_3
        );

    \I__13338\ : Odrv4
    port map (
            O => \N__54517\,
            I => comm_cmd_3
        );

    \I__13337\ : Odrv4
    port map (
            O => \N__54512\,
            I => comm_cmd_3
        );

    \I__13336\ : Odrv12
    port map (
            O => \N__54505\,
            I => comm_cmd_3
        );

    \I__13335\ : LocalMux
    port map (
            O => \N__54502\,
            I => comm_cmd_3
        );

    \I__13334\ : Odrv4
    port map (
            O => \N__54493\,
            I => comm_cmd_3
        );

    \I__13333\ : LocalMux
    port map (
            O => \N__54490\,
            I => comm_cmd_3
        );

    \I__13332\ : Odrv4
    port map (
            O => \N__54481\,
            I => comm_cmd_3
        );

    \I__13331\ : Odrv12
    port map (
            O => \N__54478\,
            I => comm_cmd_3
        );

    \I__13330\ : CascadeMux
    port map (
            O => \N__54459\,
            I => \N__54456\
        );

    \I__13329\ : InMux
    port map (
            O => \N__54456\,
            I => \N__54453\
        );

    \I__13328\ : LocalMux
    port map (
            O => \N__54453\,
            I => \N__54450\
        );

    \I__13327\ : Span4Mux_h
    port map (
            O => \N__54450\,
            I => \N__54446\
        );

    \I__13326\ : InMux
    port map (
            O => \N__54449\,
            I => \N__54443\
        );

    \I__13325\ : Odrv4
    port map (
            O => \N__54446\,
            I => comm_length_1
        );

    \I__13324\ : LocalMux
    port map (
            O => \N__54443\,
            I => comm_length_1
        );

    \I__13323\ : ClkMux
    port map (
            O => \N__54438\,
            I => \N__53928\
        );

    \I__13322\ : ClkMux
    port map (
            O => \N__54437\,
            I => \N__53928\
        );

    \I__13321\ : ClkMux
    port map (
            O => \N__54436\,
            I => \N__53928\
        );

    \I__13320\ : ClkMux
    port map (
            O => \N__54435\,
            I => \N__53928\
        );

    \I__13319\ : ClkMux
    port map (
            O => \N__54434\,
            I => \N__53928\
        );

    \I__13318\ : ClkMux
    port map (
            O => \N__54433\,
            I => \N__53928\
        );

    \I__13317\ : ClkMux
    port map (
            O => \N__54432\,
            I => \N__53928\
        );

    \I__13316\ : ClkMux
    port map (
            O => \N__54431\,
            I => \N__53928\
        );

    \I__13315\ : ClkMux
    port map (
            O => \N__54430\,
            I => \N__53928\
        );

    \I__13314\ : ClkMux
    port map (
            O => \N__54429\,
            I => \N__53928\
        );

    \I__13313\ : ClkMux
    port map (
            O => \N__54428\,
            I => \N__53928\
        );

    \I__13312\ : ClkMux
    port map (
            O => \N__54427\,
            I => \N__53928\
        );

    \I__13311\ : ClkMux
    port map (
            O => \N__54426\,
            I => \N__53928\
        );

    \I__13310\ : ClkMux
    port map (
            O => \N__54425\,
            I => \N__53928\
        );

    \I__13309\ : ClkMux
    port map (
            O => \N__54424\,
            I => \N__53928\
        );

    \I__13308\ : ClkMux
    port map (
            O => \N__54423\,
            I => \N__53928\
        );

    \I__13307\ : ClkMux
    port map (
            O => \N__54422\,
            I => \N__53928\
        );

    \I__13306\ : ClkMux
    port map (
            O => \N__54421\,
            I => \N__53928\
        );

    \I__13305\ : ClkMux
    port map (
            O => \N__54420\,
            I => \N__53928\
        );

    \I__13304\ : ClkMux
    port map (
            O => \N__54419\,
            I => \N__53928\
        );

    \I__13303\ : ClkMux
    port map (
            O => \N__54418\,
            I => \N__53928\
        );

    \I__13302\ : ClkMux
    port map (
            O => \N__54417\,
            I => \N__53928\
        );

    \I__13301\ : ClkMux
    port map (
            O => \N__54416\,
            I => \N__53928\
        );

    \I__13300\ : ClkMux
    port map (
            O => \N__54415\,
            I => \N__53928\
        );

    \I__13299\ : ClkMux
    port map (
            O => \N__54414\,
            I => \N__53928\
        );

    \I__13298\ : ClkMux
    port map (
            O => \N__54413\,
            I => \N__53928\
        );

    \I__13297\ : ClkMux
    port map (
            O => \N__54412\,
            I => \N__53928\
        );

    \I__13296\ : ClkMux
    port map (
            O => \N__54411\,
            I => \N__53928\
        );

    \I__13295\ : ClkMux
    port map (
            O => \N__54410\,
            I => \N__53928\
        );

    \I__13294\ : ClkMux
    port map (
            O => \N__54409\,
            I => \N__53928\
        );

    \I__13293\ : ClkMux
    port map (
            O => \N__54408\,
            I => \N__53928\
        );

    \I__13292\ : ClkMux
    port map (
            O => \N__54407\,
            I => \N__53928\
        );

    \I__13291\ : ClkMux
    port map (
            O => \N__54406\,
            I => \N__53928\
        );

    \I__13290\ : ClkMux
    port map (
            O => \N__54405\,
            I => \N__53928\
        );

    \I__13289\ : ClkMux
    port map (
            O => \N__54404\,
            I => \N__53928\
        );

    \I__13288\ : ClkMux
    port map (
            O => \N__54403\,
            I => \N__53928\
        );

    \I__13287\ : ClkMux
    port map (
            O => \N__54402\,
            I => \N__53928\
        );

    \I__13286\ : ClkMux
    port map (
            O => \N__54401\,
            I => \N__53928\
        );

    \I__13285\ : ClkMux
    port map (
            O => \N__54400\,
            I => \N__53928\
        );

    \I__13284\ : ClkMux
    port map (
            O => \N__54399\,
            I => \N__53928\
        );

    \I__13283\ : ClkMux
    port map (
            O => \N__54398\,
            I => \N__53928\
        );

    \I__13282\ : ClkMux
    port map (
            O => \N__54397\,
            I => \N__53928\
        );

    \I__13281\ : ClkMux
    port map (
            O => \N__54396\,
            I => \N__53928\
        );

    \I__13280\ : ClkMux
    port map (
            O => \N__54395\,
            I => \N__53928\
        );

    \I__13279\ : ClkMux
    port map (
            O => \N__54394\,
            I => \N__53928\
        );

    \I__13278\ : ClkMux
    port map (
            O => \N__54393\,
            I => \N__53928\
        );

    \I__13277\ : ClkMux
    port map (
            O => \N__54392\,
            I => \N__53928\
        );

    \I__13276\ : ClkMux
    port map (
            O => \N__54391\,
            I => \N__53928\
        );

    \I__13275\ : ClkMux
    port map (
            O => \N__54390\,
            I => \N__53928\
        );

    \I__13274\ : ClkMux
    port map (
            O => \N__54389\,
            I => \N__53928\
        );

    \I__13273\ : ClkMux
    port map (
            O => \N__54388\,
            I => \N__53928\
        );

    \I__13272\ : ClkMux
    port map (
            O => \N__54387\,
            I => \N__53928\
        );

    \I__13271\ : ClkMux
    port map (
            O => \N__54386\,
            I => \N__53928\
        );

    \I__13270\ : ClkMux
    port map (
            O => \N__54385\,
            I => \N__53928\
        );

    \I__13269\ : ClkMux
    port map (
            O => \N__54384\,
            I => \N__53928\
        );

    \I__13268\ : ClkMux
    port map (
            O => \N__54383\,
            I => \N__53928\
        );

    \I__13267\ : ClkMux
    port map (
            O => \N__54382\,
            I => \N__53928\
        );

    \I__13266\ : ClkMux
    port map (
            O => \N__54381\,
            I => \N__53928\
        );

    \I__13265\ : ClkMux
    port map (
            O => \N__54380\,
            I => \N__53928\
        );

    \I__13264\ : ClkMux
    port map (
            O => \N__54379\,
            I => \N__53928\
        );

    \I__13263\ : ClkMux
    port map (
            O => \N__54378\,
            I => \N__53928\
        );

    \I__13262\ : ClkMux
    port map (
            O => \N__54377\,
            I => \N__53928\
        );

    \I__13261\ : ClkMux
    port map (
            O => \N__54376\,
            I => \N__53928\
        );

    \I__13260\ : ClkMux
    port map (
            O => \N__54375\,
            I => \N__53928\
        );

    \I__13259\ : ClkMux
    port map (
            O => \N__54374\,
            I => \N__53928\
        );

    \I__13258\ : ClkMux
    port map (
            O => \N__54373\,
            I => \N__53928\
        );

    \I__13257\ : ClkMux
    port map (
            O => \N__54372\,
            I => \N__53928\
        );

    \I__13256\ : ClkMux
    port map (
            O => \N__54371\,
            I => \N__53928\
        );

    \I__13255\ : ClkMux
    port map (
            O => \N__54370\,
            I => \N__53928\
        );

    \I__13254\ : ClkMux
    port map (
            O => \N__54369\,
            I => \N__53928\
        );

    \I__13253\ : ClkMux
    port map (
            O => \N__54368\,
            I => \N__53928\
        );

    \I__13252\ : ClkMux
    port map (
            O => \N__54367\,
            I => \N__53928\
        );

    \I__13251\ : ClkMux
    port map (
            O => \N__54366\,
            I => \N__53928\
        );

    \I__13250\ : ClkMux
    port map (
            O => \N__54365\,
            I => \N__53928\
        );

    \I__13249\ : ClkMux
    port map (
            O => \N__54364\,
            I => \N__53928\
        );

    \I__13248\ : ClkMux
    port map (
            O => \N__54363\,
            I => \N__53928\
        );

    \I__13247\ : ClkMux
    port map (
            O => \N__54362\,
            I => \N__53928\
        );

    \I__13246\ : ClkMux
    port map (
            O => \N__54361\,
            I => \N__53928\
        );

    \I__13245\ : ClkMux
    port map (
            O => \N__54360\,
            I => \N__53928\
        );

    \I__13244\ : ClkMux
    port map (
            O => \N__54359\,
            I => \N__53928\
        );

    \I__13243\ : ClkMux
    port map (
            O => \N__54358\,
            I => \N__53928\
        );

    \I__13242\ : ClkMux
    port map (
            O => \N__54357\,
            I => \N__53928\
        );

    \I__13241\ : ClkMux
    port map (
            O => \N__54356\,
            I => \N__53928\
        );

    \I__13240\ : ClkMux
    port map (
            O => \N__54355\,
            I => \N__53928\
        );

    \I__13239\ : ClkMux
    port map (
            O => \N__54354\,
            I => \N__53928\
        );

    \I__13238\ : ClkMux
    port map (
            O => \N__54353\,
            I => \N__53928\
        );

    \I__13237\ : ClkMux
    port map (
            O => \N__54352\,
            I => \N__53928\
        );

    \I__13236\ : ClkMux
    port map (
            O => \N__54351\,
            I => \N__53928\
        );

    \I__13235\ : ClkMux
    port map (
            O => \N__54350\,
            I => \N__53928\
        );

    \I__13234\ : ClkMux
    port map (
            O => \N__54349\,
            I => \N__53928\
        );

    \I__13233\ : ClkMux
    port map (
            O => \N__54348\,
            I => \N__53928\
        );

    \I__13232\ : ClkMux
    port map (
            O => \N__54347\,
            I => \N__53928\
        );

    \I__13231\ : ClkMux
    port map (
            O => \N__54346\,
            I => \N__53928\
        );

    \I__13230\ : ClkMux
    port map (
            O => \N__54345\,
            I => \N__53928\
        );

    \I__13229\ : ClkMux
    port map (
            O => \N__54344\,
            I => \N__53928\
        );

    \I__13228\ : ClkMux
    port map (
            O => \N__54343\,
            I => \N__53928\
        );

    \I__13227\ : ClkMux
    port map (
            O => \N__54342\,
            I => \N__53928\
        );

    \I__13226\ : ClkMux
    port map (
            O => \N__54341\,
            I => \N__53928\
        );

    \I__13225\ : ClkMux
    port map (
            O => \N__54340\,
            I => \N__53928\
        );

    \I__13224\ : ClkMux
    port map (
            O => \N__54339\,
            I => \N__53928\
        );

    \I__13223\ : ClkMux
    port map (
            O => \N__54338\,
            I => \N__53928\
        );

    \I__13222\ : ClkMux
    port map (
            O => \N__54337\,
            I => \N__53928\
        );

    \I__13221\ : ClkMux
    port map (
            O => \N__54336\,
            I => \N__53928\
        );

    \I__13220\ : ClkMux
    port map (
            O => \N__54335\,
            I => \N__53928\
        );

    \I__13219\ : ClkMux
    port map (
            O => \N__54334\,
            I => \N__53928\
        );

    \I__13218\ : ClkMux
    port map (
            O => \N__54333\,
            I => \N__53928\
        );

    \I__13217\ : ClkMux
    port map (
            O => \N__54332\,
            I => \N__53928\
        );

    \I__13216\ : ClkMux
    port map (
            O => \N__54331\,
            I => \N__53928\
        );

    \I__13215\ : ClkMux
    port map (
            O => \N__54330\,
            I => \N__53928\
        );

    \I__13214\ : ClkMux
    port map (
            O => \N__54329\,
            I => \N__53928\
        );

    \I__13213\ : ClkMux
    port map (
            O => \N__54328\,
            I => \N__53928\
        );

    \I__13212\ : ClkMux
    port map (
            O => \N__54327\,
            I => \N__53928\
        );

    \I__13211\ : ClkMux
    port map (
            O => \N__54326\,
            I => \N__53928\
        );

    \I__13210\ : ClkMux
    port map (
            O => \N__54325\,
            I => \N__53928\
        );

    \I__13209\ : ClkMux
    port map (
            O => \N__54324\,
            I => \N__53928\
        );

    \I__13208\ : ClkMux
    port map (
            O => \N__54323\,
            I => \N__53928\
        );

    \I__13207\ : ClkMux
    port map (
            O => \N__54322\,
            I => \N__53928\
        );

    \I__13206\ : ClkMux
    port map (
            O => \N__54321\,
            I => \N__53928\
        );

    \I__13205\ : ClkMux
    port map (
            O => \N__54320\,
            I => \N__53928\
        );

    \I__13204\ : ClkMux
    port map (
            O => \N__54319\,
            I => \N__53928\
        );

    \I__13203\ : ClkMux
    port map (
            O => \N__54318\,
            I => \N__53928\
        );

    \I__13202\ : ClkMux
    port map (
            O => \N__54317\,
            I => \N__53928\
        );

    \I__13201\ : ClkMux
    port map (
            O => \N__54316\,
            I => \N__53928\
        );

    \I__13200\ : ClkMux
    port map (
            O => \N__54315\,
            I => \N__53928\
        );

    \I__13199\ : ClkMux
    port map (
            O => \N__54314\,
            I => \N__53928\
        );

    \I__13198\ : ClkMux
    port map (
            O => \N__54313\,
            I => \N__53928\
        );

    \I__13197\ : ClkMux
    port map (
            O => \N__54312\,
            I => \N__53928\
        );

    \I__13196\ : ClkMux
    port map (
            O => \N__54311\,
            I => \N__53928\
        );

    \I__13195\ : ClkMux
    port map (
            O => \N__54310\,
            I => \N__53928\
        );

    \I__13194\ : ClkMux
    port map (
            O => \N__54309\,
            I => \N__53928\
        );

    \I__13193\ : ClkMux
    port map (
            O => \N__54308\,
            I => \N__53928\
        );

    \I__13192\ : ClkMux
    port map (
            O => \N__54307\,
            I => \N__53928\
        );

    \I__13191\ : ClkMux
    port map (
            O => \N__54306\,
            I => \N__53928\
        );

    \I__13190\ : ClkMux
    port map (
            O => \N__54305\,
            I => \N__53928\
        );

    \I__13189\ : ClkMux
    port map (
            O => \N__54304\,
            I => \N__53928\
        );

    \I__13188\ : ClkMux
    port map (
            O => \N__54303\,
            I => \N__53928\
        );

    \I__13187\ : ClkMux
    port map (
            O => \N__54302\,
            I => \N__53928\
        );

    \I__13186\ : ClkMux
    port map (
            O => \N__54301\,
            I => \N__53928\
        );

    \I__13185\ : ClkMux
    port map (
            O => \N__54300\,
            I => \N__53928\
        );

    \I__13184\ : ClkMux
    port map (
            O => \N__54299\,
            I => \N__53928\
        );

    \I__13183\ : ClkMux
    port map (
            O => \N__54298\,
            I => \N__53928\
        );

    \I__13182\ : ClkMux
    port map (
            O => \N__54297\,
            I => \N__53928\
        );

    \I__13181\ : ClkMux
    port map (
            O => \N__54296\,
            I => \N__53928\
        );

    \I__13180\ : ClkMux
    port map (
            O => \N__54295\,
            I => \N__53928\
        );

    \I__13179\ : ClkMux
    port map (
            O => \N__54294\,
            I => \N__53928\
        );

    \I__13178\ : ClkMux
    port map (
            O => \N__54293\,
            I => \N__53928\
        );

    \I__13177\ : ClkMux
    port map (
            O => \N__54292\,
            I => \N__53928\
        );

    \I__13176\ : ClkMux
    port map (
            O => \N__54291\,
            I => \N__53928\
        );

    \I__13175\ : ClkMux
    port map (
            O => \N__54290\,
            I => \N__53928\
        );

    \I__13174\ : ClkMux
    port map (
            O => \N__54289\,
            I => \N__53928\
        );

    \I__13173\ : ClkMux
    port map (
            O => \N__54288\,
            I => \N__53928\
        );

    \I__13172\ : ClkMux
    port map (
            O => \N__54287\,
            I => \N__53928\
        );

    \I__13171\ : ClkMux
    port map (
            O => \N__54286\,
            I => \N__53928\
        );

    \I__13170\ : ClkMux
    port map (
            O => \N__54285\,
            I => \N__53928\
        );

    \I__13169\ : ClkMux
    port map (
            O => \N__54284\,
            I => \N__53928\
        );

    \I__13168\ : ClkMux
    port map (
            O => \N__54283\,
            I => \N__53928\
        );

    \I__13167\ : ClkMux
    port map (
            O => \N__54282\,
            I => \N__53928\
        );

    \I__13166\ : ClkMux
    port map (
            O => \N__54281\,
            I => \N__53928\
        );

    \I__13165\ : ClkMux
    port map (
            O => \N__54280\,
            I => \N__53928\
        );

    \I__13164\ : ClkMux
    port map (
            O => \N__54279\,
            I => \N__53928\
        );

    \I__13163\ : ClkMux
    port map (
            O => \N__54278\,
            I => \N__53928\
        );

    \I__13162\ : ClkMux
    port map (
            O => \N__54277\,
            I => \N__53928\
        );

    \I__13161\ : ClkMux
    port map (
            O => \N__54276\,
            I => \N__53928\
        );

    \I__13160\ : ClkMux
    port map (
            O => \N__54275\,
            I => \N__53928\
        );

    \I__13159\ : ClkMux
    port map (
            O => \N__54274\,
            I => \N__53928\
        );

    \I__13158\ : ClkMux
    port map (
            O => \N__54273\,
            I => \N__53928\
        );

    \I__13157\ : ClkMux
    port map (
            O => \N__54272\,
            I => \N__53928\
        );

    \I__13156\ : ClkMux
    port map (
            O => \N__54271\,
            I => \N__53928\
        );

    \I__13155\ : ClkMux
    port map (
            O => \N__54270\,
            I => \N__53928\
        );

    \I__13154\ : ClkMux
    port map (
            O => \N__54269\,
            I => \N__53928\
        );

    \I__13153\ : GlobalMux
    port map (
            O => \N__53928\,
            I => \clk_32MHz\
        );

    \I__13152\ : CEMux
    port map (
            O => \N__53925\,
            I => \N__53921\
        );

    \I__13151\ : InMux
    port map (
            O => \N__53924\,
            I => \N__53918\
        );

    \I__13150\ : LocalMux
    port map (
            O => \N__53921\,
            I => \N__53914\
        );

    \I__13149\ : LocalMux
    port map (
            O => \N__53918\,
            I => \N__53911\
        );

    \I__13148\ : InMux
    port map (
            O => \N__53917\,
            I => \N__53908\
        );

    \I__13147\ : Odrv4
    port map (
            O => \N__53914\,
            I => n11860
        );

    \I__13146\ : Odrv4
    port map (
            O => \N__53911\,
            I => n11860
        );

    \I__13145\ : LocalMux
    port map (
            O => \N__53908\,
            I => n11860
        );

    \I__13144\ : SRMux
    port map (
            O => \N__53901\,
            I => \N__53898\
        );

    \I__13143\ : LocalMux
    port map (
            O => \N__53898\,
            I => n14655
        );

    \I__13142\ : CascadeMux
    port map (
            O => \N__53895\,
            I => \N__53892\
        );

    \I__13141\ : InMux
    port map (
            O => \N__53892\,
            I => \N__53889\
        );

    \I__13140\ : LocalMux
    port map (
            O => \N__53889\,
            I => \N__53886\
        );

    \I__13139\ : Odrv4
    port map (
            O => \N__53886\,
            I => buf_data_iac_12
        );

    \I__13138\ : InMux
    port map (
            O => \N__53883\,
            I => \N__53880\
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__53880\,
            I => \N__53877\
        );

    \I__13136\ : Odrv4
    port map (
            O => \N__53877\,
            I => n21451
        );

    \I__13135\ : InMux
    port map (
            O => \N__53874\,
            I => \N__53871\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__53871\,
            I => \N__53868\
        );

    \I__13133\ : Odrv4
    port map (
            O => \N__53868\,
            I => buf_data_iac_18
        );

    \I__13132\ : CascadeMux
    port map (
            O => \N__53865\,
            I => \N__53862\
        );

    \I__13131\ : InMux
    port map (
            O => \N__53862\,
            I => \N__53859\
        );

    \I__13130\ : LocalMux
    port map (
            O => \N__53859\,
            I => \N__53856\
        );

    \I__13129\ : Span4Mux_h
    port map (
            O => \N__53856\,
            I => \N__53853\
        );

    \I__13128\ : Odrv4
    port map (
            O => \N__53853\,
            I => n21151
        );

    \I__13127\ : InMux
    port map (
            O => \N__53850\,
            I => \N__53847\
        );

    \I__13126\ : LocalMux
    port map (
            O => \N__53847\,
            I => \N__53844\
        );

    \I__13125\ : Span12Mux_h
    port map (
            O => \N__53844\,
            I => \N__53841\
        );

    \I__13124\ : Odrv12
    port map (
            O => \N__53841\,
            I => n16_adj_1496
        );

    \I__13123\ : InMux
    port map (
            O => \N__53838\,
            I => \N__53835\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__53835\,
            I => n22399
        );

    \I__13121\ : InMux
    port map (
            O => \N__53832\,
            I => \N__53828\
        );

    \I__13120\ : CascadeMux
    port map (
            O => \N__53831\,
            I => \N__53825\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__53828\,
            I => \N__53822\
        );

    \I__13118\ : InMux
    port map (
            O => \N__53825\,
            I => \N__53819\
        );

    \I__13117\ : Span4Mux_h
    port map (
            O => \N__53822\,
            I => \N__53814\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__53819\,
            I => \N__53814\
        );

    \I__13115\ : Span4Mux_v
    port map (
            O => \N__53814\,
            I => \N__53810\
        );

    \I__13114\ : InMux
    port map (
            O => \N__53813\,
            I => \N__53807\
        );

    \I__13113\ : Span4Mux_h
    port map (
            O => \N__53810\,
            I => \N__53804\
        );

    \I__13112\ : LocalMux
    port map (
            O => \N__53807\,
            I => buf_adcdata_iac_13
        );

    \I__13111\ : Odrv4
    port map (
            O => \N__53804\,
            I => buf_adcdata_iac_13
        );

    \I__13110\ : InMux
    port map (
            O => \N__53799\,
            I => \N__53772\
        );

    \I__13109\ : InMux
    port map (
            O => \N__53798\,
            I => \N__53772\
        );

    \I__13108\ : InMux
    port map (
            O => \N__53797\,
            I => \N__53768\
        );

    \I__13107\ : CascadeMux
    port map (
            O => \N__53796\,
            I => \N__53758\
        );

    \I__13106\ : CascadeMux
    port map (
            O => \N__53795\,
            I => \N__53751\
        );

    \I__13105\ : InMux
    port map (
            O => \N__53794\,
            I => \N__53746\
        );

    \I__13104\ : InMux
    port map (
            O => \N__53793\,
            I => \N__53739\
        );

    \I__13103\ : InMux
    port map (
            O => \N__53792\,
            I => \N__53739\
        );

    \I__13102\ : InMux
    port map (
            O => \N__53791\,
            I => \N__53739\
        );

    \I__13101\ : InMux
    port map (
            O => \N__53790\,
            I => \N__53730\
        );

    \I__13100\ : InMux
    port map (
            O => \N__53789\,
            I => \N__53730\
        );

    \I__13099\ : InMux
    port map (
            O => \N__53788\,
            I => \N__53730\
        );

    \I__13098\ : InMux
    port map (
            O => \N__53787\,
            I => \N__53730\
        );

    \I__13097\ : InMux
    port map (
            O => \N__53786\,
            I => \N__53724\
        );

    \I__13096\ : InMux
    port map (
            O => \N__53785\,
            I => \N__53717\
        );

    \I__13095\ : InMux
    port map (
            O => \N__53784\,
            I => \N__53710\
        );

    \I__13094\ : InMux
    port map (
            O => \N__53783\,
            I => \N__53710\
        );

    \I__13093\ : InMux
    port map (
            O => \N__53782\,
            I => \N__53710\
        );

    \I__13092\ : InMux
    port map (
            O => \N__53781\,
            I => \N__53707\
        );

    \I__13091\ : InMux
    port map (
            O => \N__53780\,
            I => \N__53704\
        );

    \I__13090\ : InMux
    port map (
            O => \N__53779\,
            I => \N__53699\
        );

    \I__13089\ : InMux
    port map (
            O => \N__53778\,
            I => \N__53699\
        );

    \I__13088\ : InMux
    port map (
            O => \N__53777\,
            I => \N__53696\
        );

    \I__13087\ : LocalMux
    port map (
            O => \N__53772\,
            I => \N__53693\
        );

    \I__13086\ : InMux
    port map (
            O => \N__53771\,
            I => \N__53690\
        );

    \I__13085\ : LocalMux
    port map (
            O => \N__53768\,
            I => \N__53687\
        );

    \I__13084\ : InMux
    port map (
            O => \N__53767\,
            I => \N__53684\
        );

    \I__13083\ : InMux
    port map (
            O => \N__53766\,
            I => \N__53676\
        );

    \I__13082\ : InMux
    port map (
            O => \N__53765\,
            I => \N__53673\
        );

    \I__13081\ : InMux
    port map (
            O => \N__53764\,
            I => \N__53659\
        );

    \I__13080\ : InMux
    port map (
            O => \N__53763\,
            I => \N__53659\
        );

    \I__13079\ : InMux
    port map (
            O => \N__53762\,
            I => \N__53659\
        );

    \I__13078\ : InMux
    port map (
            O => \N__53761\,
            I => \N__53654\
        );

    \I__13077\ : InMux
    port map (
            O => \N__53758\,
            I => \N__53654\
        );

    \I__13076\ : InMux
    port map (
            O => \N__53757\,
            I => \N__53645\
        );

    \I__13075\ : InMux
    port map (
            O => \N__53756\,
            I => \N__53645\
        );

    \I__13074\ : InMux
    port map (
            O => \N__53755\,
            I => \N__53645\
        );

    \I__13073\ : InMux
    port map (
            O => \N__53754\,
            I => \N__53645\
        );

    \I__13072\ : InMux
    port map (
            O => \N__53751\,
            I => \N__53642\
        );

    \I__13071\ : InMux
    port map (
            O => \N__53750\,
            I => \N__53637\
        );

    \I__13070\ : InMux
    port map (
            O => \N__53749\,
            I => \N__53637\
        );

    \I__13069\ : LocalMux
    port map (
            O => \N__53746\,
            I => \N__53634\
        );

    \I__13068\ : LocalMux
    port map (
            O => \N__53739\,
            I => \N__53631\
        );

    \I__13067\ : LocalMux
    port map (
            O => \N__53730\,
            I => \N__53628\
        );

    \I__13066\ : InMux
    port map (
            O => \N__53729\,
            I => \N__53621\
        );

    \I__13065\ : InMux
    port map (
            O => \N__53728\,
            I => \N__53621\
        );

    \I__13064\ : InMux
    port map (
            O => \N__53727\,
            I => \N__53621\
        );

    \I__13063\ : LocalMux
    port map (
            O => \N__53724\,
            I => \N__53618\
        );

    \I__13062\ : InMux
    port map (
            O => \N__53723\,
            I => \N__53615\
        );

    \I__13061\ : InMux
    port map (
            O => \N__53722\,
            I => \N__53608\
        );

    \I__13060\ : InMux
    port map (
            O => \N__53721\,
            I => \N__53605\
        );

    \I__13059\ : InMux
    port map (
            O => \N__53720\,
            I => \N__53602\
        );

    \I__13058\ : LocalMux
    port map (
            O => \N__53717\,
            I => \N__53597\
        );

    \I__13057\ : LocalMux
    port map (
            O => \N__53710\,
            I => \N__53597\
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__53707\,
            I => \N__53590\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__53704\,
            I => \N__53590\
        );

    \I__13054\ : LocalMux
    port map (
            O => \N__53699\,
            I => \N__53590\
        );

    \I__13053\ : LocalMux
    port map (
            O => \N__53696\,
            I => \N__53585\
        );

    \I__13052\ : Span4Mux_v
    port map (
            O => \N__53693\,
            I => \N__53585\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__53690\,
            I => \N__53580\
        );

    \I__13050\ : Span4Mux_h
    port map (
            O => \N__53687\,
            I => \N__53580\
        );

    \I__13049\ : LocalMux
    port map (
            O => \N__53684\,
            I => \N__53577\
        );

    \I__13048\ : InMux
    port map (
            O => \N__53683\,
            I => \N__53568\
        );

    \I__13047\ : InMux
    port map (
            O => \N__53682\,
            I => \N__53568\
        );

    \I__13046\ : InMux
    port map (
            O => \N__53681\,
            I => \N__53568\
        );

    \I__13045\ : InMux
    port map (
            O => \N__53680\,
            I => \N__53568\
        );

    \I__13044\ : InMux
    port map (
            O => \N__53679\,
            I => \N__53565\
        );

    \I__13043\ : LocalMux
    port map (
            O => \N__53676\,
            I => \N__53562\
        );

    \I__13042\ : LocalMux
    port map (
            O => \N__53673\,
            I => \N__53559\
        );

    \I__13041\ : InMux
    port map (
            O => \N__53672\,
            I => \N__53556\
        );

    \I__13040\ : InMux
    port map (
            O => \N__53671\,
            I => \N__53549\
        );

    \I__13039\ : InMux
    port map (
            O => \N__53670\,
            I => \N__53545\
        );

    \I__13038\ : InMux
    port map (
            O => \N__53669\,
            I => \N__53536\
        );

    \I__13037\ : InMux
    port map (
            O => \N__53668\,
            I => \N__53536\
        );

    \I__13036\ : InMux
    port map (
            O => \N__53667\,
            I => \N__53536\
        );

    \I__13035\ : InMux
    port map (
            O => \N__53666\,
            I => \N__53536\
        );

    \I__13034\ : LocalMux
    port map (
            O => \N__53659\,
            I => \N__53529\
        );

    \I__13033\ : LocalMux
    port map (
            O => \N__53654\,
            I => \N__53529\
        );

    \I__13032\ : LocalMux
    port map (
            O => \N__53645\,
            I => \N__53529\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__53642\,
            I => \N__53526\
        );

    \I__13030\ : LocalMux
    port map (
            O => \N__53637\,
            I => \N__53523\
        );

    \I__13029\ : Span4Mux_h
    port map (
            O => \N__53634\,
            I => \N__53520\
        );

    \I__13028\ : Span4Mux_h
    port map (
            O => \N__53631\,
            I => \N__53513\
        );

    \I__13027\ : Span4Mux_v
    port map (
            O => \N__53628\,
            I => \N__53513\
        );

    \I__13026\ : LocalMux
    port map (
            O => \N__53621\,
            I => \N__53513\
        );

    \I__13025\ : Span4Mux_h
    port map (
            O => \N__53618\,
            I => \N__53510\
        );

    \I__13024\ : LocalMux
    port map (
            O => \N__53615\,
            I => \N__53507\
        );

    \I__13023\ : InMux
    port map (
            O => \N__53614\,
            I => \N__53502\
        );

    \I__13022\ : InMux
    port map (
            O => \N__53613\,
            I => \N__53502\
        );

    \I__13021\ : InMux
    port map (
            O => \N__53612\,
            I => \N__53499\
        );

    \I__13020\ : InMux
    port map (
            O => \N__53611\,
            I => \N__53496\
        );

    \I__13019\ : LocalMux
    port map (
            O => \N__53608\,
            I => \N__53493\
        );

    \I__13018\ : LocalMux
    port map (
            O => \N__53605\,
            I => \N__53490\
        );

    \I__13017\ : LocalMux
    port map (
            O => \N__53602\,
            I => \N__53486\
        );

    \I__13016\ : Span4Mux_h
    port map (
            O => \N__53597\,
            I => \N__53483\
        );

    \I__13015\ : Span4Mux_h
    port map (
            O => \N__53590\,
            I => \N__53480\
        );

    \I__13014\ : Span4Mux_h
    port map (
            O => \N__53585\,
            I => \N__53475\
        );

    \I__13013\ : Span4Mux_v
    port map (
            O => \N__53580\,
            I => \N__53475\
        );

    \I__13012\ : Span4Mux_h
    port map (
            O => \N__53577\,
            I => \N__53472\
        );

    \I__13011\ : LocalMux
    port map (
            O => \N__53568\,
            I => \N__53469\
        );

    \I__13010\ : LocalMux
    port map (
            O => \N__53565\,
            I => \N__53466\
        );

    \I__13009\ : Span4Mux_h
    port map (
            O => \N__53562\,
            I => \N__53459\
        );

    \I__13008\ : Span4Mux_v
    port map (
            O => \N__53559\,
            I => \N__53459\
        );

    \I__13007\ : LocalMux
    port map (
            O => \N__53556\,
            I => \N__53459\
        );

    \I__13006\ : InMux
    port map (
            O => \N__53555\,
            I => \N__53454\
        );

    \I__13005\ : InMux
    port map (
            O => \N__53554\,
            I => \N__53447\
        );

    \I__13004\ : InMux
    port map (
            O => \N__53553\,
            I => \N__53447\
        );

    \I__13003\ : InMux
    port map (
            O => \N__53552\,
            I => \N__53447\
        );

    \I__13002\ : LocalMux
    port map (
            O => \N__53549\,
            I => \N__53444\
        );

    \I__13001\ : InMux
    port map (
            O => \N__53548\,
            I => \N__53441\
        );

    \I__13000\ : LocalMux
    port map (
            O => \N__53545\,
            I => \N__53430\
        );

    \I__12999\ : LocalMux
    port map (
            O => \N__53536\,
            I => \N__53430\
        );

    \I__12998\ : Span4Mux_v
    port map (
            O => \N__53529\,
            I => \N__53430\
        );

    \I__12997\ : Span4Mux_v
    port map (
            O => \N__53526\,
            I => \N__53430\
        );

    \I__12996\ : Span4Mux_v
    port map (
            O => \N__53523\,
            I => \N__53430\
        );

    \I__12995\ : Span4Mux_h
    port map (
            O => \N__53520\,
            I => \N__53423\
        );

    \I__12994\ : Span4Mux_h
    port map (
            O => \N__53513\,
            I => \N__53423\
        );

    \I__12993\ : Span4Mux_h
    port map (
            O => \N__53510\,
            I => \N__53423\
        );

    \I__12992\ : Span4Mux_v
    port map (
            O => \N__53507\,
            I => \N__53420\
        );

    \I__12991\ : LocalMux
    port map (
            O => \N__53502\,
            I => \N__53409\
        );

    \I__12990\ : LocalMux
    port map (
            O => \N__53499\,
            I => \N__53409\
        );

    \I__12989\ : LocalMux
    port map (
            O => \N__53496\,
            I => \N__53409\
        );

    \I__12988\ : Span12Mux_v
    port map (
            O => \N__53493\,
            I => \N__53409\
        );

    \I__12987\ : Span12Mux_v
    port map (
            O => \N__53490\,
            I => \N__53409\
        );

    \I__12986\ : InMux
    port map (
            O => \N__53489\,
            I => \N__53406\
        );

    \I__12985\ : Span4Mux_v
    port map (
            O => \N__53486\,
            I => \N__53397\
        );

    \I__12984\ : Span4Mux_h
    port map (
            O => \N__53483\,
            I => \N__53397\
        );

    \I__12983\ : Span4Mux_h
    port map (
            O => \N__53480\,
            I => \N__53397\
        );

    \I__12982\ : Span4Mux_h
    port map (
            O => \N__53475\,
            I => \N__53397\
        );

    \I__12981\ : Span4Mux_h
    port map (
            O => \N__53472\,
            I => \N__53388\
        );

    \I__12980\ : Span4Mux_h
    port map (
            O => \N__53469\,
            I => \N__53388\
        );

    \I__12979\ : Span4Mux_v
    port map (
            O => \N__53466\,
            I => \N__53388\
        );

    \I__12978\ : Span4Mux_h
    port map (
            O => \N__53459\,
            I => \N__53388\
        );

    \I__12977\ : InMux
    port map (
            O => \N__53458\,
            I => \N__53383\
        );

    \I__12976\ : InMux
    port map (
            O => \N__53457\,
            I => \N__53383\
        );

    \I__12975\ : LocalMux
    port map (
            O => \N__53454\,
            I => comm_cmd_2
        );

    \I__12974\ : LocalMux
    port map (
            O => \N__53447\,
            I => comm_cmd_2
        );

    \I__12973\ : Odrv4
    port map (
            O => \N__53444\,
            I => comm_cmd_2
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__53441\,
            I => comm_cmd_2
        );

    \I__12971\ : Odrv4
    port map (
            O => \N__53430\,
            I => comm_cmd_2
        );

    \I__12970\ : Odrv4
    port map (
            O => \N__53423\,
            I => comm_cmd_2
        );

    \I__12969\ : Odrv4
    port map (
            O => \N__53420\,
            I => comm_cmd_2
        );

    \I__12968\ : Odrv12
    port map (
            O => \N__53409\,
            I => comm_cmd_2
        );

    \I__12967\ : LocalMux
    port map (
            O => \N__53406\,
            I => comm_cmd_2
        );

    \I__12966\ : Odrv4
    port map (
            O => \N__53397\,
            I => comm_cmd_2
        );

    \I__12965\ : Odrv4
    port map (
            O => \N__53388\,
            I => comm_cmd_2
        );

    \I__12964\ : LocalMux
    port map (
            O => \N__53383\,
            I => comm_cmd_2
        );

    \I__12963\ : InMux
    port map (
            O => \N__53358\,
            I => \N__53355\
        );

    \I__12962\ : LocalMux
    port map (
            O => \N__53355\,
            I => n22402
        );

    \I__12961\ : InMux
    port map (
            O => \N__53352\,
            I => \N__53348\
        );

    \I__12960\ : InMux
    port map (
            O => \N__53351\,
            I => \N__53345\
        );

    \I__12959\ : LocalMux
    port map (
            O => \N__53348\,
            I => \N__53342\
        );

    \I__12958\ : LocalMux
    port map (
            O => \N__53345\,
            I => \N__53339\
        );

    \I__12957\ : Odrv4
    port map (
            O => \N__53342\,
            I => \ADC_VDC.genclk.n21444\
        );

    \I__12956\ : Odrv4
    port map (
            O => \N__53339\,
            I => \ADC_VDC.genclk.n21444\
        );

    \I__12955\ : SRMux
    port map (
            O => \N__53334\,
            I => \N__53331\
        );

    \I__12954\ : LocalMux
    port map (
            O => \N__53331\,
            I => \N__53328\
        );

    \I__12953\ : Odrv12
    port map (
            O => \N__53328\,
            I => \comm_spi.DOUT_7__N_747\
        );

    \I__12952\ : ClkMux
    port map (
            O => \N__53325\,
            I => \N__53321\
        );

    \I__12951\ : IoInMux
    port map (
            O => \N__53324\,
            I => \N__53315\
        );

    \I__12950\ : LocalMux
    port map (
            O => \N__53321\,
            I => \N__53312\
        );

    \I__12949\ : ClkMux
    port map (
            O => \N__53320\,
            I => \N__53309\
        );

    \I__12948\ : ClkMux
    port map (
            O => \N__53319\,
            I => \N__53306\
        );

    \I__12947\ : ClkMux
    port map (
            O => \N__53318\,
            I => \N__53303\
        );

    \I__12946\ : LocalMux
    port map (
            O => \N__53315\,
            I => \N__53295\
        );

    \I__12945\ : Span4Mux_v
    port map (
            O => \N__53312\,
            I => \N__53288\
        );

    \I__12944\ : LocalMux
    port map (
            O => \N__53309\,
            I => \N__53288\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__53306\,
            I => \N__53285\
        );

    \I__12942\ : LocalMux
    port map (
            O => \N__53303\,
            I => \N__53282\
        );

    \I__12941\ : ClkMux
    port map (
            O => \N__53302\,
            I => \N__53279\
        );

    \I__12940\ : ClkMux
    port map (
            O => \N__53301\,
            I => \N__53272\
        );

    \I__12939\ : ClkMux
    port map (
            O => \N__53300\,
            I => \N__53269\
        );

    \I__12938\ : ClkMux
    port map (
            O => \N__53299\,
            I => \N__53266\
        );

    \I__12937\ : ClkMux
    port map (
            O => \N__53298\,
            I => \N__53262\
        );

    \I__12936\ : Span4Mux_s3_h
    port map (
            O => \N__53295\,
            I => \N__53257\
        );

    \I__12935\ : ClkMux
    port map (
            O => \N__53294\,
            I => \N__53250\
        );

    \I__12934\ : ClkMux
    port map (
            O => \N__53293\,
            I => \N__53247\
        );

    \I__12933\ : Span4Mux_v
    port map (
            O => \N__53288\,
            I => \N__53244\
        );

    \I__12932\ : Span4Mux_h
    port map (
            O => \N__53285\,
            I => \N__53237\
        );

    \I__12931\ : Span4Mux_v
    port map (
            O => \N__53282\,
            I => \N__53237\
        );

    \I__12930\ : LocalMux
    port map (
            O => \N__53279\,
            I => \N__53237\
        );

    \I__12929\ : ClkMux
    port map (
            O => \N__53278\,
            I => \N__53234\
        );

    \I__12928\ : ClkMux
    port map (
            O => \N__53277\,
            I => \N__53231\
        );

    \I__12927\ : ClkMux
    port map (
            O => \N__53276\,
            I => \N__53228\
        );

    \I__12926\ : ClkMux
    port map (
            O => \N__53275\,
            I => \N__53225\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__53272\,
            I => \N__53220\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__53269\,
            I => \N__53220\
        );

    \I__12923\ : LocalMux
    port map (
            O => \N__53266\,
            I => \N__53217\
        );

    \I__12922\ : ClkMux
    port map (
            O => \N__53265\,
            I => \N__53214\
        );

    \I__12921\ : LocalMux
    port map (
            O => \N__53262\,
            I => \N__53211\
        );

    \I__12920\ : ClkMux
    port map (
            O => \N__53261\,
            I => \N__53208\
        );

    \I__12919\ : ClkMux
    port map (
            O => \N__53260\,
            I => \N__53204\
        );

    \I__12918\ : Span4Mux_h
    port map (
            O => \N__53257\,
            I => \N__53201\
        );

    \I__12917\ : ClkMux
    port map (
            O => \N__53256\,
            I => \N__53198\
        );

    \I__12916\ : ClkMux
    port map (
            O => \N__53255\,
            I => \N__53195\
        );

    \I__12915\ : ClkMux
    port map (
            O => \N__53254\,
            I => \N__53191\
        );

    \I__12914\ : ClkMux
    port map (
            O => \N__53253\,
            I => \N__53188\
        );

    \I__12913\ : LocalMux
    port map (
            O => \N__53250\,
            I => \N__53183\
        );

    \I__12912\ : LocalMux
    port map (
            O => \N__53247\,
            I => \N__53183\
        );

    \I__12911\ : Span4Mux_v
    port map (
            O => \N__53244\,
            I => \N__53176\
        );

    \I__12910\ : Span4Mux_v
    port map (
            O => \N__53237\,
            I => \N__53176\
        );

    \I__12909\ : LocalMux
    port map (
            O => \N__53234\,
            I => \N__53176\
        );

    \I__12908\ : LocalMux
    port map (
            O => \N__53231\,
            I => \N__53173\
        );

    \I__12907\ : LocalMux
    port map (
            O => \N__53228\,
            I => \N__53168\
        );

    \I__12906\ : LocalMux
    port map (
            O => \N__53225\,
            I => \N__53168\
        );

    \I__12905\ : Span4Mux_v
    port map (
            O => \N__53220\,
            I => \N__53163\
        );

    \I__12904\ : Span4Mux_v
    port map (
            O => \N__53217\,
            I => \N__53163\
        );

    \I__12903\ : LocalMux
    port map (
            O => \N__53214\,
            I => \N__53160\
        );

    \I__12902\ : Span4Mux_v
    port map (
            O => \N__53211\,
            I => \N__53155\
        );

    \I__12901\ : LocalMux
    port map (
            O => \N__53208\,
            I => \N__53155\
        );

    \I__12900\ : ClkMux
    port map (
            O => \N__53207\,
            I => \N__53152\
        );

    \I__12899\ : LocalMux
    port map (
            O => \N__53204\,
            I => \N__53149\
        );

    \I__12898\ : Span4Mux_h
    port map (
            O => \N__53201\,
            I => \N__53142\
        );

    \I__12897\ : LocalMux
    port map (
            O => \N__53198\,
            I => \N__53142\
        );

    \I__12896\ : LocalMux
    port map (
            O => \N__53195\,
            I => \N__53142\
        );

    \I__12895\ : ClkMux
    port map (
            O => \N__53194\,
            I => \N__53139\
        );

    \I__12894\ : LocalMux
    port map (
            O => \N__53191\,
            I => \N__53132\
        );

    \I__12893\ : LocalMux
    port map (
            O => \N__53188\,
            I => \N__53132\
        );

    \I__12892\ : Span4Mux_v
    port map (
            O => \N__53183\,
            I => \N__53132\
        );

    \I__12891\ : Span4Mux_h
    port map (
            O => \N__53176\,
            I => \N__53129\
        );

    \I__12890\ : Span4Mux_h
    port map (
            O => \N__53173\,
            I => \N__53124\
        );

    \I__12889\ : Span4Mux_v
    port map (
            O => \N__53168\,
            I => \N__53124\
        );

    \I__12888\ : Span4Mux_h
    port map (
            O => \N__53163\,
            I => \N__53119\
        );

    \I__12887\ : Span4Mux_v
    port map (
            O => \N__53160\,
            I => \N__53119\
        );

    \I__12886\ : Span4Mux_h
    port map (
            O => \N__53155\,
            I => \N__53114\
        );

    \I__12885\ : LocalMux
    port map (
            O => \N__53152\,
            I => \N__53114\
        );

    \I__12884\ : Span4Mux_h
    port map (
            O => \N__53149\,
            I => \N__53109\
        );

    \I__12883\ : Span4Mux_h
    port map (
            O => \N__53142\,
            I => \N__53109\
        );

    \I__12882\ : LocalMux
    port map (
            O => \N__53139\,
            I => \N__53106\
        );

    \I__12881\ : Sp12to4
    port map (
            O => \N__53132\,
            I => \N__53103\
        );

    \I__12880\ : Span4Mux_h
    port map (
            O => \N__53129\,
            I => \N__53100\
        );

    \I__12879\ : Span4Mux_h
    port map (
            O => \N__53124\,
            I => \N__53093\
        );

    \I__12878\ : Span4Mux_v
    port map (
            O => \N__53119\,
            I => \N__53093\
        );

    \I__12877\ : Span4Mux_v
    port map (
            O => \N__53114\,
            I => \N__53093\
        );

    \I__12876\ : Span4Mux_h
    port map (
            O => \N__53109\,
            I => \N__53088\
        );

    \I__12875\ : Span4Mux_v
    port map (
            O => \N__53106\,
            I => \N__53088\
        );

    \I__12874\ : Span12Mux_h
    port map (
            O => \N__53103\,
            I => \N__53085\
        );

    \I__12873\ : Span4Mux_h
    port map (
            O => \N__53100\,
            I => \N__53082\
        );

    \I__12872\ : Sp12to4
    port map (
            O => \N__53093\,
            I => \N__53079\
        );

    \I__12871\ : Span4Mux_h
    port map (
            O => \N__53088\,
            I => \N__53076\
        );

    \I__12870\ : Odrv12
    port map (
            O => \N__53085\,
            I => \VDC_CLK\
        );

    \I__12869\ : Odrv4
    port map (
            O => \N__53082\,
            I => \VDC_CLK\
        );

    \I__12868\ : Odrv12
    port map (
            O => \N__53079\,
            I => \VDC_CLK\
        );

    \I__12867\ : Odrv4
    port map (
            O => \N__53076\,
            I => \VDC_CLK\
        );

    \I__12866\ : InMux
    port map (
            O => \N__53067\,
            I => \N__53064\
        );

    \I__12865\ : LocalMux
    port map (
            O => \N__53064\,
            I => \comm_spi.n14614\
        );

    \I__12864\ : InMux
    port map (
            O => \N__53061\,
            I => \N__53058\
        );

    \I__12863\ : LocalMux
    port map (
            O => \N__53058\,
            I => \comm_spi.n14615\
        );

    \I__12862\ : InMux
    port map (
            O => \N__53055\,
            I => \N__53052\
        );

    \I__12861\ : LocalMux
    port map (
            O => \N__53052\,
            I => \N__53047\
        );

    \I__12860\ : InMux
    port map (
            O => \N__53051\,
            I => \N__53044\
        );

    \I__12859\ : InMux
    port map (
            O => \N__53050\,
            I => \N__53041\
        );

    \I__12858\ : Span4Mux_v
    port map (
            O => \N__53047\,
            I => \N__53030\
        );

    \I__12857\ : LocalMux
    port map (
            O => \N__53044\,
            I => \N__53030\
        );

    \I__12856\ : LocalMux
    port map (
            O => \N__53041\,
            I => \N__53027\
        );

    \I__12855\ : InMux
    port map (
            O => \N__53040\,
            I => \N__53022\
        );

    \I__12854\ : InMux
    port map (
            O => \N__53039\,
            I => \N__53022\
        );

    \I__12853\ : InMux
    port map (
            O => \N__53038\,
            I => \N__53019\
        );

    \I__12852\ : InMux
    port map (
            O => \N__53037\,
            I => \N__53016\
        );

    \I__12851\ : InMux
    port map (
            O => \N__53036\,
            I => \N__53013\
        );

    \I__12850\ : InMux
    port map (
            O => \N__53035\,
            I => \N__53010\
        );

    \I__12849\ : Span4Mux_v
    port map (
            O => \N__53030\,
            I => \N__53007\
        );

    \I__12848\ : Sp12to4
    port map (
            O => \N__53027\,
            I => \N__53000\
        );

    \I__12847\ : LocalMux
    port map (
            O => \N__53022\,
            I => \N__53000\
        );

    \I__12846\ : LocalMux
    port map (
            O => \N__53019\,
            I => \N__53000\
        );

    \I__12845\ : LocalMux
    port map (
            O => \N__53016\,
            I => \N__52995\
        );

    \I__12844\ : LocalMux
    port map (
            O => \N__53013\,
            I => \N__52995\
        );

    \I__12843\ : LocalMux
    port map (
            O => \N__53010\,
            I => \N__52992\
        );

    \I__12842\ : Span4Mux_h
    port map (
            O => \N__53007\,
            I => \N__52989\
        );

    \I__12841\ : Span12Mux_v
    port map (
            O => \N__53000\,
            I => \N__52986\
        );

    \I__12840\ : Span4Mux_h
    port map (
            O => \N__52995\,
            I => \N__52983\
        );

    \I__12839\ : Span4Mux_v
    port map (
            O => \N__52992\,
            I => \N__52980\
        );

    \I__12838\ : Odrv4
    port map (
            O => \N__52989\,
            I => comm_rx_buf_0
        );

    \I__12837\ : Odrv12
    port map (
            O => \N__52986\,
            I => comm_rx_buf_0
        );

    \I__12836\ : Odrv4
    port map (
            O => \N__52983\,
            I => comm_rx_buf_0
        );

    \I__12835\ : Odrv4
    port map (
            O => \N__52980\,
            I => comm_rx_buf_0
        );

    \I__12834\ : InMux
    port map (
            O => \N__52971\,
            I => \N__52966\
        );

    \I__12833\ : InMux
    port map (
            O => \N__52970\,
            I => \N__52963\
        );

    \I__12832\ : InMux
    port map (
            O => \N__52969\,
            I => \N__52960\
        );

    \I__12831\ : LocalMux
    port map (
            O => \N__52966\,
            I => \comm_spi.n22866\
        );

    \I__12830\ : LocalMux
    port map (
            O => \N__52963\,
            I => \comm_spi.n22866\
        );

    \I__12829\ : LocalMux
    port map (
            O => \N__52960\,
            I => \comm_spi.n22866\
        );

    \I__12828\ : CascadeMux
    port map (
            O => \N__52953\,
            I => \comm_spi.n22866_cascade_\
        );

    \I__12827\ : InMux
    port map (
            O => \N__52950\,
            I => \N__52945\
        );

    \I__12826\ : InMux
    port map (
            O => \N__52949\,
            I => \N__52942\
        );

    \I__12825\ : InMux
    port map (
            O => \N__52948\,
            I => \N__52939\
        );

    \I__12824\ : LocalMux
    port map (
            O => \N__52945\,
            I => \N__52934\
        );

    \I__12823\ : LocalMux
    port map (
            O => \N__52942\,
            I => \N__52934\
        );

    \I__12822\ : LocalMux
    port map (
            O => \N__52939\,
            I => \N__52931\
        );

    \I__12821\ : Span4Mux_v
    port map (
            O => \N__52934\,
            I => \N__52928\
        );

    \I__12820\ : Odrv4
    port map (
            O => \N__52931\,
            I => \comm_spi.n14601\
        );

    \I__12819\ : Odrv4
    port map (
            O => \N__52928\,
            I => \comm_spi.n14601\
        );

    \I__12818\ : CascadeMux
    port map (
            O => \N__52923\,
            I => \comm_spi.imosi_cascade_\
        );

    \I__12817\ : SRMux
    port map (
            O => \N__52920\,
            I => \N__52917\
        );

    \I__12816\ : LocalMux
    port map (
            O => \N__52917\,
            I => \N__52914\
        );

    \I__12815\ : Span4Mux_v
    port map (
            O => \N__52914\,
            I => \N__52911\
        );

    \I__12814\ : Odrv4
    port map (
            O => \N__52911\,
            I => \comm_spi.DOUT_7__N_746\
        );

    \I__12813\ : InMux
    port map (
            O => \N__52908\,
            I => \N__52901\
        );

    \I__12812\ : InMux
    port map (
            O => \N__52907\,
            I => \N__52901\
        );

    \I__12811\ : InMux
    port map (
            O => \N__52906\,
            I => \N__52898\
        );

    \I__12810\ : LocalMux
    port map (
            O => \N__52901\,
            I => \N__52895\
        );

    \I__12809\ : LocalMux
    port map (
            O => \N__52898\,
            I => \N__52890\
        );

    \I__12808\ : Span4Mux_h
    port map (
            O => \N__52895\,
            I => \N__52887\
        );

    \I__12807\ : InMux
    port map (
            O => \N__52894\,
            I => \N__52882\
        );

    \I__12806\ : InMux
    port map (
            O => \N__52893\,
            I => \N__52882\
        );

    \I__12805\ : Odrv12
    port map (
            O => \N__52890\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__12804\ : Odrv4
    port map (
            O => \N__52887\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__12803\ : LocalMux
    port map (
            O => \N__52882\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__12802\ : InMux
    port map (
            O => \N__52875\,
            I => \N__52871\
        );

    \I__12801\ : InMux
    port map (
            O => \N__52874\,
            I => \N__52868\
        );

    \I__12800\ : LocalMux
    port map (
            O => \N__52871\,
            I => \comm_spi.imosi\
        );

    \I__12799\ : LocalMux
    port map (
            O => \N__52868\,
            I => \comm_spi.imosi\
        );

    \I__12798\ : InMux
    port map (
            O => \N__52863\,
            I => \N__52859\
        );

    \I__12797\ : InMux
    port map (
            O => \N__52862\,
            I => \N__52856\
        );

    \I__12796\ : LocalMux
    port map (
            O => \N__52859\,
            I => \comm_spi.n22863\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__52856\,
            I => \comm_spi.n22863\
        );

    \I__12794\ : InMux
    port map (
            O => \N__52851\,
            I => \N__52848\
        );

    \I__12793\ : LocalMux
    port map (
            O => \N__52848\,
            I => \N__52845\
        );

    \I__12792\ : Span4Mux_h
    port map (
            O => \N__52845\,
            I => \N__52841\
        );

    \I__12791\ : InMux
    port map (
            O => \N__52844\,
            I => \N__52837\
        );

    \I__12790\ : Span4Mux_h
    port map (
            O => \N__52841\,
            I => \N__52834\
        );

    \I__12789\ : InMux
    port map (
            O => \N__52840\,
            I => \N__52831\
        );

    \I__12788\ : LocalMux
    port map (
            O => \N__52837\,
            I => req_data_cnt_5
        );

    \I__12787\ : Odrv4
    port map (
            O => \N__52834\,
            I => req_data_cnt_5
        );

    \I__12786\ : LocalMux
    port map (
            O => \N__52831\,
            I => req_data_cnt_5
        );

    \I__12785\ : CascadeMux
    port map (
            O => \N__52824\,
            I => \n22345_cascade_\
        );

    \I__12784\ : InMux
    port map (
            O => \N__52821\,
            I => \N__52818\
        );

    \I__12783\ : LocalMux
    port map (
            O => \N__52818\,
            I => \N__52815\
        );

    \I__12782\ : Span4Mux_h
    port map (
            O => \N__52815\,
            I => \N__52812\
        );

    \I__12781\ : Span4Mux_h
    port map (
            O => \N__52812\,
            I => \N__52807\
        );

    \I__12780\ : InMux
    port map (
            O => \N__52811\,
            I => \N__52802\
        );

    \I__12779\ : InMux
    port map (
            O => \N__52810\,
            I => \N__52802\
        );

    \I__12778\ : Odrv4
    port map (
            O => \N__52807\,
            I => \acadc_skipCount_5\
        );

    \I__12777\ : LocalMux
    port map (
            O => \N__52802\,
            I => \acadc_skipCount_5\
        );

    \I__12776\ : CascadeMux
    port map (
            O => \N__52797\,
            I => \n22348_cascade_\
        );

    \I__12775\ : InMux
    port map (
            O => \N__52794\,
            I => \N__52791\
        );

    \I__12774\ : LocalMux
    port map (
            O => \N__52791\,
            I => n30_adj_1500
        );

    \I__12773\ : InMux
    port map (
            O => \N__52788\,
            I => \N__52784\
        );

    \I__12772\ : InMux
    port map (
            O => \N__52787\,
            I => \N__52781\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__52784\,
            I => \N__52778\
        );

    \I__12770\ : LocalMux
    port map (
            O => \N__52781\,
            I => \N__52775\
        );

    \I__12769\ : Span4Mux_v
    port map (
            O => \N__52778\,
            I => \N__52771\
        );

    \I__12768\ : Span4Mux_h
    port map (
            O => \N__52775\,
            I => \N__52768\
        );

    \I__12767\ : InMux
    port map (
            O => \N__52774\,
            I => \N__52765\
        );

    \I__12766\ : Sp12to4
    port map (
            O => \N__52771\,
            I => \N__52762\
        );

    \I__12765\ : Span4Mux_h
    port map (
            O => \N__52768\,
            I => \N__52759\
        );

    \I__12764\ : LocalMux
    port map (
            O => \N__52765\,
            I => buf_adcdata_iac_11
        );

    \I__12763\ : Odrv12
    port map (
            O => \N__52762\,
            I => buf_adcdata_iac_11
        );

    \I__12762\ : Odrv4
    port map (
            O => \N__52759\,
            I => buf_adcdata_iac_11
        );

    \I__12761\ : InMux
    port map (
            O => \N__52752\,
            I => \N__52749\
        );

    \I__12760\ : LocalMux
    port map (
            O => \N__52749\,
            I => n16_adj_1514
        );

    \I__12759\ : InMux
    port map (
            O => \N__52746\,
            I => \N__52743\
        );

    \I__12758\ : LocalMux
    port map (
            O => \N__52743\,
            I => \N__52740\
        );

    \I__12757\ : Span4Mux_h
    port map (
            O => \N__52740\,
            I => \N__52737\
        );

    \I__12756\ : Odrv4
    port map (
            O => \N__52737\,
            I => n21126
        );

    \I__12755\ : InMux
    port map (
            O => \N__52734\,
            I => \N__52731\
        );

    \I__12754\ : LocalMux
    port map (
            O => \N__52731\,
            I => \N__52728\
        );

    \I__12753\ : Span4Mux_h
    port map (
            O => \N__52728\,
            I => \N__52725\
        );

    \I__12752\ : Odrv4
    port map (
            O => \N__52725\,
            I => buf_data_iac_10
        );

    \I__12751\ : CascadeMux
    port map (
            O => \N__52722\,
            I => \N__52719\
        );

    \I__12750\ : InMux
    port map (
            O => \N__52719\,
            I => \N__52716\
        );

    \I__12749\ : LocalMux
    port map (
            O => \N__52716\,
            I => \N__52713\
        );

    \I__12748\ : Span4Mux_v
    port map (
            O => \N__52713\,
            I => \N__52710\
        );

    \I__12747\ : Odrv4
    port map (
            O => \N__52710\,
            I => n21564
        );

    \I__12746\ : InMux
    port map (
            O => \N__52707\,
            I => \N__52704\
        );

    \I__12745\ : LocalMux
    port map (
            O => \N__52704\,
            I => \N__52701\
        );

    \I__12744\ : Span4Mux_v
    port map (
            O => \N__52701\,
            I => \N__52698\
        );

    \I__12743\ : Odrv4
    port map (
            O => \N__52698\,
            I => buf_data_iac_8
        );

    \I__12742\ : InMux
    port map (
            O => \N__52695\,
            I => \N__52692\
        );

    \I__12741\ : LocalMux
    port map (
            O => \N__52692\,
            I => \N__52689\
        );

    \I__12740\ : Span4Mux_h
    port map (
            O => \N__52689\,
            I => \N__52686\
        );

    \I__12739\ : Span4Mux_v
    port map (
            O => \N__52686\,
            I => \N__52683\
        );

    \I__12738\ : Odrv4
    port map (
            O => \N__52683\,
            I => n21218
        );

    \I__12737\ : InMux
    port map (
            O => \N__52680\,
            I => \N__52677\
        );

    \I__12736\ : LocalMux
    port map (
            O => \N__52677\,
            I => \N__52674\
        );

    \I__12735\ : Odrv4
    port map (
            O => \N__52674\,
            I => buf_data_iac_23
        );

    \I__12734\ : CascadeMux
    port map (
            O => \N__52671\,
            I => \N__52668\
        );

    \I__12733\ : InMux
    port map (
            O => \N__52668\,
            I => \N__52665\
        );

    \I__12732\ : LocalMux
    port map (
            O => \N__52665\,
            I => \N__52662\
        );

    \I__12731\ : Span12Mux_h
    port map (
            O => \N__52662\,
            I => \N__52659\
        );

    \I__12730\ : Span12Mux_h
    port map (
            O => \N__52659\,
            I => \N__52656\
        );

    \I__12729\ : Span12Mux_v
    port map (
            O => \N__52656\,
            I => \N__52653\
        );

    \I__12728\ : Odrv12
    port map (
            O => \N__52653\,
            I => n21364
        );

    \I__12727\ : CEMux
    port map (
            O => \N__52650\,
            I => \N__52647\
        );

    \I__12726\ : LocalMux
    port map (
            O => \N__52647\,
            I => \N__52644\
        );

    \I__12725\ : Odrv12
    port map (
            O => \N__52644\,
            I => \ADC_VDC.genclk.n6\
        );

    \I__12724\ : ClkMux
    port map (
            O => \N__52641\,
            I => \N__52635\
        );

    \I__12723\ : ClkMux
    port map (
            O => \N__52640\,
            I => \N__52632\
        );

    \I__12722\ : ClkMux
    port map (
            O => \N__52639\,
            I => \N__52629\
        );

    \I__12721\ : ClkMux
    port map (
            O => \N__52638\,
            I => \N__52623\
        );

    \I__12720\ : LocalMux
    port map (
            O => \N__52635\,
            I => \N__52620\
        );

    \I__12719\ : LocalMux
    port map (
            O => \N__52632\,
            I => \N__52617\
        );

    \I__12718\ : LocalMux
    port map (
            O => \N__52629\,
            I => \N__52614\
        );

    \I__12717\ : ClkMux
    port map (
            O => \N__52628\,
            I => \N__52611\
        );

    \I__12716\ : ClkMux
    port map (
            O => \N__52627\,
            I => \N__52606\
        );

    \I__12715\ : ClkMux
    port map (
            O => \N__52626\,
            I => \N__52603\
        );

    \I__12714\ : LocalMux
    port map (
            O => \N__52623\,
            I => \N__52598\
        );

    \I__12713\ : Span4Mux_v
    port map (
            O => \N__52620\,
            I => \N__52589\
        );

    \I__12712\ : Span4Mux_h
    port map (
            O => \N__52617\,
            I => \N__52589\
        );

    \I__12711\ : Span4Mux_v
    port map (
            O => \N__52614\,
            I => \N__52589\
        );

    \I__12710\ : LocalMux
    port map (
            O => \N__52611\,
            I => \N__52589\
        );

    \I__12709\ : ClkMux
    port map (
            O => \N__52610\,
            I => \N__52583\
        );

    \I__12708\ : ClkMux
    port map (
            O => \N__52609\,
            I => \N__52580\
        );

    \I__12707\ : LocalMux
    port map (
            O => \N__52606\,
            I => \N__52577\
        );

    \I__12706\ : LocalMux
    port map (
            O => \N__52603\,
            I => \N__52574\
        );

    \I__12705\ : ClkMux
    port map (
            O => \N__52602\,
            I => \N__52571\
        );

    \I__12704\ : ClkMux
    port map (
            O => \N__52601\,
            I => \N__52567\
        );

    \I__12703\ : Span4Mux_v
    port map (
            O => \N__52598\,
            I => \N__52562\
        );

    \I__12702\ : Span4Mux_v
    port map (
            O => \N__52589\,
            I => \N__52562\
        );

    \I__12701\ : ClkMux
    port map (
            O => \N__52588\,
            I => \N__52559\
        );

    \I__12700\ : ClkMux
    port map (
            O => \N__52587\,
            I => \N__52556\
        );

    \I__12699\ : ClkMux
    port map (
            O => \N__52586\,
            I => \N__52553\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__52583\,
            I => \N__52549\
        );

    \I__12697\ : LocalMux
    port map (
            O => \N__52580\,
            I => \N__52543\
        );

    \I__12696\ : Span4Mux_h
    port map (
            O => \N__52577\,
            I => \N__52538\
        );

    \I__12695\ : Span4Mux_v
    port map (
            O => \N__52574\,
            I => \N__52538\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__52571\,
            I => \N__52535\
        );

    \I__12693\ : ClkMux
    port map (
            O => \N__52570\,
            I => \N__52532\
        );

    \I__12692\ : LocalMux
    port map (
            O => \N__52567\,
            I => \N__52528\
        );

    \I__12691\ : Span4Mux_h
    port map (
            O => \N__52562\,
            I => \N__52523\
        );

    \I__12690\ : LocalMux
    port map (
            O => \N__52559\,
            I => \N__52523\
        );

    \I__12689\ : LocalMux
    port map (
            O => \N__52556\,
            I => \N__52518\
        );

    \I__12688\ : LocalMux
    port map (
            O => \N__52553\,
            I => \N__52518\
        );

    \I__12687\ : ClkMux
    port map (
            O => \N__52552\,
            I => \N__52515\
        );

    \I__12686\ : Span4Mux_h
    port map (
            O => \N__52549\,
            I => \N__52512\
        );

    \I__12685\ : ClkMux
    port map (
            O => \N__52548\,
            I => \N__52509\
        );

    \I__12684\ : ClkMux
    port map (
            O => \N__52547\,
            I => \N__52506\
        );

    \I__12683\ : ClkMux
    port map (
            O => \N__52546\,
            I => \N__52503\
        );

    \I__12682\ : Span4Mux_h
    port map (
            O => \N__52543\,
            I => \N__52499\
        );

    \I__12681\ : Span4Mux_h
    port map (
            O => \N__52538\,
            I => \N__52495\
        );

    \I__12680\ : Span4Mux_v
    port map (
            O => \N__52535\,
            I => \N__52490\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__52532\,
            I => \N__52490\
        );

    \I__12678\ : ClkMux
    port map (
            O => \N__52531\,
            I => \N__52487\
        );

    \I__12677\ : Span4Mux_h
    port map (
            O => \N__52528\,
            I => \N__52482\
        );

    \I__12676\ : Span4Mux_h
    port map (
            O => \N__52523\,
            I => \N__52482\
        );

    \I__12675\ : Span4Mux_v
    port map (
            O => \N__52518\,
            I => \N__52473\
        );

    \I__12674\ : LocalMux
    port map (
            O => \N__52515\,
            I => \N__52473\
        );

    \I__12673\ : Span4Mux_v
    port map (
            O => \N__52512\,
            I => \N__52473\
        );

    \I__12672\ : LocalMux
    port map (
            O => \N__52509\,
            I => \N__52473\
        );

    \I__12671\ : LocalMux
    port map (
            O => \N__52506\,
            I => \N__52468\
        );

    \I__12670\ : LocalMux
    port map (
            O => \N__52503\,
            I => \N__52468\
        );

    \I__12669\ : ClkMux
    port map (
            O => \N__52502\,
            I => \N__52465\
        );

    \I__12668\ : Span4Mux_h
    port map (
            O => \N__52499\,
            I => \N__52462\
        );

    \I__12667\ : ClkMux
    port map (
            O => \N__52498\,
            I => \N__52459\
        );

    \I__12666\ : Sp12to4
    port map (
            O => \N__52495\,
            I => \N__52452\
        );

    \I__12665\ : Sp12to4
    port map (
            O => \N__52490\,
            I => \N__52452\
        );

    \I__12664\ : LocalMux
    port map (
            O => \N__52487\,
            I => \N__52452\
        );

    \I__12663\ : Span4Mux_v
    port map (
            O => \N__52482\,
            I => \N__52449\
        );

    \I__12662\ : Span4Mux_h
    port map (
            O => \N__52473\,
            I => \N__52442\
        );

    \I__12661\ : Span4Mux_v
    port map (
            O => \N__52468\,
            I => \N__52442\
        );

    \I__12660\ : LocalMux
    port map (
            O => \N__52465\,
            I => \N__52442\
        );

    \I__12659\ : Span4Mux_v
    port map (
            O => \N__52462\,
            I => \N__52437\
        );

    \I__12658\ : LocalMux
    port map (
            O => \N__52459\,
            I => \N__52437\
        );

    \I__12657\ : Odrv12
    port map (
            O => \N__52452\,
            I => \comm_spi.iclk\
        );

    \I__12656\ : Odrv4
    port map (
            O => \N__52449\,
            I => \comm_spi.iclk\
        );

    \I__12655\ : Odrv4
    port map (
            O => \N__52442\,
            I => \comm_spi.iclk\
        );

    \I__12654\ : Odrv4
    port map (
            O => \N__52437\,
            I => \comm_spi.iclk\
        );

    \I__12653\ : InMux
    port map (
            O => \N__52428\,
            I => \N__52425\
        );

    \I__12652\ : LocalMux
    port map (
            O => \N__52425\,
            I => \N__52422\
        );

    \I__12651\ : Span4Mux_h
    port map (
            O => \N__52422\,
            I => \N__52419\
        );

    \I__12650\ : Odrv4
    port map (
            O => \N__52419\,
            I => n4_adj_1600
        );

    \I__12649\ : CascadeMux
    port map (
            O => \N__52416\,
            I => \n4_adj_1600_cascade_\
        );

    \I__12648\ : InMux
    port map (
            O => \N__52413\,
            I => \N__52401\
        );

    \I__12647\ : InMux
    port map (
            O => \N__52412\,
            I => \N__52398\
        );

    \I__12646\ : InMux
    port map (
            O => \N__52411\,
            I => \N__52395\
        );

    \I__12645\ : InMux
    port map (
            O => \N__52410\,
            I => \N__52392\
        );

    \I__12644\ : InMux
    port map (
            O => \N__52409\,
            I => \N__52389\
        );

    \I__12643\ : InMux
    port map (
            O => \N__52408\,
            I => \N__52383\
        );

    \I__12642\ : InMux
    port map (
            O => \N__52407\,
            I => \N__52374\
        );

    \I__12641\ : InMux
    port map (
            O => \N__52406\,
            I => \N__52374\
        );

    \I__12640\ : InMux
    port map (
            O => \N__52405\,
            I => \N__52374\
        );

    \I__12639\ : InMux
    port map (
            O => \N__52404\,
            I => \N__52374\
        );

    \I__12638\ : LocalMux
    port map (
            O => \N__52401\,
            I => \N__52371\
        );

    \I__12637\ : LocalMux
    port map (
            O => \N__52398\,
            I => \N__52367\
        );

    \I__12636\ : LocalMux
    port map (
            O => \N__52395\,
            I => \N__52362\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__52392\,
            I => \N__52362\
        );

    \I__12634\ : LocalMux
    port map (
            O => \N__52389\,
            I => \N__52359\
        );

    \I__12633\ : InMux
    port map (
            O => \N__52388\,
            I => \N__52356\
        );

    \I__12632\ : InMux
    port map (
            O => \N__52387\,
            I => \N__52351\
        );

    \I__12631\ : InMux
    port map (
            O => \N__52386\,
            I => \N__52348\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__52383\,
            I => \N__52339\
        );

    \I__12629\ : LocalMux
    port map (
            O => \N__52374\,
            I => \N__52339\
        );

    \I__12628\ : Span4Mux_v
    port map (
            O => \N__52371\,
            I => \N__52336\
        );

    \I__12627\ : InMux
    port map (
            O => \N__52370\,
            I => \N__52333\
        );

    \I__12626\ : Span4Mux_v
    port map (
            O => \N__52367\,
            I => \N__52321\
        );

    \I__12625\ : Span4Mux_v
    port map (
            O => \N__52362\,
            I => \N__52321\
        );

    \I__12624\ : Span4Mux_h
    port map (
            O => \N__52359\,
            I => \N__52321\
        );

    \I__12623\ : LocalMux
    port map (
            O => \N__52356\,
            I => \N__52321\
        );

    \I__12622\ : InMux
    port map (
            O => \N__52355\,
            I => \N__52316\
        );

    \I__12621\ : InMux
    port map (
            O => \N__52354\,
            I => \N__52316\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__52351\,
            I => \N__52311\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__52348\,
            I => \N__52311\
        );

    \I__12618\ : InMux
    port map (
            O => \N__52347\,
            I => \N__52302\
        );

    \I__12617\ : InMux
    port map (
            O => \N__52346\,
            I => \N__52302\
        );

    \I__12616\ : InMux
    port map (
            O => \N__52345\,
            I => \N__52302\
        );

    \I__12615\ : InMux
    port map (
            O => \N__52344\,
            I => \N__52302\
        );

    \I__12614\ : Span4Mux_h
    port map (
            O => \N__52339\,
            I => \N__52299\
        );

    \I__12613\ : Span4Mux_v
    port map (
            O => \N__52336\,
            I => \N__52294\
        );

    \I__12612\ : LocalMux
    port map (
            O => \N__52333\,
            I => \N__52294\
        );

    \I__12611\ : InMux
    port map (
            O => \N__52332\,
            I => \N__52287\
        );

    \I__12610\ : InMux
    port map (
            O => \N__52331\,
            I => \N__52287\
        );

    \I__12609\ : InMux
    port map (
            O => \N__52330\,
            I => \N__52287\
        );

    \I__12608\ : Span4Mux_h
    port map (
            O => \N__52321\,
            I => \N__52284\
        );

    \I__12607\ : LocalMux
    port map (
            O => \N__52316\,
            I => comm_index_1
        );

    \I__12606\ : Odrv4
    port map (
            O => \N__52311\,
            I => comm_index_1
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__52302\,
            I => comm_index_1
        );

    \I__12604\ : Odrv4
    port map (
            O => \N__52299\,
            I => comm_index_1
        );

    \I__12603\ : Odrv4
    port map (
            O => \N__52294\,
            I => comm_index_1
        );

    \I__12602\ : LocalMux
    port map (
            O => \N__52287\,
            I => comm_index_1
        );

    \I__12601\ : Odrv4
    port map (
            O => \N__52284\,
            I => comm_index_1
        );

    \I__12600\ : CascadeMux
    port map (
            O => \N__52269\,
            I => \n5_cascade_\
        );

    \I__12599\ : InMux
    port map (
            O => \N__52266\,
            I => \N__52262\
        );

    \I__12598\ : InMux
    port map (
            O => \N__52265\,
            I => \N__52259\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__52262\,
            I => \N__52255\
        );

    \I__12596\ : LocalMux
    port map (
            O => \N__52259\,
            I => \N__52251\
        );

    \I__12595\ : InMux
    port map (
            O => \N__52258\,
            I => \N__52248\
        );

    \I__12594\ : Span4Mux_h
    port map (
            O => \N__52255\,
            I => \N__52245\
        );

    \I__12593\ : InMux
    port map (
            O => \N__52254\,
            I => \N__52240\
        );

    \I__12592\ : Span4Mux_h
    port map (
            O => \N__52251\,
            I => \N__52237\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__52248\,
            I => \N__52234\
        );

    \I__12590\ : Span4Mux_h
    port map (
            O => \N__52245\,
            I => \N__52231\
        );

    \I__12589\ : InMux
    port map (
            O => \N__52244\,
            I => \N__52228\
        );

    \I__12588\ : InMux
    port map (
            O => \N__52243\,
            I => \N__52225\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__52240\,
            I => comm_cmd_7
        );

    \I__12586\ : Odrv4
    port map (
            O => \N__52237\,
            I => comm_cmd_7
        );

    \I__12585\ : Odrv4
    port map (
            O => \N__52234\,
            I => comm_cmd_7
        );

    \I__12584\ : Odrv4
    port map (
            O => \N__52231\,
            I => comm_cmd_7
        );

    \I__12583\ : LocalMux
    port map (
            O => \N__52228\,
            I => comm_cmd_7
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__52225\,
            I => comm_cmd_7
        );

    \I__12581\ : InMux
    port map (
            O => \N__52212\,
            I => \N__52209\
        );

    \I__12580\ : LocalMux
    port map (
            O => \N__52209\,
            I => \N__52206\
        );

    \I__12579\ : Span4Mux_h
    port map (
            O => \N__52206\,
            I => \N__52203\
        );

    \I__12578\ : Span4Mux_h
    port map (
            O => \N__52203\,
            I => \N__52200\
        );

    \I__12577\ : Odrv4
    port map (
            O => \N__52200\,
            I => n21888
        );

    \I__12576\ : CascadeMux
    port map (
            O => \N__52197\,
            I => \N__52194\
        );

    \I__12575\ : InMux
    port map (
            O => \N__52194\,
            I => \N__52191\
        );

    \I__12574\ : LocalMux
    port map (
            O => \N__52191\,
            I => n21317
        );

    \I__12573\ : InMux
    port map (
            O => \N__52188\,
            I => \N__52184\
        );

    \I__12572\ : InMux
    port map (
            O => \N__52187\,
            I => \N__52181\
        );

    \I__12571\ : LocalMux
    port map (
            O => \N__52184\,
            I => \N__52178\
        );

    \I__12570\ : LocalMux
    port map (
            O => \N__52181\,
            I => \N__52174\
        );

    \I__12569\ : Span4Mux_v
    port map (
            O => \N__52178\,
            I => \N__52171\
        );

    \I__12568\ : CascadeMux
    port map (
            O => \N__52177\,
            I => \N__52168\
        );

    \I__12567\ : Span12Mux_v
    port map (
            O => \N__52174\,
            I => \N__52165\
        );

    \I__12566\ : Sp12to4
    port map (
            O => \N__52171\,
            I => \N__52162\
        );

    \I__12565\ : InMux
    port map (
            O => \N__52168\,
            I => \N__52159\
        );

    \I__12564\ : Span12Mux_h
    port map (
            O => \N__52165\,
            I => \N__52156\
        );

    \I__12563\ : Span12Mux_h
    port map (
            O => \N__52162\,
            I => \N__52153\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__52159\,
            I => buf_adcdata_iac_15
        );

    \I__12561\ : Odrv12
    port map (
            O => \N__52156\,
            I => buf_adcdata_iac_15
        );

    \I__12560\ : Odrv12
    port map (
            O => \N__52153\,
            I => buf_adcdata_iac_15
        );

    \I__12559\ : InMux
    port map (
            O => \N__52146\,
            I => \N__52143\
        );

    \I__12558\ : LocalMux
    port map (
            O => \N__52143\,
            I => \N__52140\
        );

    \I__12557\ : Sp12to4
    port map (
            O => \N__52140\,
            I => \N__52137\
        );

    \I__12556\ : Odrv12
    port map (
            O => \N__52137\,
            I => n16_adj_1504
        );

    \I__12555\ : InMux
    port map (
            O => \N__52134\,
            I => \N__52131\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__52131\,
            I => \N__52128\
        );

    \I__12553\ : Odrv4
    port map (
            O => \N__52128\,
            I => n21048
        );

    \I__12552\ : CascadeMux
    port map (
            O => \N__52125\,
            I => \N__52121\
        );

    \I__12551\ : InMux
    port map (
            O => \N__52124\,
            I => \N__52118\
        );

    \I__12550\ : InMux
    port map (
            O => \N__52121\,
            I => \N__52114\
        );

    \I__12549\ : LocalMux
    port map (
            O => \N__52118\,
            I => \N__52108\
        );

    \I__12548\ : InMux
    port map (
            O => \N__52117\,
            I => \N__52105\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__52114\,
            I => \N__52102\
        );

    \I__12546\ : InMux
    port map (
            O => \N__52113\,
            I => \N__52099\
        );

    \I__12545\ : InMux
    port map (
            O => \N__52112\,
            I => \N__52096\
        );

    \I__12544\ : InMux
    port map (
            O => \N__52111\,
            I => \N__52093\
        );

    \I__12543\ : Span4Mux_h
    port map (
            O => \N__52108\,
            I => \N__52087\
        );

    \I__12542\ : LocalMux
    port map (
            O => \N__52105\,
            I => \N__52087\
        );

    \I__12541\ : Span4Mux_h
    port map (
            O => \N__52102\,
            I => \N__52084\
        );

    \I__12540\ : LocalMux
    port map (
            O => \N__52099\,
            I => \N__52079\
        );

    \I__12539\ : LocalMux
    port map (
            O => \N__52096\,
            I => \N__52079\
        );

    \I__12538\ : LocalMux
    port map (
            O => \N__52093\,
            I => \N__52076\
        );

    \I__12537\ : InMux
    port map (
            O => \N__52092\,
            I => \N__52073\
        );

    \I__12536\ : Sp12to4
    port map (
            O => \N__52087\,
            I => \N__52066\
        );

    \I__12535\ : Sp12to4
    port map (
            O => \N__52084\,
            I => \N__52066\
        );

    \I__12534\ : Sp12to4
    port map (
            O => \N__52079\,
            I => \N__52066\
        );

    \I__12533\ : Span4Mux_v
    port map (
            O => \N__52076\,
            I => \N__52063\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__52073\,
            I => \N__52060\
        );

    \I__12531\ : Span12Mux_v
    port map (
            O => \N__52066\,
            I => \N__52055\
        );

    \I__12530\ : Span4Mux_h
    port map (
            O => \N__52063\,
            I => \N__52052\
        );

    \I__12529\ : Span4Mux_v
    port map (
            O => \N__52060\,
            I => \N__52049\
        );

    \I__12528\ : InMux
    port map (
            O => \N__52059\,
            I => \N__52046\
        );

    \I__12527\ : InMux
    port map (
            O => \N__52058\,
            I => \N__52043\
        );

    \I__12526\ : Odrv12
    port map (
            O => \N__52055\,
            I => comm_rx_buf_5
        );

    \I__12525\ : Odrv4
    port map (
            O => \N__52052\,
            I => comm_rx_buf_5
        );

    \I__12524\ : Odrv4
    port map (
            O => \N__52049\,
            I => comm_rx_buf_5
        );

    \I__12523\ : LocalMux
    port map (
            O => \N__52046\,
            I => comm_rx_buf_5
        );

    \I__12522\ : LocalMux
    port map (
            O => \N__52043\,
            I => comm_rx_buf_5
        );

    \I__12521\ : InMux
    port map (
            O => \N__52032\,
            I => \N__52029\
        );

    \I__12520\ : LocalMux
    port map (
            O => \N__52029\,
            I => \N__52023\
        );

    \I__12519\ : InMux
    port map (
            O => \N__52028\,
            I => \N__52004\
        );

    \I__12518\ : InMux
    port map (
            O => \N__52027\,
            I => \N__52001\
        );

    \I__12517\ : InMux
    port map (
            O => \N__52026\,
            I => \N__51989\
        );

    \I__12516\ : Span4Mux_v
    port map (
            O => \N__52023\,
            I => \N__51986\
        );

    \I__12515\ : InMux
    port map (
            O => \N__52022\,
            I => \N__51983\
        );

    \I__12514\ : InMux
    port map (
            O => \N__52021\,
            I => \N__51978\
        );

    \I__12513\ : InMux
    port map (
            O => \N__52020\,
            I => \N__51978\
        );

    \I__12512\ : InMux
    port map (
            O => \N__52019\,
            I => \N__51961\
        );

    \I__12511\ : InMux
    port map (
            O => \N__52018\,
            I => \N__51961\
        );

    \I__12510\ : InMux
    port map (
            O => \N__52017\,
            I => \N__51961\
        );

    \I__12509\ : InMux
    port map (
            O => \N__52016\,
            I => \N__51961\
        );

    \I__12508\ : InMux
    port map (
            O => \N__52015\,
            I => \N__51961\
        );

    \I__12507\ : InMux
    port map (
            O => \N__52014\,
            I => \N__51961\
        );

    \I__12506\ : InMux
    port map (
            O => \N__52013\,
            I => \N__51961\
        );

    \I__12505\ : InMux
    port map (
            O => \N__52012\,
            I => \N__51961\
        );

    \I__12504\ : InMux
    port map (
            O => \N__52011\,
            I => \N__51951\
        );

    \I__12503\ : InMux
    port map (
            O => \N__52010\,
            I => \N__51951\
        );

    \I__12502\ : InMux
    port map (
            O => \N__52009\,
            I => \N__51951\
        );

    \I__12501\ : InMux
    port map (
            O => \N__52008\,
            I => \N__51940\
        );

    \I__12500\ : InMux
    port map (
            O => \N__52007\,
            I => \N__51937\
        );

    \I__12499\ : LocalMux
    port map (
            O => \N__52004\,
            I => \N__51932\
        );

    \I__12498\ : LocalMux
    port map (
            O => \N__52001\,
            I => \N__51932\
        );

    \I__12497\ : InMux
    port map (
            O => \N__52000\,
            I => \N__51929\
        );

    \I__12496\ : InMux
    port map (
            O => \N__51999\,
            I => \N__51926\
        );

    \I__12495\ : InMux
    port map (
            O => \N__51998\,
            I => \N__51921\
        );

    \I__12494\ : InMux
    port map (
            O => \N__51997\,
            I => \N__51918\
        );

    \I__12493\ : CascadeMux
    port map (
            O => \N__51996\,
            I => \N__51913\
        );

    \I__12492\ : CascadeMux
    port map (
            O => \N__51995\,
            I => \N__51910\
        );

    \I__12491\ : InMux
    port map (
            O => \N__51994\,
            I => \N__51906\
        );

    \I__12490\ : InMux
    port map (
            O => \N__51993\,
            I => \N__51901\
        );

    \I__12489\ : InMux
    port map (
            O => \N__51992\,
            I => \N__51898\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__51989\,
            I => \N__51887\
        );

    \I__12487\ : Span4Mux_h
    port map (
            O => \N__51986\,
            I => \N__51887\
        );

    \I__12486\ : LocalMux
    port map (
            O => \N__51983\,
            I => \N__51887\
        );

    \I__12485\ : LocalMux
    port map (
            O => \N__51978\,
            I => \N__51887\
        );

    \I__12484\ : LocalMux
    port map (
            O => \N__51961\,
            I => \N__51887\
        );

    \I__12483\ : InMux
    port map (
            O => \N__51960\,
            I => \N__51884\
        );

    \I__12482\ : InMux
    port map (
            O => \N__51959\,
            I => \N__51881\
        );

    \I__12481\ : CascadeMux
    port map (
            O => \N__51958\,
            I => \N__51873\
        );

    \I__12480\ : LocalMux
    port map (
            O => \N__51951\,
            I => \N__51855\
        );

    \I__12479\ : InMux
    port map (
            O => \N__51950\,
            I => \N__51838\
        );

    \I__12478\ : InMux
    port map (
            O => \N__51949\,
            I => \N__51838\
        );

    \I__12477\ : InMux
    port map (
            O => \N__51948\,
            I => \N__51838\
        );

    \I__12476\ : InMux
    port map (
            O => \N__51947\,
            I => \N__51838\
        );

    \I__12475\ : InMux
    port map (
            O => \N__51946\,
            I => \N__51838\
        );

    \I__12474\ : InMux
    port map (
            O => \N__51945\,
            I => \N__51838\
        );

    \I__12473\ : InMux
    port map (
            O => \N__51944\,
            I => \N__51838\
        );

    \I__12472\ : InMux
    port map (
            O => \N__51943\,
            I => \N__51838\
        );

    \I__12471\ : LocalMux
    port map (
            O => \N__51940\,
            I => \N__51827\
        );

    \I__12470\ : LocalMux
    port map (
            O => \N__51937\,
            I => \N__51827\
        );

    \I__12469\ : Span4Mux_v
    port map (
            O => \N__51932\,
            I => \N__51827\
        );

    \I__12468\ : LocalMux
    port map (
            O => \N__51929\,
            I => \N__51827\
        );

    \I__12467\ : LocalMux
    port map (
            O => \N__51926\,
            I => \N__51827\
        );

    \I__12466\ : InMux
    port map (
            O => \N__51925\,
            I => \N__51821\
        );

    \I__12465\ : InMux
    port map (
            O => \N__51924\,
            I => \N__51818\
        );

    \I__12464\ : LocalMux
    port map (
            O => \N__51921\,
            I => \N__51813\
        );

    \I__12463\ : LocalMux
    port map (
            O => \N__51918\,
            I => \N__51813\
        );

    \I__12462\ : InMux
    port map (
            O => \N__51917\,
            I => \N__51808\
        );

    \I__12461\ : InMux
    port map (
            O => \N__51916\,
            I => \N__51808\
        );

    \I__12460\ : InMux
    port map (
            O => \N__51913\,
            I => \N__51801\
        );

    \I__12459\ : InMux
    port map (
            O => \N__51910\,
            I => \N__51801\
        );

    \I__12458\ : InMux
    port map (
            O => \N__51909\,
            I => \N__51801\
        );

    \I__12457\ : LocalMux
    port map (
            O => \N__51906\,
            I => \N__51796\
        );

    \I__12456\ : InMux
    port map (
            O => \N__51905\,
            I => \N__51793\
        );

    \I__12455\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51789\
        );

    \I__12454\ : LocalMux
    port map (
            O => \N__51901\,
            I => \N__51778\
        );

    \I__12453\ : LocalMux
    port map (
            O => \N__51898\,
            I => \N__51778\
        );

    \I__12452\ : Span4Mux_v
    port map (
            O => \N__51887\,
            I => \N__51778\
        );

    \I__12451\ : LocalMux
    port map (
            O => \N__51884\,
            I => \N__51778\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__51881\,
            I => \N__51778\
        );

    \I__12449\ : InMux
    port map (
            O => \N__51880\,
            I => \N__51775\
        );

    \I__12448\ : InMux
    port map (
            O => \N__51879\,
            I => \N__51772\
        );

    \I__12447\ : InMux
    port map (
            O => \N__51878\,
            I => \N__51769\
        );

    \I__12446\ : InMux
    port map (
            O => \N__51877\,
            I => \N__51762\
        );

    \I__12445\ : InMux
    port map (
            O => \N__51876\,
            I => \N__51762\
        );

    \I__12444\ : InMux
    port map (
            O => \N__51873\,
            I => \N__51762\
        );

    \I__12443\ : InMux
    port map (
            O => \N__51872\,
            I => \N__51755\
        );

    \I__12442\ : InMux
    port map (
            O => \N__51871\,
            I => \N__51740\
        );

    \I__12441\ : InMux
    port map (
            O => \N__51870\,
            I => \N__51740\
        );

    \I__12440\ : InMux
    port map (
            O => \N__51869\,
            I => \N__51740\
        );

    \I__12439\ : InMux
    port map (
            O => \N__51868\,
            I => \N__51740\
        );

    \I__12438\ : InMux
    port map (
            O => \N__51867\,
            I => \N__51740\
        );

    \I__12437\ : InMux
    port map (
            O => \N__51866\,
            I => \N__51740\
        );

    \I__12436\ : InMux
    port map (
            O => \N__51865\,
            I => \N__51740\
        );

    \I__12435\ : InMux
    port map (
            O => \N__51864\,
            I => \N__51731\
        );

    \I__12434\ : InMux
    port map (
            O => \N__51863\,
            I => \N__51731\
        );

    \I__12433\ : InMux
    port map (
            O => \N__51862\,
            I => \N__51731\
        );

    \I__12432\ : InMux
    port map (
            O => \N__51861\,
            I => \N__51731\
        );

    \I__12431\ : InMux
    port map (
            O => \N__51860\,
            I => \N__51728\
        );

    \I__12430\ : CascadeMux
    port map (
            O => \N__51859\,
            I => \N__51715\
        );

    \I__12429\ : InMux
    port map (
            O => \N__51858\,
            I => \N__51711\
        );

    \I__12428\ : Span4Mux_v
    port map (
            O => \N__51855\,
            I => \N__51708\
        );

    \I__12427\ : LocalMux
    port map (
            O => \N__51838\,
            I => \N__51703\
        );

    \I__12426\ : Span4Mux_v
    port map (
            O => \N__51827\,
            I => \N__51703\
        );

    \I__12425\ : InMux
    port map (
            O => \N__51826\,
            I => \N__51696\
        );

    \I__12424\ : InMux
    port map (
            O => \N__51825\,
            I => \N__51696\
        );

    \I__12423\ : InMux
    port map (
            O => \N__51824\,
            I => \N__51696\
        );

    \I__12422\ : LocalMux
    port map (
            O => \N__51821\,
            I => \N__51685\
        );

    \I__12421\ : LocalMux
    port map (
            O => \N__51818\,
            I => \N__51685\
        );

    \I__12420\ : Span4Mux_v
    port map (
            O => \N__51813\,
            I => \N__51685\
        );

    \I__12419\ : LocalMux
    port map (
            O => \N__51808\,
            I => \N__51685\
        );

    \I__12418\ : LocalMux
    port map (
            O => \N__51801\,
            I => \N__51685\
        );

    \I__12417\ : InMux
    port map (
            O => \N__51800\,
            I => \N__51682\
        );

    \I__12416\ : InMux
    port map (
            O => \N__51799\,
            I => \N__51679\
        );

    \I__12415\ : Span4Mux_v
    port map (
            O => \N__51796\,
            I => \N__51674\
        );

    \I__12414\ : LocalMux
    port map (
            O => \N__51793\,
            I => \N__51674\
        );

    \I__12413\ : InMux
    port map (
            O => \N__51792\,
            I => \N__51671\
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__51789\,
            I => \N__51666\
        );

    \I__12411\ : Span4Mux_v
    port map (
            O => \N__51778\,
            I => \N__51666\
        );

    \I__12410\ : LocalMux
    port map (
            O => \N__51775\,
            I => \N__51657\
        );

    \I__12409\ : LocalMux
    port map (
            O => \N__51772\,
            I => \N__51657\
        );

    \I__12408\ : LocalMux
    port map (
            O => \N__51769\,
            I => \N__51657\
        );

    \I__12407\ : LocalMux
    port map (
            O => \N__51762\,
            I => \N__51657\
        );

    \I__12406\ : InMux
    port map (
            O => \N__51761\,
            I => \N__51646\
        );

    \I__12405\ : CascadeMux
    port map (
            O => \N__51760\,
            I => \N__51638\
        );

    \I__12404\ : CascadeMux
    port map (
            O => \N__51759\,
            I => \N__51633\
        );

    \I__12403\ : InMux
    port map (
            O => \N__51758\,
            I => \N__51629\
        );

    \I__12402\ : LocalMux
    port map (
            O => \N__51755\,
            I => \N__51626\
        );

    \I__12401\ : LocalMux
    port map (
            O => \N__51740\,
            I => \N__51623\
        );

    \I__12400\ : LocalMux
    port map (
            O => \N__51731\,
            I => \N__51620\
        );

    \I__12399\ : LocalMux
    port map (
            O => \N__51728\,
            I => \N__51617\
        );

    \I__12398\ : InMux
    port map (
            O => \N__51727\,
            I => \N__51614\
        );

    \I__12397\ : InMux
    port map (
            O => \N__51726\,
            I => \N__51611\
        );

    \I__12396\ : InMux
    port map (
            O => \N__51725\,
            I => \N__51604\
        );

    \I__12395\ : InMux
    port map (
            O => \N__51724\,
            I => \N__51604\
        );

    \I__12394\ : InMux
    port map (
            O => \N__51723\,
            I => \N__51604\
        );

    \I__12393\ : InMux
    port map (
            O => \N__51722\,
            I => \N__51599\
        );

    \I__12392\ : InMux
    port map (
            O => \N__51721\,
            I => \N__51599\
        );

    \I__12391\ : InMux
    port map (
            O => \N__51720\,
            I => \N__51596\
        );

    \I__12390\ : InMux
    port map (
            O => \N__51719\,
            I => \N__51587\
        );

    \I__12389\ : InMux
    port map (
            O => \N__51718\,
            I => \N__51587\
        );

    \I__12388\ : InMux
    port map (
            O => \N__51715\,
            I => \N__51587\
        );

    \I__12387\ : InMux
    port map (
            O => \N__51714\,
            I => \N__51587\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__51711\,
            I => \N__51578\
        );

    \I__12385\ : Span4Mux_h
    port map (
            O => \N__51708\,
            I => \N__51578\
        );

    \I__12384\ : Span4Mux_h
    port map (
            O => \N__51703\,
            I => \N__51578\
        );

    \I__12383\ : LocalMux
    port map (
            O => \N__51696\,
            I => \N__51578\
        );

    \I__12382\ : Span4Mux_v
    port map (
            O => \N__51685\,
            I => \N__51575\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__51682\,
            I => \N__51569\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__51679\,
            I => \N__51566\
        );

    \I__12379\ : Span4Mux_v
    port map (
            O => \N__51674\,
            I => \N__51563\
        );

    \I__12378\ : LocalMux
    port map (
            O => \N__51671\,
            I => \N__51556\
        );

    \I__12377\ : Span4Mux_h
    port map (
            O => \N__51666\,
            I => \N__51556\
        );

    \I__12376\ : Span4Mux_v
    port map (
            O => \N__51657\,
            I => \N__51556\
        );

    \I__12375\ : InMux
    port map (
            O => \N__51656\,
            I => \N__51539\
        );

    \I__12374\ : InMux
    port map (
            O => \N__51655\,
            I => \N__51539\
        );

    \I__12373\ : InMux
    port map (
            O => \N__51654\,
            I => \N__51539\
        );

    \I__12372\ : InMux
    port map (
            O => \N__51653\,
            I => \N__51539\
        );

    \I__12371\ : InMux
    port map (
            O => \N__51652\,
            I => \N__51539\
        );

    \I__12370\ : InMux
    port map (
            O => \N__51651\,
            I => \N__51539\
        );

    \I__12369\ : InMux
    port map (
            O => \N__51650\,
            I => \N__51539\
        );

    \I__12368\ : InMux
    port map (
            O => \N__51649\,
            I => \N__51539\
        );

    \I__12367\ : LocalMux
    port map (
            O => \N__51646\,
            I => \N__51536\
        );

    \I__12366\ : InMux
    port map (
            O => \N__51645\,
            I => \N__51533\
        );

    \I__12365\ : InMux
    port map (
            O => \N__51644\,
            I => \N__51526\
        );

    \I__12364\ : InMux
    port map (
            O => \N__51643\,
            I => \N__51526\
        );

    \I__12363\ : InMux
    port map (
            O => \N__51642\,
            I => \N__51526\
        );

    \I__12362\ : InMux
    port map (
            O => \N__51641\,
            I => \N__51519\
        );

    \I__12361\ : InMux
    port map (
            O => \N__51638\,
            I => \N__51519\
        );

    \I__12360\ : InMux
    port map (
            O => \N__51637\,
            I => \N__51519\
        );

    \I__12359\ : InMux
    port map (
            O => \N__51636\,
            I => \N__51512\
        );

    \I__12358\ : InMux
    port map (
            O => \N__51633\,
            I => \N__51512\
        );

    \I__12357\ : InMux
    port map (
            O => \N__51632\,
            I => \N__51512\
        );

    \I__12356\ : LocalMux
    port map (
            O => \N__51629\,
            I => \N__51503\
        );

    \I__12355\ : Span4Mux_h
    port map (
            O => \N__51626\,
            I => \N__51503\
        );

    \I__12354\ : Span4Mux_h
    port map (
            O => \N__51623\,
            I => \N__51503\
        );

    \I__12353\ : Span4Mux_v
    port map (
            O => \N__51620\,
            I => \N__51503\
        );

    \I__12352\ : Span12Mux_v
    port map (
            O => \N__51617\,
            I => \N__51496\
        );

    \I__12351\ : LocalMux
    port map (
            O => \N__51614\,
            I => \N__51496\
        );

    \I__12350\ : LocalMux
    port map (
            O => \N__51611\,
            I => \N__51496\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__51604\,
            I => \N__51491\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__51599\,
            I => \N__51491\
        );

    \I__12347\ : LocalMux
    port map (
            O => \N__51596\,
            I => \N__51486\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__51587\,
            I => \N__51486\
        );

    \I__12345\ : Span4Mux_v
    port map (
            O => \N__51578\,
            I => \N__51481\
        );

    \I__12344\ : Span4Mux_h
    port map (
            O => \N__51575\,
            I => \N__51481\
        );

    \I__12343\ : InMux
    port map (
            O => \N__51574\,
            I => \N__51474\
        );

    \I__12342\ : InMux
    port map (
            O => \N__51573\,
            I => \N__51474\
        );

    \I__12341\ : InMux
    port map (
            O => \N__51572\,
            I => \N__51474\
        );

    \I__12340\ : Span4Mux_v
    port map (
            O => \N__51569\,
            I => \N__51465\
        );

    \I__12339\ : Span4Mux_v
    port map (
            O => \N__51566\,
            I => \N__51465\
        );

    \I__12338\ : Span4Mux_h
    port map (
            O => \N__51563\,
            I => \N__51465\
        );

    \I__12337\ : Span4Mux_v
    port map (
            O => \N__51556\,
            I => \N__51465\
        );

    \I__12336\ : LocalMux
    port map (
            O => \N__51539\,
            I => comm_state_1
        );

    \I__12335\ : Odrv4
    port map (
            O => \N__51536\,
            I => comm_state_1
        );

    \I__12334\ : LocalMux
    port map (
            O => \N__51533\,
            I => comm_state_1
        );

    \I__12333\ : LocalMux
    port map (
            O => \N__51526\,
            I => comm_state_1
        );

    \I__12332\ : LocalMux
    port map (
            O => \N__51519\,
            I => comm_state_1
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__51512\,
            I => comm_state_1
        );

    \I__12330\ : Odrv4
    port map (
            O => \N__51503\,
            I => comm_state_1
        );

    \I__12329\ : Odrv12
    port map (
            O => \N__51496\,
            I => comm_state_1
        );

    \I__12328\ : Odrv12
    port map (
            O => \N__51491\,
            I => comm_state_1
        );

    \I__12327\ : Odrv4
    port map (
            O => \N__51486\,
            I => comm_state_1
        );

    \I__12326\ : Odrv4
    port map (
            O => \N__51481\,
            I => comm_state_1
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__51474\,
            I => comm_state_1
        );

    \I__12324\ : Odrv4
    port map (
            O => \N__51465\,
            I => comm_state_1
        );

    \I__12323\ : InMux
    port map (
            O => \N__51438\,
            I => \N__51432\
        );

    \I__12322\ : InMux
    port map (
            O => \N__51437\,
            I => \N__51429\
        );

    \I__12321\ : InMux
    port map (
            O => \N__51436\,
            I => \N__51425\
        );

    \I__12320\ : InMux
    port map (
            O => \N__51435\,
            I => \N__51422\
        );

    \I__12319\ : LocalMux
    port map (
            O => \N__51432\,
            I => \N__51419\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__51429\,
            I => \N__51416\
        );

    \I__12317\ : InMux
    port map (
            O => \N__51428\,
            I => \N__51413\
        );

    \I__12316\ : LocalMux
    port map (
            O => \N__51425\,
            I => \N__51410\
        );

    \I__12315\ : LocalMux
    port map (
            O => \N__51422\,
            I => \N__51407\
        );

    \I__12314\ : Span4Mux_v
    port map (
            O => \N__51419\,
            I => \N__51400\
        );

    \I__12313\ : Span4Mux_h
    port map (
            O => \N__51416\,
            I => \N__51400\
        );

    \I__12312\ : LocalMux
    port map (
            O => \N__51413\,
            I => \N__51400\
        );

    \I__12311\ : Span4Mux_v
    port map (
            O => \N__51410\,
            I => \N__51397\
        );

    \I__12310\ : Span12Mux_v
    port map (
            O => \N__51407\,
            I => \N__51394\
        );

    \I__12309\ : Span4Mux_h
    port map (
            O => \N__51400\,
            I => \N__51389\
        );

    \I__12308\ : Span4Mux_v
    port map (
            O => \N__51397\,
            I => \N__51389\
        );

    \I__12307\ : Odrv12
    port map (
            O => \N__51394\,
            I => comm_buf_1_5
        );

    \I__12306\ : Odrv4
    port map (
            O => \N__51389\,
            I => comm_buf_1_5
        );

    \I__12305\ : CEMux
    port map (
            O => \N__51384\,
            I => \N__51378\
        );

    \I__12304\ : CEMux
    port map (
            O => \N__51383\,
            I => \N__51375\
        );

    \I__12303\ : CEMux
    port map (
            O => \N__51382\,
            I => \N__51371\
        );

    \I__12302\ : CEMux
    port map (
            O => \N__51381\,
            I => \N__51368\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__51378\,
            I => \N__51365\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__51375\,
            I => \N__51362\
        );

    \I__12299\ : CEMux
    port map (
            O => \N__51374\,
            I => \N__51359\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__51371\,
            I => \N__51353\
        );

    \I__12297\ : LocalMux
    port map (
            O => \N__51368\,
            I => \N__51350\
        );

    \I__12296\ : Span4Mux_h
    port map (
            O => \N__51365\,
            I => \N__51347\
        );

    \I__12295\ : Span4Mux_h
    port map (
            O => \N__51362\,
            I => \N__51342\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__51359\,
            I => \N__51342\
        );

    \I__12293\ : CEMux
    port map (
            O => \N__51358\,
            I => \N__51339\
        );

    \I__12292\ : CEMux
    port map (
            O => \N__51357\,
            I => \N__51336\
        );

    \I__12291\ : CEMux
    port map (
            O => \N__51356\,
            I => \N__51333\
        );

    \I__12290\ : Span4Mux_h
    port map (
            O => \N__51353\,
            I => \N__51330\
        );

    \I__12289\ : Span4Mux_v
    port map (
            O => \N__51350\,
            I => \N__51327\
        );

    \I__12288\ : Sp12to4
    port map (
            O => \N__51347\,
            I => \N__51324\
        );

    \I__12287\ : Span4Mux_v
    port map (
            O => \N__51342\,
            I => \N__51321\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__51339\,
            I => n11991
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__51336\,
            I => n11991
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__51333\,
            I => n11991
        );

    \I__12283\ : Odrv4
    port map (
            O => \N__51330\,
            I => n11991
        );

    \I__12282\ : Odrv4
    port map (
            O => \N__51327\,
            I => n11991
        );

    \I__12281\ : Odrv12
    port map (
            O => \N__51324\,
            I => n11991
        );

    \I__12280\ : Odrv4
    port map (
            O => \N__51321\,
            I => n11991
        );

    \I__12279\ : SRMux
    port map (
            O => \N__51306\,
            I => \N__51303\
        );

    \I__12278\ : LocalMux
    port map (
            O => \N__51303\,
            I => \N__51296\
        );

    \I__12277\ : SRMux
    port map (
            O => \N__51302\,
            I => \N__51293\
        );

    \I__12276\ : SRMux
    port map (
            O => \N__51301\,
            I => \N__51290\
        );

    \I__12275\ : SRMux
    port map (
            O => \N__51300\,
            I => \N__51287\
        );

    \I__12274\ : SRMux
    port map (
            O => \N__51299\,
            I => \N__51284\
        );

    \I__12273\ : Span4Mux_h
    port map (
            O => \N__51296\,
            I => \N__51278\
        );

    \I__12272\ : LocalMux
    port map (
            O => \N__51293\,
            I => \N__51278\
        );

    \I__12271\ : LocalMux
    port map (
            O => \N__51290\,
            I => \N__51270\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__51287\,
            I => \N__51270\
        );

    \I__12269\ : LocalMux
    port map (
            O => \N__51284\,
            I => \N__51270\
        );

    \I__12268\ : SRMux
    port map (
            O => \N__51283\,
            I => \N__51267\
        );

    \I__12267\ : Span4Mux_h
    port map (
            O => \N__51278\,
            I => \N__51264\
        );

    \I__12266\ : SRMux
    port map (
            O => \N__51277\,
            I => \N__51261\
        );

    \I__12265\ : Span4Mux_v
    port map (
            O => \N__51270\,
            I => \N__51258\
        );

    \I__12264\ : LocalMux
    port map (
            O => \N__51267\,
            I => \N__51250\
        );

    \I__12263\ : Span4Mux_h
    port map (
            O => \N__51264\,
            I => \N__51250\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__51261\,
            I => \N__51250\
        );

    \I__12261\ : Span4Mux_h
    port map (
            O => \N__51258\,
            I => \N__51247\
        );

    \I__12260\ : SRMux
    port map (
            O => \N__51257\,
            I => \N__51244\
        );

    \I__12259\ : Span4Mux_v
    port map (
            O => \N__51250\,
            I => \N__51241\
        );

    \I__12258\ : Sp12to4
    port map (
            O => \N__51247\,
            I => \N__51238\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__51244\,
            I => \N__51233\
        );

    \I__12256\ : Sp12to4
    port map (
            O => \N__51241\,
            I => \N__51233\
        );

    \I__12255\ : Odrv12
    port map (
            O => \N__51238\,
            I => n14757
        );

    \I__12254\ : Odrv12
    port map (
            O => \N__51233\,
            I => n14757
        );

    \I__12253\ : InMux
    port map (
            O => \N__51228\,
            I => \N__51225\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__51225\,
            I => \N__51222\
        );

    \I__12251\ : Span4Mux_v
    port map (
            O => \N__51222\,
            I => \N__51219\
        );

    \I__12250\ : Span4Mux_h
    port map (
            O => \N__51219\,
            I => \N__51216\
        );

    \I__12249\ : Span4Mux_h
    port map (
            O => \N__51216\,
            I => \N__51213\
        );

    \I__12248\ : Odrv4
    port map (
            O => \N__51213\,
            I => n19_adj_1497
        );

    \I__12247\ : CascadeMux
    port map (
            O => \N__51210\,
            I => \N__51207\
        );

    \I__12246\ : InMux
    port map (
            O => \N__51207\,
            I => \N__51204\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__51204\,
            I => \N__51201\
        );

    \I__12244\ : Span4Mux_v
    port map (
            O => \N__51201\,
            I => \N__51198\
        );

    \I__12243\ : Span4Mux_h
    port map (
            O => \N__51198\,
            I => \N__51195\
        );

    \I__12242\ : Span4Mux_h
    port map (
            O => \N__51195\,
            I => \N__51191\
        );

    \I__12241\ : CascadeMux
    port map (
            O => \N__51194\,
            I => \N__51188\
        );

    \I__12240\ : Span4Mux_h
    port map (
            O => \N__51191\,
            I => \N__51185\
        );

    \I__12239\ : InMux
    port map (
            O => \N__51188\,
            I => \N__51182\
        );

    \I__12238\ : Odrv4
    port map (
            O => \N__51185\,
            I => \buf_readRTD_5\
        );

    \I__12237\ : LocalMux
    port map (
            O => \N__51182\,
            I => \buf_readRTD_5\
        );

    \I__12236\ : InMux
    port map (
            O => \N__51177\,
            I => \N__51173\
        );

    \I__12235\ : CascadeMux
    port map (
            O => \N__51176\,
            I => \N__51170\
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__51173\,
            I => \N__51167\
        );

    \I__12233\ : InMux
    port map (
            O => \N__51170\,
            I => \N__51164\
        );

    \I__12232\ : Span4Mux_h
    port map (
            O => \N__51167\,
            I => \N__51161\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__51164\,
            I => data_idxvec_5
        );

    \I__12230\ : Odrv4
    port map (
            O => \N__51161\,
            I => data_idxvec_5
        );

    \I__12229\ : InMux
    port map (
            O => \N__51156\,
            I => \N__51152\
        );

    \I__12228\ : InMux
    port map (
            O => \N__51155\,
            I => \N__51148\
        );

    \I__12227\ : LocalMux
    port map (
            O => \N__51152\,
            I => \N__51145\
        );

    \I__12226\ : InMux
    port map (
            O => \N__51151\,
            I => \N__51142\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__51148\,
            I => \N__51139\
        );

    \I__12224\ : Span4Mux_h
    port map (
            O => \N__51145\,
            I => \N__51136\
        );

    \I__12223\ : LocalMux
    port map (
            O => \N__51142\,
            I => data_cntvec_5
        );

    \I__12222\ : Odrv4
    port map (
            O => \N__51139\,
            I => data_cntvec_5
        );

    \I__12221\ : Odrv4
    port map (
            O => \N__51136\,
            I => data_cntvec_5
        );

    \I__12220\ : CascadeMux
    port map (
            O => \N__51129\,
            I => \n26_adj_1498_cascade_\
        );

    \I__12219\ : CascadeMux
    port map (
            O => \N__51126\,
            I => \n21132_cascade_\
        );

    \I__12218\ : InMux
    port map (
            O => \N__51123\,
            I => \N__51120\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__51120\,
            I => n21127
        );

    \I__12216\ : CascadeMux
    port map (
            O => \N__51117\,
            I => \n22333_cascade_\
        );

    \I__12215\ : InMux
    port map (
            O => \N__51114\,
            I => \N__51111\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__51111\,
            I => \N__51103\
        );

    \I__12213\ : InMux
    port map (
            O => \N__51110\,
            I => \N__51100\
        );

    \I__12212\ : InMux
    port map (
            O => \N__51109\,
            I => \N__51097\
        );

    \I__12211\ : InMux
    port map (
            O => \N__51108\,
            I => \N__51094\
        );

    \I__12210\ : InMux
    port map (
            O => \N__51107\,
            I => \N__51091\
        );

    \I__12209\ : CascadeMux
    port map (
            O => \N__51106\,
            I => \N__51088\
        );

    \I__12208\ : Span4Mux_v
    port map (
            O => \N__51103\,
            I => \N__51083\
        );

    \I__12207\ : LocalMux
    port map (
            O => \N__51100\,
            I => \N__51083\
        );

    \I__12206\ : LocalMux
    port map (
            O => \N__51097\,
            I => \N__51078\
        );

    \I__12205\ : LocalMux
    port map (
            O => \N__51094\,
            I => \N__51078\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__51091\,
            I => \N__51075\
        );

    \I__12203\ : InMux
    port map (
            O => \N__51088\,
            I => \N__51072\
        );

    \I__12202\ : Span4Mux_v
    port map (
            O => \N__51083\,
            I => \N__51068\
        );

    \I__12201\ : Span4Mux_v
    port map (
            O => \N__51078\,
            I => \N__51065\
        );

    \I__12200\ : Span4Mux_v
    port map (
            O => \N__51075\,
            I => \N__51062\
        );

    \I__12199\ : LocalMux
    port map (
            O => \N__51072\,
            I => \N__51059\
        );

    \I__12198\ : InMux
    port map (
            O => \N__51071\,
            I => \N__51056\
        );

    \I__12197\ : Sp12to4
    port map (
            O => \N__51068\,
            I => \N__51049\
        );

    \I__12196\ : Sp12to4
    port map (
            O => \N__51065\,
            I => \N__51049\
        );

    \I__12195\ : Span4Mux_h
    port map (
            O => \N__51062\,
            I => \N__51046\
        );

    \I__12194\ : Span4Mux_v
    port map (
            O => \N__51059\,
            I => \N__51041\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__51056\,
            I => \N__51041\
        );

    \I__12192\ : InMux
    port map (
            O => \N__51055\,
            I => \N__51038\
        );

    \I__12191\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51035\
        );

    \I__12190\ : Odrv12
    port map (
            O => \N__51049\,
            I => comm_rx_buf_3
        );

    \I__12189\ : Odrv4
    port map (
            O => \N__51046\,
            I => comm_rx_buf_3
        );

    \I__12188\ : Odrv4
    port map (
            O => \N__51041\,
            I => comm_rx_buf_3
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__51038\,
            I => comm_rx_buf_3
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__51035\,
            I => comm_rx_buf_3
        );

    \I__12185\ : CascadeMux
    port map (
            O => \N__51024\,
            I => \n22336_cascade_\
        );

    \I__12184\ : CascadeMux
    port map (
            O => \N__51021\,
            I => \N__51016\
        );

    \I__12183\ : CascadeMux
    port map (
            O => \N__51020\,
            I => \N__51013\
        );

    \I__12182\ : InMux
    port map (
            O => \N__51019\,
            I => \N__51009\
        );

    \I__12181\ : InMux
    port map (
            O => \N__51016\,
            I => \N__51006\
        );

    \I__12180\ : InMux
    port map (
            O => \N__51013\,
            I => \N__51003\
        );

    \I__12179\ : InMux
    port map (
            O => \N__51012\,
            I => \N__51000\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__51009\,
            I => \N__50996\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__51006\,
            I => \N__50993\
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__51003\,
            I => \N__50990\
        );

    \I__12175\ : LocalMux
    port map (
            O => \N__51000\,
            I => \N__50987\
        );

    \I__12174\ : InMux
    port map (
            O => \N__50999\,
            I => \N__50984\
        );

    \I__12173\ : Span4Mux_v
    port map (
            O => \N__50996\,
            I => \N__50981\
        );

    \I__12172\ : Span4Mux_v
    port map (
            O => \N__50993\,
            I => \N__50978\
        );

    \I__12171\ : Span4Mux_v
    port map (
            O => \N__50990\,
            I => \N__50973\
        );

    \I__12170\ : Span4Mux_v
    port map (
            O => \N__50987\,
            I => \N__50973\
        );

    \I__12169\ : LocalMux
    port map (
            O => \N__50984\,
            I => \N__50970\
        );

    \I__12168\ : Span4Mux_v
    port map (
            O => \N__50981\,
            I => \N__50967\
        );

    \I__12167\ : Span4Mux_v
    port map (
            O => \N__50978\,
            I => \N__50962\
        );

    \I__12166\ : Span4Mux_h
    port map (
            O => \N__50973\,
            I => \N__50962\
        );

    \I__12165\ : Sp12to4
    port map (
            O => \N__50970\,
            I => \N__50959\
        );

    \I__12164\ : Span4Mux_h
    port map (
            O => \N__50967\,
            I => \N__50956\
        );

    \I__12163\ : Odrv4
    port map (
            O => \N__50962\,
            I => comm_buf_1_3
        );

    \I__12162\ : Odrv12
    port map (
            O => \N__50959\,
            I => comm_buf_1_3
        );

    \I__12161\ : Odrv4
    port map (
            O => \N__50956\,
            I => comm_buf_1_3
        );

    \I__12160\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50946\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__50946\,
            I => \N__50943\
        );

    \I__12158\ : Span4Mux_v
    port map (
            O => \N__50943\,
            I => \N__50940\
        );

    \I__12157\ : Span4Mux_h
    port map (
            O => \N__50940\,
            I => \N__50936\
        );

    \I__12156\ : CascadeMux
    port map (
            O => \N__50939\,
            I => \N__50933\
        );

    \I__12155\ : Span4Mux_h
    port map (
            O => \N__50936\,
            I => \N__50930\
        );

    \I__12154\ : InMux
    port map (
            O => \N__50933\,
            I => \N__50927\
        );

    \I__12153\ : Odrv4
    port map (
            O => \N__50930\,
            I => buf_adcdata_vdc_11
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__50927\,
            I => buf_adcdata_vdc_11
        );

    \I__12151\ : InMux
    port map (
            O => \N__50922\,
            I => \N__50917\
        );

    \I__12150\ : InMux
    port map (
            O => \N__50921\,
            I => \N__50914\
        );

    \I__12149\ : CascadeMux
    port map (
            O => \N__50920\,
            I => \N__50911\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__50917\,
            I => \N__50908\
        );

    \I__12147\ : LocalMux
    port map (
            O => \N__50914\,
            I => \N__50905\
        );

    \I__12146\ : InMux
    port map (
            O => \N__50911\,
            I => \N__50902\
        );

    \I__12145\ : Span12Mux_v
    port map (
            O => \N__50908\,
            I => \N__50899\
        );

    \I__12144\ : Span12Mux_h
    port map (
            O => \N__50905\,
            I => \N__50896\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__50902\,
            I => buf_adcdata_vac_11
        );

    \I__12142\ : Odrv12
    port map (
            O => \N__50899\,
            I => buf_adcdata_vac_11
        );

    \I__12141\ : Odrv12
    port map (
            O => \N__50896\,
            I => buf_adcdata_vac_11
        );

    \I__12140\ : InMux
    port map (
            O => \N__50889\,
            I => \N__50886\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__50886\,
            I => n19_adj_1515
        );

    \I__12138\ : InMux
    port map (
            O => \N__50883\,
            I => \N__50879\
        );

    \I__12137\ : CascadeMux
    port map (
            O => \N__50882\,
            I => \N__50876\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__50879\,
            I => \N__50873\
        );

    \I__12135\ : InMux
    port map (
            O => \N__50876\,
            I => \N__50870\
        );

    \I__12134\ : Span4Mux_v
    port map (
            O => \N__50873\,
            I => \N__50867\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__50870\,
            I => data_idxvec_3
        );

    \I__12132\ : Odrv4
    port map (
            O => \N__50867\,
            I => data_idxvec_3
        );

    \I__12131\ : InMux
    port map (
            O => \N__50862\,
            I => \N__50858\
        );

    \I__12130\ : InMux
    port map (
            O => \N__50861\,
            I => \N__50855\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__50858\,
            I => \N__50851\
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__50855\,
            I => \N__50848\
        );

    \I__12127\ : InMux
    port map (
            O => \N__50854\,
            I => \N__50845\
        );

    \I__12126\ : Span4Mux_h
    port map (
            O => \N__50851\,
            I => \N__50840\
        );

    \I__12125\ : Span4Mux_h
    port map (
            O => \N__50848\,
            I => \N__50840\
        );

    \I__12124\ : LocalMux
    port map (
            O => \N__50845\,
            I => data_cntvec_3
        );

    \I__12123\ : Odrv4
    port map (
            O => \N__50840\,
            I => data_cntvec_3
        );

    \I__12122\ : InMux
    port map (
            O => \N__50835\,
            I => \N__50832\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__50832\,
            I => \N__50829\
        );

    \I__12120\ : Span4Mux_h
    port map (
            O => \N__50829\,
            I => \N__50826\
        );

    \I__12119\ : Span4Mux_v
    port map (
            O => \N__50826\,
            I => \N__50823\
        );

    \I__12118\ : Odrv4
    port map (
            O => \N__50823\,
            I => buf_data_iac_11
        );

    \I__12117\ : CascadeMux
    port map (
            O => \N__50820\,
            I => \n26_adj_1516_cascade_\
        );

    \I__12116\ : InMux
    port map (
            O => \N__50817\,
            I => \N__50814\
        );

    \I__12115\ : LocalMux
    port map (
            O => \N__50814\,
            I => n21133
        );

    \I__12114\ : CascadeMux
    port map (
            O => \N__50811\,
            I => \n21316_cascade_\
        );

    \I__12113\ : InMux
    port map (
            O => \N__50808\,
            I => \N__50802\
        );

    \I__12112\ : InMux
    port map (
            O => \N__50807\,
            I => \N__50802\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__50802\,
            I => comm_length_2
        );

    \I__12110\ : CascadeMux
    port map (
            O => \N__50799\,
            I => \N__50787\
        );

    \I__12109\ : CascadeMux
    port map (
            O => \N__50798\,
            I => \N__50783\
        );

    \I__12108\ : InMux
    port map (
            O => \N__50797\,
            I => \N__50768\
        );

    \I__12107\ : InMux
    port map (
            O => \N__50796\,
            I => \N__50768\
        );

    \I__12106\ : InMux
    port map (
            O => \N__50795\,
            I => \N__50768\
        );

    \I__12105\ : InMux
    port map (
            O => \N__50794\,
            I => \N__50768\
        );

    \I__12104\ : InMux
    port map (
            O => \N__50793\,
            I => \N__50761\
        );

    \I__12103\ : InMux
    port map (
            O => \N__50792\,
            I => \N__50761\
        );

    \I__12102\ : InMux
    port map (
            O => \N__50791\,
            I => \N__50761\
        );

    \I__12101\ : InMux
    port map (
            O => \N__50790\,
            I => \N__50758\
        );

    \I__12100\ : InMux
    port map (
            O => \N__50787\,
            I => \N__50748\
        );

    \I__12099\ : InMux
    port map (
            O => \N__50786\,
            I => \N__50743\
        );

    \I__12098\ : InMux
    port map (
            O => \N__50783\,
            I => \N__50743\
        );

    \I__12097\ : InMux
    port map (
            O => \N__50782\,
            I => \N__50740\
        );

    \I__12096\ : CascadeMux
    port map (
            O => \N__50781\,
            I => \N__50737\
        );

    \I__12095\ : CascadeMux
    port map (
            O => \N__50780\,
            I => \N__50734\
        );

    \I__12094\ : InMux
    port map (
            O => \N__50779\,
            I => \N__50726\
        );

    \I__12093\ : InMux
    port map (
            O => \N__50778\,
            I => \N__50721\
        );

    \I__12092\ : InMux
    port map (
            O => \N__50777\,
            I => \N__50721\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__50768\,
            I => \N__50714\
        );

    \I__12090\ : LocalMux
    port map (
            O => \N__50761\,
            I => \N__50714\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__50758\,
            I => \N__50714\
        );

    \I__12088\ : InMux
    port map (
            O => \N__50757\,
            I => \N__50705\
        );

    \I__12087\ : InMux
    port map (
            O => \N__50756\,
            I => \N__50705\
        );

    \I__12086\ : InMux
    port map (
            O => \N__50755\,
            I => \N__50705\
        );

    \I__12085\ : InMux
    port map (
            O => \N__50754\,
            I => \N__50705\
        );

    \I__12084\ : InMux
    port map (
            O => \N__50753\,
            I => \N__50702\
        );

    \I__12083\ : InMux
    port map (
            O => \N__50752\,
            I => \N__50697\
        );

    \I__12082\ : InMux
    port map (
            O => \N__50751\,
            I => \N__50697\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__50748\,
            I => \N__50694\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__50743\,
            I => \N__50689\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__50740\,
            I => \N__50689\
        );

    \I__12078\ : InMux
    port map (
            O => \N__50737\,
            I => \N__50681\
        );

    \I__12077\ : InMux
    port map (
            O => \N__50734\,
            I => \N__50681\
        );

    \I__12076\ : InMux
    port map (
            O => \N__50733\,
            I => \N__50681\
        );

    \I__12075\ : InMux
    port map (
            O => \N__50732\,
            I => \N__50672\
        );

    \I__12074\ : InMux
    port map (
            O => \N__50731\,
            I => \N__50672\
        );

    \I__12073\ : InMux
    port map (
            O => \N__50730\,
            I => \N__50672\
        );

    \I__12072\ : InMux
    port map (
            O => \N__50729\,
            I => \N__50672\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__50726\,
            I => \N__50659\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__50721\,
            I => \N__50659\
        );

    \I__12069\ : Span4Mux_v
    port map (
            O => \N__50714\,
            I => \N__50659\
        );

    \I__12068\ : LocalMux
    port map (
            O => \N__50705\,
            I => \N__50659\
        );

    \I__12067\ : LocalMux
    port map (
            O => \N__50702\,
            I => \N__50654\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__50697\,
            I => \N__50647\
        );

    \I__12065\ : Span4Mux_h
    port map (
            O => \N__50694\,
            I => \N__50647\
        );

    \I__12064\ : Span4Mux_v
    port map (
            O => \N__50689\,
            I => \N__50647\
        );

    \I__12063\ : InMux
    port map (
            O => \N__50688\,
            I => \N__50644\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__50681\,
            I => \N__50639\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__50672\,
            I => \N__50639\
        );

    \I__12060\ : InMux
    port map (
            O => \N__50671\,
            I => \N__50630\
        );

    \I__12059\ : InMux
    port map (
            O => \N__50670\,
            I => \N__50630\
        );

    \I__12058\ : InMux
    port map (
            O => \N__50669\,
            I => \N__50630\
        );

    \I__12057\ : InMux
    port map (
            O => \N__50668\,
            I => \N__50630\
        );

    \I__12056\ : Span4Mux_h
    port map (
            O => \N__50659\,
            I => \N__50627\
        );

    \I__12055\ : InMux
    port map (
            O => \N__50658\,
            I => \N__50622\
        );

    \I__12054\ : InMux
    port map (
            O => \N__50657\,
            I => \N__50622\
        );

    \I__12053\ : Span4Mux_h
    port map (
            O => \N__50654\,
            I => \N__50617\
        );

    \I__12052\ : Span4Mux_h
    port map (
            O => \N__50647\,
            I => \N__50617\
        );

    \I__12051\ : LocalMux
    port map (
            O => \N__50644\,
            I => comm_index_0
        );

    \I__12050\ : Odrv4
    port map (
            O => \N__50639\,
            I => comm_index_0
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__50630\,
            I => comm_index_0
        );

    \I__12048\ : Odrv4
    port map (
            O => \N__50627\,
            I => comm_index_0
        );

    \I__12047\ : LocalMux
    port map (
            O => \N__50622\,
            I => comm_index_0
        );

    \I__12046\ : Odrv4
    port map (
            O => \N__50617\,
            I => comm_index_0
        );

    \I__12045\ : InMux
    port map (
            O => \N__50604\,
            I => \N__50588\
        );

    \I__12044\ : InMux
    port map (
            O => \N__50603\,
            I => \N__50588\
        );

    \I__12043\ : InMux
    port map (
            O => \N__50602\,
            I => \N__50585\
        );

    \I__12042\ : InMux
    port map (
            O => \N__50601\,
            I => \N__50581\
        );

    \I__12041\ : InMux
    port map (
            O => \N__50600\,
            I => \N__50573\
        );

    \I__12040\ : InMux
    port map (
            O => \N__50599\,
            I => \N__50573\
        );

    \I__12039\ : InMux
    port map (
            O => \N__50598\,
            I => \N__50566\
        );

    \I__12038\ : InMux
    port map (
            O => \N__50597\,
            I => \N__50566\
        );

    \I__12037\ : InMux
    port map (
            O => \N__50596\,
            I => \N__50557\
        );

    \I__12036\ : InMux
    port map (
            O => \N__50595\,
            I => \N__50557\
        );

    \I__12035\ : InMux
    port map (
            O => \N__50594\,
            I => \N__50557\
        );

    \I__12034\ : InMux
    port map (
            O => \N__50593\,
            I => \N__50557\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__50588\,
            I => \N__50552\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__50585\,
            I => \N__50552\
        );

    \I__12031\ : InMux
    port map (
            O => \N__50584\,
            I => \N__50549\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__50581\,
            I => \N__50546\
        );

    \I__12029\ : InMux
    port map (
            O => \N__50580\,
            I => \N__50543\
        );

    \I__12028\ : InMux
    port map (
            O => \N__50579\,
            I => \N__50540\
        );

    \I__12027\ : InMux
    port map (
            O => \N__50578\,
            I => \N__50535\
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__50573\,
            I => \N__50532\
        );

    \I__12025\ : InMux
    port map (
            O => \N__50572\,
            I => \N__50527\
        );

    \I__12024\ : InMux
    port map (
            O => \N__50571\,
            I => \N__50527\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__50566\,
            I => \N__50522\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__50557\,
            I => \N__50522\
        );

    \I__12021\ : Span4Mux_v
    port map (
            O => \N__50552\,
            I => \N__50515\
        );

    \I__12020\ : LocalMux
    port map (
            O => \N__50549\,
            I => \N__50515\
        );

    \I__12019\ : Span4Mux_v
    port map (
            O => \N__50546\,
            I => \N__50515\
        );

    \I__12018\ : LocalMux
    port map (
            O => \N__50543\,
            I => \N__50510\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__50540\,
            I => \N__50510\
        );

    \I__12016\ : InMux
    port map (
            O => \N__50539\,
            I => \N__50505\
        );

    \I__12015\ : InMux
    port map (
            O => \N__50538\,
            I => \N__50505\
        );

    \I__12014\ : LocalMux
    port map (
            O => \N__50535\,
            I => \N__50498\
        );

    \I__12013\ : Span4Mux_h
    port map (
            O => \N__50532\,
            I => \N__50498\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__50527\,
            I => \N__50498\
        );

    \I__12011\ : Span4Mux_h
    port map (
            O => \N__50522\,
            I => \N__50495\
        );

    \I__12010\ : Span4Mux_h
    port map (
            O => \N__50515\,
            I => \N__50490\
        );

    \I__12009\ : Span4Mux_v
    port map (
            O => \N__50510\,
            I => \N__50490\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__50505\,
            I => comm_index_2
        );

    \I__12007\ : Odrv4
    port map (
            O => \N__50498\,
            I => comm_index_2
        );

    \I__12006\ : Odrv4
    port map (
            O => \N__50495\,
            I => comm_index_2
        );

    \I__12005\ : Odrv4
    port map (
            O => \N__50490\,
            I => comm_index_2
        );

    \I__12004\ : CascadeMux
    port map (
            O => \N__50481\,
            I => \n22267_cascade_\
        );

    \I__12003\ : InMux
    port map (
            O => \N__50478\,
            I => \N__50474\
        );

    \I__12002\ : CascadeMux
    port map (
            O => \N__50477\,
            I => \N__50471\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__50474\,
            I => \N__50468\
        );

    \I__12000\ : InMux
    port map (
            O => \N__50471\,
            I => \N__50465\
        );

    \I__11999\ : Span4Mux_h
    port map (
            O => \N__50468\,
            I => \N__50462\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__50465\,
            I => data_idxvec_7
        );

    \I__11997\ : Odrv4
    port map (
            O => \N__50462\,
            I => data_idxvec_7
        );

    \I__11996\ : InMux
    port map (
            O => \N__50457\,
            I => \N__50454\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__50454\,
            I => \N__50449\
        );

    \I__11994\ : InMux
    port map (
            O => \N__50453\,
            I => \N__50446\
        );

    \I__11993\ : InMux
    port map (
            O => \N__50452\,
            I => \N__50443\
        );

    \I__11992\ : Span12Mux_h
    port map (
            O => \N__50449\,
            I => \N__50440\
        );

    \I__11991\ : LocalMux
    port map (
            O => \N__50446\,
            I => data_cntvec_7
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__50443\,
            I => data_cntvec_7
        );

    \I__11989\ : Odrv12
    port map (
            O => \N__50440\,
            I => data_cntvec_7
        );

    \I__11988\ : InMux
    port map (
            O => \N__50433\,
            I => \N__50430\
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__50430\,
            I => \N__50427\
        );

    \I__11986\ : Span12Mux_h
    port map (
            O => \N__50427\,
            I => \N__50424\
        );

    \I__11985\ : Odrv12
    port map (
            O => \N__50424\,
            I => buf_data_iac_15
        );

    \I__11984\ : CascadeMux
    port map (
            O => \N__50421\,
            I => \n26_adj_1502_cascade_\
        );

    \I__11983\ : InMux
    port map (
            O => \N__50418\,
            I => \N__50415\
        );

    \I__11982\ : LocalMux
    port map (
            O => \N__50415\,
            I => n21055
        );

    \I__11981\ : CascadeMux
    port map (
            O => \N__50412\,
            I => \N__50405\
        );

    \I__11980\ : InMux
    port map (
            O => \N__50411\,
            I => \N__50402\
        );

    \I__11979\ : InMux
    port map (
            O => \N__50410\,
            I => \N__50399\
        );

    \I__11978\ : InMux
    port map (
            O => \N__50409\,
            I => \N__50396\
        );

    \I__11977\ : InMux
    port map (
            O => \N__50408\,
            I => \N__50393\
        );

    \I__11976\ : InMux
    port map (
            O => \N__50405\,
            I => \N__50390\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__50402\,
            I => \N__50384\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__50399\,
            I => \N__50384\
        );

    \I__11973\ : LocalMux
    port map (
            O => \N__50396\,
            I => \N__50381\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__50393\,
            I => \N__50377\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__50390\,
            I => \N__50374\
        );

    \I__11970\ : InMux
    port map (
            O => \N__50389\,
            I => \N__50371\
        );

    \I__11969\ : Span4Mux_v
    port map (
            O => \N__50384\,
            I => \N__50366\
        );

    \I__11968\ : Span4Mux_h
    port map (
            O => \N__50381\,
            I => \N__50366\
        );

    \I__11967\ : InMux
    port map (
            O => \N__50380\,
            I => \N__50363\
        );

    \I__11966\ : Span4Mux_v
    port map (
            O => \N__50377\,
            I => \N__50358\
        );

    \I__11965\ : Span4Mux_v
    port map (
            O => \N__50374\,
            I => \N__50358\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__50371\,
            I => \N__50355\
        );

    \I__11963\ : Span4Mux_h
    port map (
            O => \N__50366\,
            I => \N__50350\
        );

    \I__11962\ : LocalMux
    port map (
            O => \N__50363\,
            I => \N__50350\
        );

    \I__11961\ : Sp12to4
    port map (
            O => \N__50358\,
            I => \N__50346\
        );

    \I__11960\ : Span4Mux_v
    port map (
            O => \N__50355\,
            I => \N__50343\
        );

    \I__11959\ : Span4Mux_v
    port map (
            O => \N__50350\,
            I => \N__50340\
        );

    \I__11958\ : InMux
    port map (
            O => \N__50349\,
            I => \N__50337\
        );

    \I__11957\ : Odrv12
    port map (
            O => \N__50346\,
            I => comm_rx_buf_7
        );

    \I__11956\ : Odrv4
    port map (
            O => \N__50343\,
            I => comm_rx_buf_7
        );

    \I__11955\ : Odrv4
    port map (
            O => \N__50340\,
            I => comm_rx_buf_7
        );

    \I__11954\ : LocalMux
    port map (
            O => \N__50337\,
            I => comm_rx_buf_7
        );

    \I__11953\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50325\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__50325\,
            I => n22270
        );

    \I__11951\ : CascadeMux
    port map (
            O => \N__50322\,
            I => \N__50315\
        );

    \I__11950\ : CascadeMux
    port map (
            O => \N__50321\,
            I => \N__50312\
        );

    \I__11949\ : CascadeMux
    port map (
            O => \N__50320\,
            I => \N__50309\
        );

    \I__11948\ : InMux
    port map (
            O => \N__50319\,
            I => \N__50306\
        );

    \I__11947\ : InMux
    port map (
            O => \N__50318\,
            I => \N__50303\
        );

    \I__11946\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50299\
        );

    \I__11945\ : InMux
    port map (
            O => \N__50312\,
            I => \N__50296\
        );

    \I__11944\ : InMux
    port map (
            O => \N__50309\,
            I => \N__50293\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__50306\,
            I => \N__50290\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__50303\,
            I => \N__50287\
        );

    \I__11941\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50284\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__50299\,
            I => \N__50281\
        );

    \I__11939\ : LocalMux
    port map (
            O => \N__50296\,
            I => \N__50278\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__50293\,
            I => \N__50275\
        );

    \I__11937\ : Span4Mux_v
    port map (
            O => \N__50290\,
            I => \N__50272\
        );

    \I__11936\ : Span4Mux_h
    port map (
            O => \N__50287\,
            I => \N__50267\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__50284\,
            I => \N__50267\
        );

    \I__11934\ : Span4Mux_h
    port map (
            O => \N__50281\,
            I => \N__50264\
        );

    \I__11933\ : Span4Mux_v
    port map (
            O => \N__50278\,
            I => \N__50257\
        );

    \I__11932\ : Span4Mux_v
    port map (
            O => \N__50275\,
            I => \N__50257\
        );

    \I__11931\ : Span4Mux_h
    port map (
            O => \N__50272\,
            I => \N__50257\
        );

    \I__11930\ : Span4Mux_h
    port map (
            O => \N__50267\,
            I => \N__50254\
        );

    \I__11929\ : Span4Mux_v
    port map (
            O => \N__50264\,
            I => \N__50251\
        );

    \I__11928\ : Sp12to4
    port map (
            O => \N__50257\,
            I => \N__50248\
        );

    \I__11927\ : Span4Mux_v
    port map (
            O => \N__50254\,
            I => \N__50245\
        );

    \I__11926\ : Odrv4
    port map (
            O => \N__50251\,
            I => comm_buf_1_7
        );

    \I__11925\ : Odrv12
    port map (
            O => \N__50248\,
            I => comm_buf_1_7
        );

    \I__11924\ : Odrv4
    port map (
            O => \N__50245\,
            I => comm_buf_1_7
        );

    \I__11923\ : InMux
    port map (
            O => \N__50238\,
            I => \N__50235\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__50235\,
            I => \N__50232\
        );

    \I__11921\ : Span12Mux_h
    port map (
            O => \N__50232\,
            I => \N__50228\
        );

    \I__11920\ : InMux
    port map (
            O => \N__50231\,
            I => \N__50225\
        );

    \I__11919\ : Odrv12
    port map (
            O => \N__50228\,
            I => buf_adcdata_vdc_15
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__50225\,
            I => buf_adcdata_vdc_15
        );

    \I__11917\ : InMux
    port map (
            O => \N__50220\,
            I => \N__50217\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__50217\,
            I => \N__50213\
        );

    \I__11915\ : InMux
    port map (
            O => \N__50216\,
            I => \N__50210\
        );

    \I__11914\ : Span4Mux_v
    port map (
            O => \N__50213\,
            I => \N__50205\
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__50210\,
            I => \N__50205\
        );

    \I__11912\ : Span4Mux_h
    port map (
            O => \N__50205\,
            I => \N__50202\
        );

    \I__11911\ : Span4Mux_h
    port map (
            O => \N__50202\,
            I => \N__50198\
        );

    \I__11910\ : InMux
    port map (
            O => \N__50201\,
            I => \N__50195\
        );

    \I__11909\ : Span4Mux_h
    port map (
            O => \N__50198\,
            I => \N__50192\
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__50195\,
            I => buf_adcdata_vac_15
        );

    \I__11907\ : Odrv4
    port map (
            O => \N__50192\,
            I => buf_adcdata_vac_15
        );

    \I__11906\ : CascadeMux
    port map (
            O => \N__50187\,
            I => \n19_adj_1503_cascade_\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50184\,
            I => \N__50181\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__50181\,
            I => \N__50178\
        );

    \I__11903\ : Span12Mux_s11_h
    port map (
            O => \N__50178\,
            I => \N__50174\
        );

    \I__11902\ : CascadeMux
    port map (
            O => \N__50177\,
            I => \N__50171\
        );

    \I__11901\ : Span12Mux_h
    port map (
            O => \N__50174\,
            I => \N__50168\
        );

    \I__11900\ : InMux
    port map (
            O => \N__50171\,
            I => \N__50165\
        );

    \I__11899\ : Odrv12
    port map (
            O => \N__50168\,
            I => \buf_readRTD_7\
        );

    \I__11898\ : LocalMux
    port map (
            O => \N__50165\,
            I => \buf_readRTD_7\
        );

    \I__11897\ : InMux
    port map (
            O => \N__50160\,
            I => \N__50157\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__50157\,
            I => n21049
        );

    \I__11895\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50151\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__50151\,
            I => \N__50148\
        );

    \I__11893\ : Span4Mux_v
    port map (
            O => \N__50148\,
            I => \N__50145\
        );

    \I__11892\ : Span4Mux_h
    port map (
            O => \N__50145\,
            I => \N__50142\
        );

    \I__11891\ : Span4Mux_h
    port map (
            O => \N__50142\,
            I => \N__50138\
        );

    \I__11890\ : CascadeMux
    port map (
            O => \N__50141\,
            I => \N__50135\
        );

    \I__11889\ : Span4Mux_h
    port map (
            O => \N__50138\,
            I => \N__50132\
        );

    \I__11888\ : InMux
    port map (
            O => \N__50135\,
            I => \N__50129\
        );

    \I__11887\ : Odrv4
    port map (
            O => \N__50132\,
            I => \buf_readRTD_3\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__50129\,
            I => \buf_readRTD_3\
        );

    \I__11885\ : InMux
    port map (
            O => \N__50124\,
            I => \N__50121\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__50121\,
            I => \N__50118\
        );

    \I__11883\ : Span4Mux_h
    port map (
            O => \N__50118\,
            I => \N__50114\
        );

    \I__11882\ : CascadeMux
    port map (
            O => \N__50117\,
            I => \N__50110\
        );

    \I__11881\ : Span4Mux_v
    port map (
            O => \N__50114\,
            I => \N__50107\
        );

    \I__11880\ : CascadeMux
    port map (
            O => \N__50113\,
            I => \N__50104\
        );

    \I__11879\ : InMux
    port map (
            O => \N__50110\,
            I => \N__50101\
        );

    \I__11878\ : Span4Mux_h
    port map (
            O => \N__50107\,
            I => \N__50098\
        );

    \I__11877\ : InMux
    port map (
            O => \N__50104\,
            I => \N__50095\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__50101\,
            I => req_data_cnt_3
        );

    \I__11875\ : Odrv4
    port map (
            O => \N__50098\,
            I => req_data_cnt_3
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__50095\,
            I => req_data_cnt_3
        );

    \I__11873\ : InMux
    port map (
            O => \N__50088\,
            I => \N__50084\
        );

    \I__11872\ : CascadeMux
    port map (
            O => \N__50087\,
            I => \N__50081\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__50084\,
            I => \N__50077\
        );

    \I__11870\ : InMux
    port map (
            O => \N__50081\,
            I => \N__50074\
        );

    \I__11869\ : InMux
    port map (
            O => \N__50080\,
            I => \N__50071\
        );

    \I__11868\ : Span12Mux_h
    port map (
            O => \N__50077\,
            I => \N__50068\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__50074\,
            I => \N__50065\
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__50071\,
            I => \acadc_skipCount_3\
        );

    \I__11865\ : Odrv12
    port map (
            O => \N__50068\,
            I => \acadc_skipCount_3\
        );

    \I__11864\ : Odrv4
    port map (
            O => \N__50065\,
            I => \acadc_skipCount_3\
        );

    \I__11863\ : InMux
    port map (
            O => \N__50058\,
            I => \N__50055\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__50055\,
            I => n12_adj_1548
        );

    \I__11861\ : InMux
    port map (
            O => \N__50052\,
            I => \N__50048\
        );

    \I__11860\ : CascadeMux
    port map (
            O => \N__50051\,
            I => \N__50042\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__50048\,
            I => \N__50039\
        );

    \I__11858\ : CascadeMux
    port map (
            O => \N__50047\,
            I => \N__50032\
        );

    \I__11857\ : CascadeMux
    port map (
            O => \N__50046\,
            I => \N__50027\
        );

    \I__11856\ : InMux
    port map (
            O => \N__50045\,
            I => \N__50023\
        );

    \I__11855\ : InMux
    port map (
            O => \N__50042\,
            I => \N__50020\
        );

    \I__11854\ : Span4Mux_h
    port map (
            O => \N__50039\,
            I => \N__50017\
        );

    \I__11853\ : InMux
    port map (
            O => \N__50038\,
            I => \N__50014\
        );

    \I__11852\ : CascadeMux
    port map (
            O => \N__50037\,
            I => \N__50009\
        );

    \I__11851\ : InMux
    port map (
            O => \N__50036\,
            I => \N__50001\
        );

    \I__11850\ : InMux
    port map (
            O => \N__50035\,
            I => \N__50001\
        );

    \I__11849\ : InMux
    port map (
            O => \N__50032\,
            I => \N__50001\
        );

    \I__11848\ : CascadeMux
    port map (
            O => \N__50031\,
            I => \N__49998\
        );

    \I__11847\ : CascadeMux
    port map (
            O => \N__50030\,
            I => \N__49995\
        );

    \I__11846\ : InMux
    port map (
            O => \N__50027\,
            I => \N__49990\
        );

    \I__11845\ : InMux
    port map (
            O => \N__50026\,
            I => \N__49987\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__50023\,
            I => \N__49984\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__50020\,
            I => \N__49981\
        );

    \I__11842\ : Span4Mux_v
    port map (
            O => \N__50017\,
            I => \N__49976\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__50014\,
            I => \N__49976\
        );

    \I__11840\ : InMux
    port map (
            O => \N__50013\,
            I => \N__49973\
        );

    \I__11839\ : InMux
    port map (
            O => \N__50012\,
            I => \N__49966\
        );

    \I__11838\ : InMux
    port map (
            O => \N__50009\,
            I => \N__49966\
        );

    \I__11837\ : InMux
    port map (
            O => \N__50008\,
            I => \N__49966\
        );

    \I__11836\ : LocalMux
    port map (
            O => \N__50001\,
            I => \N__49961\
        );

    \I__11835\ : InMux
    port map (
            O => \N__49998\,
            I => \N__49952\
        );

    \I__11834\ : InMux
    port map (
            O => \N__49995\,
            I => \N__49952\
        );

    \I__11833\ : InMux
    port map (
            O => \N__49994\,
            I => \N__49952\
        );

    \I__11832\ : InMux
    port map (
            O => \N__49993\,
            I => \N__49952\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__49990\,
            I => \N__49949\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__49987\,
            I => \N__49946\
        );

    \I__11829\ : Span4Mux_h
    port map (
            O => \N__49984\,
            I => \N__49941\
        );

    \I__11828\ : Span4Mux_h
    port map (
            O => \N__49981\,
            I => \N__49941\
        );

    \I__11827\ : Span4Mux_v
    port map (
            O => \N__49976\,
            I => \N__49936\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__49973\,
            I => \N__49936\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__49966\,
            I => \N__49933\
        );

    \I__11824\ : InMux
    port map (
            O => \N__49965\,
            I => \N__49928\
        );

    \I__11823\ : InMux
    port map (
            O => \N__49964\,
            I => \N__49928\
        );

    \I__11822\ : Span4Mux_v
    port map (
            O => \N__49961\,
            I => \N__49921\
        );

    \I__11821\ : LocalMux
    port map (
            O => \N__49952\,
            I => \N__49921\
        );

    \I__11820\ : Span4Mux_v
    port map (
            O => \N__49949\,
            I => \N__49921\
        );

    \I__11819\ : Span4Mux_v
    port map (
            O => \N__49946\,
            I => \N__49918\
        );

    \I__11818\ : Span4Mux_v
    port map (
            O => \N__49941\,
            I => \N__49913\
        );

    \I__11817\ : Span4Mux_h
    port map (
            O => \N__49936\,
            I => \N__49913\
        );

    \I__11816\ : Span12Mux_v
    port map (
            O => \N__49933\,
            I => \N__49908\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__49928\,
            I => \N__49908\
        );

    \I__11814\ : Sp12to4
    port map (
            O => \N__49921\,
            I => \N__49905\
        );

    \I__11813\ : Sp12to4
    port map (
            O => \N__49918\,
            I => \N__49900\
        );

    \I__11812\ : Sp12to4
    port map (
            O => \N__49913\,
            I => \N__49900\
        );

    \I__11811\ : Span12Mux_v
    port map (
            O => \N__49908\,
            I => \N__49897\
        );

    \I__11810\ : Span12Mux_h
    port map (
            O => \N__49905\,
            I => \N__49894\
        );

    \I__11809\ : Span12Mux_v
    port map (
            O => \N__49900\,
            I => \N__49891\
        );

    \I__11808\ : Span12Mux_h
    port map (
            O => \N__49897\,
            I => \N__49886\
        );

    \I__11807\ : Span12Mux_v
    port map (
            O => \N__49894\,
            I => \N__49886\
        );

    \I__11806\ : Odrv12
    port map (
            O => \N__49891\,
            I => \ICE_SPI_CE0\
        );

    \I__11805\ : Odrv12
    port map (
            O => \N__49886\,
            I => \ICE_SPI_CE0\
        );

    \I__11804\ : InMux
    port map (
            O => \N__49881\,
            I => \N__49878\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__49878\,
            I => \N__49868\
        );

    \I__11802\ : CascadeMux
    port map (
            O => \N__49877\,
            I => \N__49864\
        );

    \I__11801\ : InMux
    port map (
            O => \N__49876\,
            I => \N__49859\
        );

    \I__11800\ : InMux
    port map (
            O => \N__49875\,
            I => \N__49859\
        );

    \I__11799\ : InMux
    port map (
            O => \N__49874\,
            I => \N__49850\
        );

    \I__11798\ : InMux
    port map (
            O => \N__49873\,
            I => \N__49850\
        );

    \I__11797\ : InMux
    port map (
            O => \N__49872\,
            I => \N__49850\
        );

    \I__11796\ : InMux
    port map (
            O => \N__49871\,
            I => \N__49850\
        );

    \I__11795\ : Span4Mux_v
    port map (
            O => \N__49868\,
            I => \N__49843\
        );

    \I__11794\ : InMux
    port map (
            O => \N__49867\,
            I => \N__49840\
        );

    \I__11793\ : InMux
    port map (
            O => \N__49864\,
            I => \N__49837\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__49859\,
            I => \N__49832\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__49850\,
            I => \N__49832\
        );

    \I__11790\ : InMux
    port map (
            O => \N__49849\,
            I => \N__49829\
        );

    \I__11789\ : InMux
    port map (
            O => \N__49848\,
            I => \N__49826\
        );

    \I__11788\ : InMux
    port map (
            O => \N__49847\,
            I => \N__49823\
        );

    \I__11787\ : InMux
    port map (
            O => \N__49846\,
            I => \N__49820\
        );

    \I__11786\ : Sp12to4
    port map (
            O => \N__49843\,
            I => \N__49813\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__49840\,
            I => \N__49813\
        );

    \I__11784\ : LocalMux
    port map (
            O => \N__49837\,
            I => \N__49813\
        );

    \I__11783\ : Odrv4
    port map (
            O => \N__49832\,
            I => comm_data_vld
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49829\,
            I => comm_data_vld
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__49826\,
            I => comm_data_vld
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__49823\,
            I => comm_data_vld
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__49820\,
            I => comm_data_vld
        );

    \I__11778\ : Odrv12
    port map (
            O => \N__49813\,
            I => comm_data_vld
        );

    \I__11777\ : InMux
    port map (
            O => \N__49800\,
            I => \N__49797\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__49797\,
            I => n18984
        );

    \I__11775\ : InMux
    port map (
            O => \N__49794\,
            I => \N__49790\
        );

    \I__11774\ : InMux
    port map (
            O => \N__49793\,
            I => \N__49787\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__49790\,
            I => \N__49781\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__49787\,
            I => \N__49781\
        );

    \I__11771\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49778\
        );

    \I__11770\ : Span4Mux_v
    port map (
            O => \N__49781\,
            I => \N__49773\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__49778\,
            I => \N__49770\
        );

    \I__11768\ : InMux
    port map (
            O => \N__49777\,
            I => \N__49767\
        );

    \I__11767\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49764\
        );

    \I__11766\ : Span4Mux_h
    port map (
            O => \N__49773\,
            I => \N__49761\
        );

    \I__11765\ : Sp12to4
    port map (
            O => \N__49770\,
            I => \N__49756\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__49767\,
            I => \N__49756\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__49764\,
            I => comm_cmd_4
        );

    \I__11762\ : Odrv4
    port map (
            O => \N__49761\,
            I => comm_cmd_4
        );

    \I__11761\ : Odrv12
    port map (
            O => \N__49756\,
            I => comm_cmd_4
        );

    \I__11760\ : InMux
    port map (
            O => \N__49749\,
            I => \N__49745\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49748\,
            I => \N__49742\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__49745\,
            I => \N__49737\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__49742\,
            I => \N__49737\
        );

    \I__11756\ : Span4Mux_h
    port map (
            O => \N__49737\,
            I => \N__49734\
        );

    \I__11755\ : Span4Mux_h
    port map (
            O => \N__49734\,
            I => \N__49728\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49733\,
            I => \N__49723\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49732\,
            I => \N__49723\
        );

    \I__11752\ : InMux
    port map (
            O => \N__49731\,
            I => \N__49720\
        );

    \I__11751\ : Odrv4
    port map (
            O => \N__49728\,
            I => comm_cmd_6
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__49723\,
            I => comm_cmd_6
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__49720\,
            I => comm_cmd_6
        );

    \I__11748\ : InMux
    port map (
            O => \N__49713\,
            I => \N__49709\
        );

    \I__11747\ : InMux
    port map (
            O => \N__49712\,
            I => \N__49706\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__49709\,
            I => \N__49701\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__49706\,
            I => \N__49701\
        );

    \I__11744\ : Span4Mux_h
    port map (
            O => \N__49701\,
            I => \N__49697\
        );

    \I__11743\ : InMux
    port map (
            O => \N__49700\,
            I => \N__49692\
        );

    \I__11742\ : Span4Mux_v
    port map (
            O => \N__49697\,
            I => \N__49689\
        );

    \I__11741\ : InMux
    port map (
            O => \N__49696\,
            I => \N__49686\
        );

    \I__11740\ : InMux
    port map (
            O => \N__49695\,
            I => \N__49683\
        );

    \I__11739\ : LocalMux
    port map (
            O => \N__49692\,
            I => comm_cmd_5
        );

    \I__11738\ : Odrv4
    port map (
            O => \N__49689\,
            I => comm_cmd_5
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__49686\,
            I => comm_cmd_5
        );

    \I__11736\ : LocalMux
    port map (
            O => \N__49683\,
            I => comm_cmd_5
        );

    \I__11735\ : CascadeMux
    port map (
            O => \N__49674\,
            I => \N__49671\
        );

    \I__11734\ : InMux
    port map (
            O => \N__49671\,
            I => \N__49668\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__49668\,
            I => n21546
        );

    \I__11732\ : InMux
    port map (
            O => \N__49665\,
            I => \N__49662\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__49662\,
            I => \N__49659\
        );

    \I__11730\ : Odrv4
    port map (
            O => \N__49659\,
            I => n12092
        );

    \I__11729\ : InMux
    port map (
            O => \N__49656\,
            I => \N__49650\
        );

    \I__11728\ : InMux
    port map (
            O => \N__49655\,
            I => \N__49643\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49654\,
            I => \N__49643\
        );

    \I__11726\ : InMux
    port map (
            O => \N__49653\,
            I => \N__49643\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__49650\,
            I => \N__49640\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__49643\,
            I => \N__49637\
        );

    \I__11723\ : Span4Mux_h
    port map (
            O => \N__49640\,
            I => \N__49634\
        );

    \I__11722\ : Span4Mux_v
    port map (
            O => \N__49637\,
            I => \N__49629\
        );

    \I__11721\ : Span4Mux_h
    port map (
            O => \N__49634\,
            I => \N__49629\
        );

    \I__11720\ : Span4Mux_h
    port map (
            O => \N__49629\,
            I => \N__49626\
        );

    \I__11719\ : Odrv4
    port map (
            O => \N__49626\,
            I => n12219
        );

    \I__11718\ : InMux
    port map (
            O => \N__49623\,
            I => \N__49620\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__49620\,
            I => \N__49616\
        );

    \I__11716\ : InMux
    port map (
            O => \N__49619\,
            I => \N__49613\
        );

    \I__11715\ : Span4Mux_h
    port map (
            O => \N__49616\,
            I => \N__49610\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__49613\,
            I => n9255
        );

    \I__11713\ : Odrv4
    port map (
            O => \N__49610\,
            I => n9255
        );

    \I__11712\ : CascadeMux
    port map (
            O => \N__49605\,
            I => \n11853_cascade_\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49602\,
            I => \N__49598\
        );

    \I__11710\ : InMux
    port map (
            O => \N__49601\,
            I => \N__49595\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__49598\,
            I => \N__49592\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__49595\,
            I => \N__49582\
        );

    \I__11707\ : Span4Mux_v
    port map (
            O => \N__49592\,
            I => \N__49579\
        );

    \I__11706\ : CascadeMux
    port map (
            O => \N__49591\,
            I => \N__49576\
        );

    \I__11705\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49567\
        );

    \I__11704\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49567\
        );

    \I__11703\ : InMux
    port map (
            O => \N__49588\,
            I => \N__49567\
        );

    \I__11702\ : InMux
    port map (
            O => \N__49587\,
            I => \N__49563\
        );

    \I__11701\ : InMux
    port map (
            O => \N__49586\,
            I => \N__49559\
        );

    \I__11700\ : InMux
    port map (
            O => \N__49585\,
            I => \N__49556\
        );

    \I__11699\ : Span4Mux_v
    port map (
            O => \N__49582\,
            I => \N__49553\
        );

    \I__11698\ : Span4Mux_h
    port map (
            O => \N__49579\,
            I => \N__49550\
        );

    \I__11697\ : InMux
    port map (
            O => \N__49576\,
            I => \N__49543\
        );

    \I__11696\ : InMux
    port map (
            O => \N__49575\,
            I => \N__49543\
        );

    \I__11695\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49543\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__49567\,
            I => \N__49540\
        );

    \I__11693\ : InMux
    port map (
            O => \N__49566\,
            I => \N__49537\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__49563\,
            I => \N__49534\
        );

    \I__11691\ : InMux
    port map (
            O => \N__49562\,
            I => \N__49531\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__49559\,
            I => \N__49526\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__49556\,
            I => \N__49526\
        );

    \I__11688\ : Span4Mux_h
    port map (
            O => \N__49553\,
            I => \N__49519\
        );

    \I__11687\ : Span4Mux_v
    port map (
            O => \N__49550\,
            I => \N__49519\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__49543\,
            I => \N__49519\
        );

    \I__11685\ : Span4Mux_h
    port map (
            O => \N__49540\,
            I => \N__49512\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__49537\,
            I => \N__49512\
        );

    \I__11683\ : Span4Mux_h
    port map (
            O => \N__49534\,
            I => \N__49512\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__49531\,
            I => n12226
        );

    \I__11681\ : Odrv12
    port map (
            O => \N__49526\,
            I => n12226
        );

    \I__11680\ : Odrv4
    port map (
            O => \N__49519\,
            I => n12226
        );

    \I__11679\ : Odrv4
    port map (
            O => \N__49512\,
            I => n12226
        );

    \I__11678\ : InMux
    port map (
            O => \N__49503\,
            I => \N__49500\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__49500\,
            I => \N__49478\
        );

    \I__11676\ : InMux
    port map (
            O => \N__49499\,
            I => \N__49471\
        );

    \I__11675\ : InMux
    port map (
            O => \N__49498\,
            I => \N__49471\
        );

    \I__11674\ : InMux
    port map (
            O => \N__49497\,
            I => \N__49471\
        );

    \I__11673\ : CascadeMux
    port map (
            O => \N__49496\,
            I => \N__49468\
        );

    \I__11672\ : CascadeMux
    port map (
            O => \N__49495\,
            I => \N__49465\
        );

    \I__11671\ : CascadeMux
    port map (
            O => \N__49494\,
            I => \N__49460\
        );

    \I__11670\ : InMux
    port map (
            O => \N__49493\,
            I => \N__49457\
        );

    \I__11669\ : InMux
    port map (
            O => \N__49492\,
            I => \N__49454\
        );

    \I__11668\ : InMux
    port map (
            O => \N__49491\,
            I => \N__49449\
        );

    \I__11667\ : InMux
    port map (
            O => \N__49490\,
            I => \N__49449\
        );

    \I__11666\ : InMux
    port map (
            O => \N__49489\,
            I => \N__49446\
        );

    \I__11665\ : InMux
    port map (
            O => \N__49488\,
            I => \N__49439\
        );

    \I__11664\ : InMux
    port map (
            O => \N__49487\,
            I => \N__49439\
        );

    \I__11663\ : InMux
    port map (
            O => \N__49486\,
            I => \N__49439\
        );

    \I__11662\ : InMux
    port map (
            O => \N__49485\,
            I => \N__49430\
        );

    \I__11661\ : InMux
    port map (
            O => \N__49484\,
            I => \N__49430\
        );

    \I__11660\ : InMux
    port map (
            O => \N__49483\,
            I => \N__49430\
        );

    \I__11659\ : InMux
    port map (
            O => \N__49482\,
            I => \N__49430\
        );

    \I__11658\ : InMux
    port map (
            O => \N__49481\,
            I => \N__49427\
        );

    \I__11657\ : Span4Mux_v
    port map (
            O => \N__49478\,
            I => \N__49420\
        );

    \I__11656\ : LocalMux
    port map (
            O => \N__49471\,
            I => \N__49420\
        );

    \I__11655\ : InMux
    port map (
            O => \N__49468\,
            I => \N__49417\
        );

    \I__11654\ : InMux
    port map (
            O => \N__49465\,
            I => \N__49414\
        );

    \I__11653\ : InMux
    port map (
            O => \N__49464\,
            I => \N__49394\
        );

    \I__11652\ : InMux
    port map (
            O => \N__49463\,
            I => \N__49394\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49460\,
            I => \N__49394\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__49457\,
            I => \N__49391\
        );

    \I__11649\ : LocalMux
    port map (
            O => \N__49454\,
            I => \N__49388\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__49449\,
            I => \N__49385\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__49446\,
            I => \N__49380\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__49439\,
            I => \N__49380\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__49430\,
            I => \N__49375\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__49427\,
            I => \N__49375\
        );

    \I__11643\ : InMux
    port map (
            O => \N__49426\,
            I => \N__49372\
        );

    \I__11642\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49369\
        );

    \I__11641\ : Span4Mux_h
    port map (
            O => \N__49420\,
            I => \N__49362\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__49417\,
            I => \N__49362\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__49414\,
            I => \N__49362\
        );

    \I__11638\ : InMux
    port map (
            O => \N__49413\,
            I => \N__49353\
        );

    \I__11637\ : InMux
    port map (
            O => \N__49412\,
            I => \N__49353\
        );

    \I__11636\ : InMux
    port map (
            O => \N__49411\,
            I => \N__49353\
        );

    \I__11635\ : InMux
    port map (
            O => \N__49410\,
            I => \N__49353\
        );

    \I__11634\ : InMux
    port map (
            O => \N__49409\,
            I => \N__49348\
        );

    \I__11633\ : InMux
    port map (
            O => \N__49408\,
            I => \N__49348\
        );

    \I__11632\ : InMux
    port map (
            O => \N__49407\,
            I => \N__49339\
        );

    \I__11631\ : InMux
    port map (
            O => \N__49406\,
            I => \N__49339\
        );

    \I__11630\ : InMux
    port map (
            O => \N__49405\,
            I => \N__49339\
        );

    \I__11629\ : InMux
    port map (
            O => \N__49404\,
            I => \N__49339\
        );

    \I__11628\ : InMux
    port map (
            O => \N__49403\,
            I => \N__49332\
        );

    \I__11627\ : InMux
    port map (
            O => \N__49402\,
            I => \N__49332\
        );

    \I__11626\ : InMux
    port map (
            O => \N__49401\,
            I => \N__49332\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__49394\,
            I => \N__49327\
        );

    \I__11624\ : Span12Mux_v
    port map (
            O => \N__49391\,
            I => \N__49327\
        );

    \I__11623\ : Span12Mux_h
    port map (
            O => \N__49388\,
            I => \N__49324\
        );

    \I__11622\ : Span4Mux_h
    port map (
            O => \N__49385\,
            I => \N__49317\
        );

    \I__11621\ : Span4Mux_h
    port map (
            O => \N__49380\,
            I => \N__49317\
        );

    \I__11620\ : Span4Mux_v
    port map (
            O => \N__49375\,
            I => \N__49317\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__49372\,
            I => \N__49310\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__49369\,
            I => \N__49310\
        );

    \I__11617\ : Sp12to4
    port map (
            O => \N__49362\,
            I => \N__49310\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__49353\,
            I => comm_state_0
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__49348\,
            I => comm_state_0
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__49339\,
            I => comm_state_0
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__49332\,
            I => comm_state_0
        );

    \I__11612\ : Odrv12
    port map (
            O => \N__49327\,
            I => comm_state_0
        );

    \I__11611\ : Odrv12
    port map (
            O => \N__49324\,
            I => comm_state_0
        );

    \I__11610\ : Odrv4
    port map (
            O => \N__49317\,
            I => comm_state_0
        );

    \I__11609\ : Odrv12
    port map (
            O => \N__49310\,
            I => comm_state_0
        );

    \I__11608\ : InMux
    port map (
            O => \N__49293\,
            I => \N__49289\
        );

    \I__11607\ : InMux
    port map (
            O => \N__49292\,
            I => \N__49286\
        );

    \I__11606\ : LocalMux
    port map (
            O => \N__49289\,
            I => n18991
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__49286\,
            I => n18991
        );

    \I__11604\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49272\
        );

    \I__11603\ : InMux
    port map (
            O => \N__49280\,
            I => \N__49272\
        );

    \I__11602\ : InMux
    port map (
            O => \N__49279\,
            I => \N__49272\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__49272\,
            I => \N__49268\
        );

    \I__11600\ : InMux
    port map (
            O => \N__49271\,
            I => \N__49265\
        );

    \I__11599\ : Span12Mux_h
    port map (
            O => \N__49268\,
            I => \N__49262\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__49265\,
            I => \N__49259\
        );

    \I__11597\ : Odrv12
    port map (
            O => \N__49262\,
            I => n20804
        );

    \I__11596\ : Odrv4
    port map (
            O => \N__49259\,
            I => n20804
        );

    \I__11595\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49251\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__49251\,
            I => \N__49248\
        );

    \I__11593\ : Span4Mux_v
    port map (
            O => \N__49248\,
            I => \N__49245\
        );

    \I__11592\ : Span4Mux_v
    port map (
            O => \N__49245\,
            I => \N__49242\
        );

    \I__11591\ : Odrv4
    port map (
            O => \N__49242\,
            I => n21341
        );

    \I__11590\ : CascadeMux
    port map (
            O => \N__49239\,
            I => \n21339_cascade_\
        );

    \I__11589\ : InMux
    port map (
            O => \N__49236\,
            I => \N__49233\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__49233\,
            I => n38_adj_1608
        );

    \I__11587\ : CascadeMux
    port map (
            O => \N__49230\,
            I => \N__49227\
        );

    \I__11586\ : InMux
    port map (
            O => \N__49227\,
            I => \N__49224\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__49224\,
            I => \N__49221\
        );

    \I__11584\ : Span4Mux_v
    port map (
            O => \N__49221\,
            I => \N__49218\
        );

    \I__11583\ : Odrv4
    port map (
            O => \N__49218\,
            I => n21054
        );

    \I__11582\ : InMux
    port map (
            O => \N__49215\,
            I => \ADC_VDC.genclk.n19723\
        );

    \I__11581\ : InMux
    port map (
            O => \N__49212\,
            I => \N__49208\
        );

    \I__11580\ : InMux
    port map (
            O => \N__49211\,
            I => \N__49205\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__49208\,
            I => \N__49202\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__49205\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__11577\ : Odrv4
    port map (
            O => \N__49202\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__11576\ : CEMux
    port map (
            O => \N__49197\,
            I => \N__49193\
        );

    \I__11575\ : CEMux
    port map (
            O => \N__49196\,
            I => \N__49190\
        );

    \I__11574\ : LocalMux
    port map (
            O => \N__49193\,
            I => \N__49187\
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__49190\,
            I => \N__49184\
        );

    \I__11572\ : Span4Mux_h
    port map (
            O => \N__49187\,
            I => \N__49181\
        );

    \I__11571\ : Odrv12
    port map (
            O => \N__49184\,
            I => \ADC_VDC.genclk.n11735\
        );

    \I__11570\ : Odrv4
    port map (
            O => \N__49181\,
            I => \ADC_VDC.genclk.n11735\
        );

    \I__11569\ : InMux
    port map (
            O => \N__49176\,
            I => \N__49173\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__49173\,
            I => \N__49168\
        );

    \I__11567\ : CascadeMux
    port map (
            O => \N__49172\,
            I => \N__49164\
        );

    \I__11566\ : InMux
    port map (
            O => \N__49171\,
            I => \N__49161\
        );

    \I__11565\ : Span4Mux_h
    port map (
            O => \N__49168\,
            I => \N__49158\
        );

    \I__11564\ : InMux
    port map (
            O => \N__49167\,
            I => \N__49155\
        );

    \I__11563\ : InMux
    port map (
            O => \N__49164\,
            I => \N__49152\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__49161\,
            I => n14529
        );

    \I__11561\ : Odrv4
    port map (
            O => \N__49158\,
            I => n14529
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__49155\,
            I => n14529
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__49152\,
            I => n14529
        );

    \I__11558\ : InMux
    port map (
            O => \N__49143\,
            I => \N__49140\
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__49140\,
            I => \N__49137\
        );

    \I__11556\ : Span4Mux_h
    port map (
            O => \N__49137\,
            I => \N__49134\
        );

    \I__11555\ : Span4Mux_h
    port map (
            O => \N__49134\,
            I => \N__49131\
        );

    \I__11554\ : Odrv4
    port map (
            O => \N__49131\,
            I => n17815
        );

    \I__11553\ : InMux
    port map (
            O => \N__49128\,
            I => \N__49125\
        );

    \I__11552\ : LocalMux
    port map (
            O => \N__49125\,
            I => \N__49122\
        );

    \I__11551\ : Span4Mux_v
    port map (
            O => \N__49122\,
            I => \N__49119\
        );

    \I__11550\ : Span4Mux_h
    port map (
            O => \N__49119\,
            I => \N__49116\
        );

    \I__11549\ : Odrv4
    port map (
            O => \N__49116\,
            I => n23_adj_1620
        );

    \I__11548\ : CascadeMux
    port map (
            O => \N__49113\,
            I => \n21_adj_1598_cascade_\
        );

    \I__11547\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49107\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__49107\,
            I => \N__49104\
        );

    \I__11545\ : Span4Mux_h
    port map (
            O => \N__49104\,
            I => \N__49101\
        );

    \I__11544\ : Span4Mux_h
    port map (
            O => \N__49101\,
            I => \N__49098\
        );

    \I__11543\ : Span4Mux_h
    port map (
            O => \N__49098\,
            I => \N__49095\
        );

    \I__11542\ : Odrv4
    port map (
            O => \N__49095\,
            I => n17564
        );

    \I__11541\ : InMux
    port map (
            O => \N__49092\,
            I => \N__49089\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__49089\,
            I => \N__49083\
        );

    \I__11539\ : InMux
    port map (
            O => \N__49088\,
            I => \N__49080\
        );

    \I__11538\ : InMux
    port map (
            O => \N__49087\,
            I => \N__49077\
        );

    \I__11537\ : InMux
    port map (
            O => \N__49086\,
            I => \N__49074\
        );

    \I__11536\ : Span4Mux_v
    port map (
            O => \N__49083\,
            I => \N__49071\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__49080\,
            I => \N__49068\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__49077\,
            I => \N__49063\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__49074\,
            I => \N__49063\
        );

    \I__11532\ : Span4Mux_h
    port map (
            O => \N__49071\,
            I => \N__49058\
        );

    \I__11531\ : Span4Mux_v
    port map (
            O => \N__49068\,
            I => \N__49058\
        );

    \I__11530\ : Span4Mux_h
    port map (
            O => \N__49063\,
            I => \N__49055\
        );

    \I__11529\ : Odrv4
    port map (
            O => \N__49058\,
            I => n2358
        );

    \I__11528\ : Odrv4
    port map (
            O => \N__49055\,
            I => n2358
        );

    \I__11527\ : InMux
    port map (
            O => \N__49050\,
            I => \N__49047\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__49047\,
            I => \N__49044\
        );

    \I__11525\ : Sp12to4
    port map (
            O => \N__49044\,
            I => \N__49041\
        );

    \I__11524\ : Span12Mux_h
    port map (
            O => \N__49041\,
            I => \N__49038\
        );

    \I__11523\ : Odrv12
    port map (
            O => \N__49038\,
            I => n20856
        );

    \I__11522\ : CascadeMux
    port map (
            O => \N__49035\,
            I => \n15_cascade_\
        );

    \I__11521\ : CEMux
    port map (
            O => \N__49032\,
            I => \N__49029\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__49029\,
            I => n18_adj_1619
        );

    \I__11519\ : CascadeMux
    port map (
            O => \N__49026\,
            I => \N__49023\
        );

    \I__11518\ : InMux
    port map (
            O => \N__49023\,
            I => \N__49020\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__49020\,
            I => n14130
        );

    \I__11516\ : InMux
    port map (
            O => \N__49017\,
            I => \N__49014\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__49014\,
            I => n20880
        );

    \I__11514\ : CascadeMux
    port map (
            O => \N__49011\,
            I => \n20880_cascade_\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__49008\,
            I => \N__49004\
        );

    \I__11512\ : InMux
    port map (
            O => \N__49007\,
            I => \N__49001\
        );

    \I__11511\ : InMux
    port map (
            O => \N__49004\,
            I => \N__48998\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__49001\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__11509\ : LocalMux
    port map (
            O => \N__48998\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__11508\ : InMux
    port map (
            O => \N__48993\,
            I => \ADC_VDC.genclk.n19715\
        );

    \I__11507\ : InMux
    port map (
            O => \N__48990\,
            I => \N__48986\
        );

    \I__11506\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48983\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__48986\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__11504\ : LocalMux
    port map (
            O => \N__48983\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__11503\ : InMux
    port map (
            O => \N__48978\,
            I => \bfn_19_8_0_\
        );

    \I__11502\ : CascadeMux
    port map (
            O => \N__48975\,
            I => \N__48971\
        );

    \I__11501\ : CascadeMux
    port map (
            O => \N__48974\,
            I => \N__48968\
        );

    \I__11500\ : InMux
    port map (
            O => \N__48971\,
            I => \N__48965\
        );

    \I__11499\ : InMux
    port map (
            O => \N__48968\,
            I => \N__48962\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__48965\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__48962\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__11496\ : InMux
    port map (
            O => \N__48957\,
            I => \ADC_VDC.genclk.n19717\
        );

    \I__11495\ : InMux
    port map (
            O => \N__48954\,
            I => \N__48950\
        );

    \I__11494\ : InMux
    port map (
            O => \N__48953\,
            I => \N__48947\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__48950\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__48947\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__11491\ : InMux
    port map (
            O => \N__48942\,
            I => \ADC_VDC.genclk.n19718\
        );

    \I__11490\ : CascadeMux
    port map (
            O => \N__48939\,
            I => \N__48936\
        );

    \I__11489\ : InMux
    port map (
            O => \N__48936\,
            I => \N__48932\
        );

    \I__11488\ : InMux
    port map (
            O => \N__48935\,
            I => \N__48929\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__48932\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__48929\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48924\,
            I => \ADC_VDC.genclk.n19719\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48921\,
            I => \N__48917\
        );

    \I__11483\ : InMux
    port map (
            O => \N__48920\,
            I => \N__48914\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__48917\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__48914\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__11480\ : InMux
    port map (
            O => \N__48909\,
            I => \ADC_VDC.genclk.n19720\
        );

    \I__11479\ : CascadeMux
    port map (
            O => \N__48906\,
            I => \N__48903\
        );

    \I__11478\ : InMux
    port map (
            O => \N__48903\,
            I => \N__48899\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48902\,
            I => \N__48896\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__48899\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__48896\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48891\,
            I => \ADC_VDC.genclk.n19721\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48888\,
            I => \N__48884\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48887\,
            I => \N__48881\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__48884\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__11470\ : LocalMux
    port map (
            O => \N__48881\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48876\,
            I => \ADC_VDC.genclk.n19722\
        );

    \I__11468\ : CascadeMux
    port map (
            O => \N__48873\,
            I => \N__48859\
        );

    \I__11467\ : CascadeMux
    port map (
            O => \N__48872\,
            I => \N__48856\
        );

    \I__11466\ : CascadeMux
    port map (
            O => \N__48871\,
            I => \N__48848\
        );

    \I__11465\ : CascadeMux
    port map (
            O => \N__48870\,
            I => \N__48840\
        );

    \I__11464\ : CascadeMux
    port map (
            O => \N__48869\,
            I => \N__48837\
        );

    \I__11463\ : InMux
    port map (
            O => \N__48868\,
            I => \N__48817\
        );

    \I__11462\ : InMux
    port map (
            O => \N__48867\,
            I => \N__48817\
        );

    \I__11461\ : InMux
    port map (
            O => \N__48866\,
            I => \N__48817\
        );

    \I__11460\ : InMux
    port map (
            O => \N__48865\,
            I => \N__48817\
        );

    \I__11459\ : InMux
    port map (
            O => \N__48864\,
            I => \N__48817\
        );

    \I__11458\ : InMux
    port map (
            O => \N__48863\,
            I => \N__48817\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48862\,
            I => \N__48817\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48859\,
            I => \N__48806\
        );

    \I__11455\ : InMux
    port map (
            O => \N__48856\,
            I => \N__48806\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48855\,
            I => \N__48806\
        );

    \I__11453\ : InMux
    port map (
            O => \N__48854\,
            I => \N__48806\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48853\,
            I => \N__48806\
        );

    \I__11451\ : CascadeMux
    port map (
            O => \N__48852\,
            I => \N__48801\
        );

    \I__11450\ : CascadeMux
    port map (
            O => \N__48851\,
            I => \N__48793\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48848\,
            I => \N__48787\
        );

    \I__11448\ : InMux
    port map (
            O => \N__48847\,
            I => \N__48787\
        );

    \I__11447\ : InMux
    port map (
            O => \N__48846\,
            I => \N__48779\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48845\,
            I => \N__48779\
        );

    \I__11445\ : CascadeMux
    port map (
            O => \N__48844\,
            I => \N__48775\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48843\,
            I => \N__48769\
        );

    \I__11443\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48764\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48837\,
            I => \N__48764\
        );

    \I__11441\ : CascadeMux
    port map (
            O => \N__48836\,
            I => \N__48761\
        );

    \I__11440\ : CascadeMux
    port map (
            O => \N__48835\,
            I => \N__48755\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48747\
        );

    \I__11438\ : InMux
    port map (
            O => \N__48833\,
            I => \N__48747\
        );

    \I__11437\ : InMux
    port map (
            O => \N__48832\,
            I => \N__48747\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48817\,
            I => \N__48742\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48806\,
            I => \N__48742\
        );

    \I__11434\ : InMux
    port map (
            O => \N__48805\,
            I => \N__48735\
        );

    \I__11433\ : InMux
    port map (
            O => \N__48804\,
            I => \N__48735\
        );

    \I__11432\ : InMux
    port map (
            O => \N__48801\,
            I => \N__48735\
        );

    \I__11431\ : InMux
    port map (
            O => \N__48800\,
            I => \N__48728\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48799\,
            I => \N__48728\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48798\,
            I => \N__48728\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48797\,
            I => \N__48721\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48796\,
            I => \N__48721\
        );

    \I__11426\ : InMux
    port map (
            O => \N__48793\,
            I => \N__48721\
        );

    \I__11425\ : InMux
    port map (
            O => \N__48792\,
            I => \N__48718\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__48787\,
            I => \N__48715\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48786\,
            I => \N__48710\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48785\,
            I => \N__48710\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48784\,
            I => \N__48706\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__48779\,
            I => \N__48703\
        );

    \I__11419\ : InMux
    port map (
            O => \N__48778\,
            I => \N__48696\
        );

    \I__11418\ : InMux
    port map (
            O => \N__48775\,
            I => \N__48696\
        );

    \I__11417\ : InMux
    port map (
            O => \N__48774\,
            I => \N__48696\
        );

    \I__11416\ : CascadeMux
    port map (
            O => \N__48773\,
            I => \N__48693\
        );

    \I__11415\ : CascadeMux
    port map (
            O => \N__48772\,
            I => \N__48690\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__48769\,
            I => \N__48684\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__48764\,
            I => \N__48684\
        );

    \I__11412\ : InMux
    port map (
            O => \N__48761\,
            I => \N__48681\
        );

    \I__11411\ : InMux
    port map (
            O => \N__48760\,
            I => \N__48678\
        );

    \I__11410\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48675\
        );

    \I__11409\ : InMux
    port map (
            O => \N__48758\,
            I => \N__48668\
        );

    \I__11408\ : InMux
    port map (
            O => \N__48755\,
            I => \N__48668\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48668\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48747\,
            I => \N__48657\
        );

    \I__11405\ : Span4Mux_v
    port map (
            O => \N__48742\,
            I => \N__48657\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48735\,
            I => \N__48657\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__48728\,
            I => \N__48657\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__48721\,
            I => \N__48657\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48718\,
            I => \N__48654\
        );

    \I__11400\ : Span4Mux_v
    port map (
            O => \N__48715\,
            I => \N__48651\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__48710\,
            I => \N__48648\
        );

    \I__11398\ : InMux
    port map (
            O => \N__48709\,
            I => \N__48645\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48706\,
            I => \N__48640\
        );

    \I__11396\ : Span4Mux_h
    port map (
            O => \N__48703\,
            I => \N__48640\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48696\,
            I => \N__48637\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48693\,
            I => \N__48634\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48690\,
            I => \N__48629\
        );

    \I__11392\ : InMux
    port map (
            O => \N__48689\,
            I => \N__48629\
        );

    \I__11391\ : Span12Mux_h
    port map (
            O => \N__48684\,
            I => \N__48626\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__48681\,
            I => \N__48613\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48613\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__48675\,
            I => \N__48613\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__48668\,
            I => \N__48613\
        );

    \I__11386\ : Span4Mux_v
    port map (
            O => \N__48657\,
            I => \N__48613\
        );

    \I__11385\ : Span4Mux_v
    port map (
            O => \N__48654\,
            I => \N__48613\
        );

    \I__11384\ : Sp12to4
    port map (
            O => \N__48651\,
            I => \N__48608\
        );

    \I__11383\ : Span12Mux_v
    port map (
            O => \N__48648\,
            I => \N__48608\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__48645\,
            I => adc_state_2
        );

    \I__11381\ : Odrv4
    port map (
            O => \N__48640\,
            I => adc_state_2
        );

    \I__11380\ : Odrv4
    port map (
            O => \N__48637\,
            I => adc_state_2
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__48634\,
            I => adc_state_2
        );

    \I__11378\ : LocalMux
    port map (
            O => \N__48629\,
            I => adc_state_2
        );

    \I__11377\ : Odrv12
    port map (
            O => \N__48626\,
            I => adc_state_2
        );

    \I__11376\ : Odrv4
    port map (
            O => \N__48613\,
            I => adc_state_2
        );

    \I__11375\ : Odrv12
    port map (
            O => \N__48608\,
            I => adc_state_2
        );

    \I__11374\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48570\
        );

    \I__11373\ : InMux
    port map (
            O => \N__48590\,
            I => \N__48570\
        );

    \I__11372\ : InMux
    port map (
            O => \N__48589\,
            I => \N__48539\
        );

    \I__11371\ : InMux
    port map (
            O => \N__48588\,
            I => \N__48539\
        );

    \I__11370\ : InMux
    port map (
            O => \N__48587\,
            I => \N__48539\
        );

    \I__11369\ : InMux
    port map (
            O => \N__48586\,
            I => \N__48539\
        );

    \I__11368\ : InMux
    port map (
            O => \N__48585\,
            I => \N__48539\
        );

    \I__11367\ : InMux
    port map (
            O => \N__48584\,
            I => \N__48539\
        );

    \I__11366\ : InMux
    port map (
            O => \N__48583\,
            I => \N__48539\
        );

    \I__11365\ : InMux
    port map (
            O => \N__48582\,
            I => \N__48539\
        );

    \I__11364\ : InMux
    port map (
            O => \N__48581\,
            I => \N__48531\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48580\,
            I => \N__48531\
        );

    \I__11362\ : InMux
    port map (
            O => \N__48579\,
            I => \N__48517\
        );

    \I__11361\ : InMux
    port map (
            O => \N__48578\,
            I => \N__48517\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48577\,
            I => \N__48517\
        );

    \I__11359\ : InMux
    port map (
            O => \N__48576\,
            I => \N__48517\
        );

    \I__11358\ : InMux
    port map (
            O => \N__48575\,
            I => \N__48517\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__48570\,
            I => \N__48514\
        );

    \I__11356\ : InMux
    port map (
            O => \N__48569\,
            I => \N__48509\
        );

    \I__11355\ : InMux
    port map (
            O => \N__48568\,
            I => \N__48509\
        );

    \I__11354\ : InMux
    port map (
            O => \N__48567\,
            I => \N__48502\
        );

    \I__11353\ : InMux
    port map (
            O => \N__48566\,
            I => \N__48502\
        );

    \I__11352\ : InMux
    port map (
            O => \N__48565\,
            I => \N__48502\
        );

    \I__11351\ : InMux
    port map (
            O => \N__48564\,
            I => \N__48497\
        );

    \I__11350\ : InMux
    port map (
            O => \N__48563\,
            I => \N__48497\
        );

    \I__11349\ : InMux
    port map (
            O => \N__48562\,
            I => \N__48482\
        );

    \I__11348\ : InMux
    port map (
            O => \N__48561\,
            I => \N__48482\
        );

    \I__11347\ : InMux
    port map (
            O => \N__48560\,
            I => \N__48482\
        );

    \I__11346\ : InMux
    port map (
            O => \N__48559\,
            I => \N__48482\
        );

    \I__11345\ : InMux
    port map (
            O => \N__48558\,
            I => \N__48482\
        );

    \I__11344\ : InMux
    port map (
            O => \N__48557\,
            I => \N__48482\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48556\,
            I => \N__48482\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__48539\,
            I => \N__48476\
        );

    \I__11341\ : InMux
    port map (
            O => \N__48538\,
            I => \N__48473\
        );

    \I__11340\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48470\
        );

    \I__11339\ : InMux
    port map (
            O => \N__48536\,
            I => \N__48467\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__48531\,
            I => \N__48461\
        );

    \I__11337\ : InMux
    port map (
            O => \N__48530\,
            I => \N__48458\
        );

    \I__11336\ : CascadeMux
    port map (
            O => \N__48529\,
            I => \N__48452\
        );

    \I__11335\ : InMux
    port map (
            O => \N__48528\,
            I => \N__48449\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__48517\,
            I => \N__48444\
        );

    \I__11333\ : Span4Mux_v
    port map (
            O => \N__48514\,
            I => \N__48444\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__48509\,
            I => \N__48441\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__48502\,
            I => \N__48434\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__48497\,
            I => \N__48434\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__48482\,
            I => \N__48434\
        );

    \I__11328\ : InMux
    port map (
            O => \N__48481\,
            I => \N__48431\
        );

    \I__11327\ : InMux
    port map (
            O => \N__48480\,
            I => \N__48426\
        );

    \I__11326\ : InMux
    port map (
            O => \N__48479\,
            I => \N__48426\
        );

    \I__11325\ : Span4Mux_h
    port map (
            O => \N__48476\,
            I => \N__48419\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__48473\,
            I => \N__48419\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__48470\,
            I => \N__48419\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__48467\,
            I => \N__48416\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48466\,
            I => \N__48409\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48409\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48464\,
            I => \N__48409\
        );

    \I__11318\ : Span4Mux_v
    port map (
            O => \N__48461\,
            I => \N__48406\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__48458\,
            I => \N__48403\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48457\,
            I => \N__48400\
        );

    \I__11315\ : InMux
    port map (
            O => \N__48456\,
            I => \N__48393\
        );

    \I__11314\ : InMux
    port map (
            O => \N__48455\,
            I => \N__48393\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48452\,
            I => \N__48393\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__48449\,
            I => \N__48384\
        );

    \I__11311\ : Span4Mux_v
    port map (
            O => \N__48444\,
            I => \N__48384\
        );

    \I__11310\ : Span4Mux_v
    port map (
            O => \N__48441\,
            I => \N__48384\
        );

    \I__11309\ : Span4Mux_v
    port map (
            O => \N__48434\,
            I => \N__48384\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__48431\,
            I => \N__48371\
        );

    \I__11307\ : LocalMux
    port map (
            O => \N__48426\,
            I => \N__48371\
        );

    \I__11306\ : Span4Mux_v
    port map (
            O => \N__48419\,
            I => \N__48371\
        );

    \I__11305\ : Span4Mux_v
    port map (
            O => \N__48416\,
            I => \N__48371\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__48409\,
            I => \N__48371\
        );

    \I__11303\ : Span4Mux_h
    port map (
            O => \N__48406\,
            I => \N__48371\
        );

    \I__11302\ : Odrv4
    port map (
            O => \N__48403\,
            I => adc_state_3
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__48400\,
            I => adc_state_3
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__48393\,
            I => adc_state_3
        );

    \I__11299\ : Odrv4
    port map (
            O => \N__48384\,
            I => adc_state_3
        );

    \I__11298\ : Odrv4
    port map (
            O => \N__48371\,
            I => adc_state_3
        );

    \I__11297\ : CascadeMux
    port map (
            O => \N__48360\,
            I => \ADC_VDC.n62_cascade_\
        );

    \I__11296\ : CascadeMux
    port map (
            O => \N__48357\,
            I => \N__48351\
        );

    \I__11295\ : InMux
    port map (
            O => \N__48356\,
            I => \N__48340\
        );

    \I__11294\ : InMux
    port map (
            O => \N__48355\,
            I => \N__48340\
        );

    \I__11293\ : InMux
    port map (
            O => \N__48354\,
            I => \N__48331\
        );

    \I__11292\ : InMux
    port map (
            O => \N__48351\,
            I => \N__48331\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48350\,
            I => \N__48331\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48349\,
            I => \N__48328\
        );

    \I__11289\ : InMux
    port map (
            O => \N__48348\,
            I => \N__48323\
        );

    \I__11288\ : InMux
    port map (
            O => \N__48347\,
            I => \N__48323\
        );

    \I__11287\ : InMux
    port map (
            O => \N__48346\,
            I => \N__48320\
        );

    \I__11286\ : InMux
    port map (
            O => \N__48345\,
            I => \N__48317\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__48340\,
            I => \N__48314\
        );

    \I__11284\ : InMux
    port map (
            O => \N__48339\,
            I => \N__48309\
        );

    \I__11283\ : InMux
    port map (
            O => \N__48338\,
            I => \N__48309\
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__48331\,
            I => \N__48306\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__48328\,
            I => \N__48301\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__48323\,
            I => \N__48301\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__48320\,
            I => \N__48292\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__48317\,
            I => \N__48292\
        );

    \I__11277\ : Span4Mux_v
    port map (
            O => \N__48314\,
            I => \N__48289\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__48309\,
            I => \N__48280\
        );

    \I__11275\ : Span4Mux_v
    port map (
            O => \N__48306\,
            I => \N__48280\
        );

    \I__11274\ : Span4Mux_v
    port map (
            O => \N__48301\,
            I => \N__48280\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48300\,
            I => \N__48272\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48269\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48298\,
            I => \N__48266\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48297\,
            I => \N__48263\
        );

    \I__11269\ : Span4Mux_v
    port map (
            O => \N__48292\,
            I => \N__48258\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__48289\,
            I => \N__48258\
        );

    \I__11267\ : InMux
    port map (
            O => \N__48288\,
            I => \N__48253\
        );

    \I__11266\ : InMux
    port map (
            O => \N__48287\,
            I => \N__48253\
        );

    \I__11265\ : Span4Mux_h
    port map (
            O => \N__48280\,
            I => \N__48250\
        );

    \I__11264\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48245\
        );

    \I__11263\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48245\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48277\,
            I => \N__48238\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48276\,
            I => \N__48238\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48275\,
            I => \N__48238\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48272\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__48269\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__48266\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__48263\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11255\ : Odrv4
    port map (
            O => \N__48258\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__48253\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11253\ : Odrv4
    port map (
            O => \N__48250\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__48245\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__48238\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__11250\ : InMux
    port map (
            O => \N__48219\,
            I => \N__48216\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48216\,
            I => \N__48213\
        );

    \I__11248\ : Span4Mux_h
    port map (
            O => \N__48213\,
            I => \N__48210\
        );

    \I__11247\ : Odrv4
    port map (
            O => \N__48210\,
            I => \ADC_VDC.n11\
        );

    \I__11246\ : InMux
    port map (
            O => \N__48207\,
            I => \N__48203\
        );

    \I__11245\ : InMux
    port map (
            O => \N__48206\,
            I => \N__48200\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__48203\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__48200\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__11242\ : InMux
    port map (
            O => \N__48195\,
            I => \bfn_19_7_0_\
        );

    \I__11241\ : InMux
    port map (
            O => \N__48192\,
            I => \N__48188\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48185\
        );

    \I__11239\ : LocalMux
    port map (
            O => \N__48188\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__48185\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48180\,
            I => \ADC_VDC.genclk.n19709\
        );

    \I__11236\ : CascadeMux
    port map (
            O => \N__48177\,
            I => \N__48174\
        );

    \I__11235\ : InMux
    port map (
            O => \N__48174\,
            I => \N__48170\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48173\,
            I => \N__48167\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__48170\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__48167\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__11231\ : InMux
    port map (
            O => \N__48162\,
            I => \ADC_VDC.genclk.n19710\
        );

    \I__11230\ : InMux
    port map (
            O => \N__48159\,
            I => \N__48155\
        );

    \I__11229\ : InMux
    port map (
            O => \N__48158\,
            I => \N__48152\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__48155\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__48152\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__11226\ : InMux
    port map (
            O => \N__48147\,
            I => \ADC_VDC.genclk.n19711\
        );

    \I__11225\ : CascadeMux
    port map (
            O => \N__48144\,
            I => \N__48140\
        );

    \I__11224\ : CascadeMux
    port map (
            O => \N__48143\,
            I => \N__48137\
        );

    \I__11223\ : InMux
    port map (
            O => \N__48140\,
            I => \N__48134\
        );

    \I__11222\ : InMux
    port map (
            O => \N__48137\,
            I => \N__48131\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__48134\,
            I => \N__48128\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48131\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__11219\ : Odrv4
    port map (
            O => \N__48128\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__11218\ : InMux
    port map (
            O => \N__48123\,
            I => \ADC_VDC.genclk.n19712\
        );

    \I__11217\ : CascadeMux
    port map (
            O => \N__48120\,
            I => \N__48116\
        );

    \I__11216\ : InMux
    port map (
            O => \N__48119\,
            I => \N__48113\
        );

    \I__11215\ : InMux
    port map (
            O => \N__48116\,
            I => \N__48110\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__48113\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__48110\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__11212\ : InMux
    port map (
            O => \N__48105\,
            I => \ADC_VDC.genclk.n19713\
        );

    \I__11211\ : CascadeMux
    port map (
            O => \N__48102\,
            I => \N__48099\
        );

    \I__11210\ : InMux
    port map (
            O => \N__48099\,
            I => \N__48095\
        );

    \I__11209\ : InMux
    port map (
            O => \N__48098\,
            I => \N__48092\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__48095\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__48092\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__11206\ : InMux
    port map (
            O => \N__48087\,
            I => \ADC_VDC.genclk.n19714\
        );

    \I__11205\ : InMux
    port map (
            O => \N__48084\,
            I => \N__48081\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__48081\,
            I => \N__48077\
        );

    \I__11203\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48074\
        );

    \I__11202\ : Span4Mux_v
    port map (
            O => \N__48077\,
            I => \N__48069\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__48074\,
            I => \N__48069\
        );

    \I__11200\ : Span4Mux_h
    port map (
            O => \N__48069\,
            I => \N__48063\
        );

    \I__11199\ : InMux
    port map (
            O => \N__48068\,
            I => \N__48060\
        );

    \I__11198\ : CascadeMux
    port map (
            O => \N__48067\,
            I => \N__48056\
        );

    \I__11197\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48053\
        );

    \I__11196\ : Span4Mux_v
    port map (
            O => \N__48063\,
            I => \N__48048\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__48060\,
            I => \N__48048\
        );

    \I__11194\ : InMux
    port map (
            O => \N__48059\,
            I => \N__48045\
        );

    \I__11193\ : InMux
    port map (
            O => \N__48056\,
            I => \N__48042\
        );

    \I__11192\ : LocalMux
    port map (
            O => \N__48053\,
            I => \N__48035\
        );

    \I__11191\ : Span4Mux_v
    port map (
            O => \N__48048\,
            I => \N__48035\
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__48045\,
            I => \N__48035\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__48042\,
            I => \N__48030\
        );

    \I__11188\ : Span4Mux_h
    port map (
            O => \N__48035\,
            I => \N__48030\
        );

    \I__11187\ : Odrv4
    port map (
            O => \N__48030\,
            I => comm_buf_1_2
        );

    \I__11186\ : InMux
    port map (
            O => \N__48027\,
            I => \N__48021\
        );

    \I__11185\ : InMux
    port map (
            O => \N__48026\,
            I => \N__48018\
        );

    \I__11184\ : InMux
    port map (
            O => \N__48025\,
            I => \N__48013\
        );

    \I__11183\ : InMux
    port map (
            O => \N__48024\,
            I => \N__48013\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__48021\,
            I => \N__48006\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__48018\,
            I => \N__48001\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__48013\,
            I => \N__48001\
        );

    \I__11179\ : InMux
    port map (
            O => \N__48012\,
            I => \N__47998\
        );

    \I__11178\ : InMux
    port map (
            O => \N__48011\,
            I => \N__47992\
        );

    \I__11177\ : InMux
    port map (
            O => \N__48010\,
            I => \N__47987\
        );

    \I__11176\ : InMux
    port map (
            O => \N__48009\,
            I => \N__47987\
        );

    \I__11175\ : Span4Mux_v
    port map (
            O => \N__48006\,
            I => \N__47981\
        );

    \I__11174\ : Span4Mux_v
    port map (
            O => \N__48001\,
            I => \N__47981\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__47998\,
            I => \N__47978\
        );

    \I__11172\ : InMux
    port map (
            O => \N__47997\,
            I => \N__47975\
        );

    \I__11171\ : InMux
    port map (
            O => \N__47996\,
            I => \N__47970\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47995\,
            I => \N__47970\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__47992\,
            I => \N__47964\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__47987\,
            I => \N__47961\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47986\,
            I => \N__47958\
        );

    \I__11166\ : Span4Mux_h
    port map (
            O => \N__47981\,
            I => \N__47951\
        );

    \I__11165\ : Span4Mux_v
    port map (
            O => \N__47978\,
            I => \N__47951\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__47975\,
            I => \N__47951\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__47970\,
            I => \N__47948\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47969\,
            I => \N__47941\
        );

    \I__11161\ : InMux
    port map (
            O => \N__47968\,
            I => \N__47941\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47941\
        );

    \I__11159\ : Odrv12
    port map (
            O => \N__47964\,
            I => n12367
        );

    \I__11158\ : Odrv12
    port map (
            O => \N__47961\,
            I => n12367
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__47958\,
            I => n12367
        );

    \I__11156\ : Odrv4
    port map (
            O => \N__47951\,
            I => n12367
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__47948\,
            I => n12367
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__47941\,
            I => n12367
        );

    \I__11153\ : CascadeMux
    port map (
            O => \N__47928\,
            I => \N__47925\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47922\
        );

    \I__11151\ : LocalMux
    port map (
            O => \N__47922\,
            I => \N__47919\
        );

    \I__11150\ : Span4Mux_v
    port map (
            O => \N__47919\,
            I => \N__47916\
        );

    \I__11149\ : Span4Mux_h
    port map (
            O => \N__47916\,
            I => \N__47911\
        );

    \I__11148\ : InMux
    port map (
            O => \N__47915\,
            I => \N__47906\
        );

    \I__11147\ : InMux
    port map (
            O => \N__47914\,
            I => \N__47906\
        );

    \I__11146\ : Odrv4
    port map (
            O => \N__47911\,
            I => buf_dds0_2
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__47906\,
            I => buf_dds0_2
        );

    \I__11144\ : CascadeMux
    port map (
            O => \N__47901\,
            I => \N__47898\
        );

    \I__11143\ : InMux
    port map (
            O => \N__47898\,
            I => \N__47892\
        );

    \I__11142\ : CascadeMux
    port map (
            O => \N__47897\,
            I => \N__47888\
        );

    \I__11141\ : CascadeMux
    port map (
            O => \N__47896\,
            I => \N__47885\
        );

    \I__11140\ : InMux
    port map (
            O => \N__47895\,
            I => \N__47882\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__47892\,
            I => \N__47879\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47891\,
            I => \N__47875\
        );

    \I__11137\ : InMux
    port map (
            O => \N__47888\,
            I => \N__47872\
        );

    \I__11136\ : InMux
    port map (
            O => \N__47885\,
            I => \N__47869\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47866\
        );

    \I__11134\ : Span4Mux_h
    port map (
            O => \N__47879\,
            I => \N__47863\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47878\,
            I => \N__47860\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__47875\,
            I => \N__47857\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__47872\,
            I => \N__47850\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47869\,
            I => \N__47850\
        );

    \I__11129\ : Span4Mux_v
    port map (
            O => \N__47866\,
            I => \N__47850\
        );

    \I__11128\ : Span4Mux_v
    port map (
            O => \N__47863\,
            I => \N__47847\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__47860\,
            I => \N__47844\
        );

    \I__11126\ : Span4Mux_v
    port map (
            O => \N__47857\,
            I => \N__47839\
        );

    \I__11125\ : Span4Mux_h
    port map (
            O => \N__47850\,
            I => \N__47839\
        );

    \I__11124\ : Odrv4
    port map (
            O => \N__47847\,
            I => comm_buf_1_6
        );

    \I__11123\ : Odrv12
    port map (
            O => \N__47844\,
            I => comm_buf_1_6
        );

    \I__11122\ : Odrv4
    port map (
            O => \N__47839\,
            I => comm_buf_1_6
        );

    \I__11121\ : InMux
    port map (
            O => \N__47832\,
            I => \N__47829\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47829\,
            I => \N__47825\
        );

    \I__11119\ : InMux
    port map (
            O => \N__47828\,
            I => \N__47822\
        );

    \I__11118\ : Span4Mux_v
    port map (
            O => \N__47825\,
            I => \N__47819\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__47822\,
            I => \N__47816\
        );

    \I__11116\ : Span4Mux_h
    port map (
            O => \N__47819\,
            I => \N__47813\
        );

    \I__11115\ : Span4Mux_h
    port map (
            O => \N__47816\,
            I => \N__47810\
        );

    \I__11114\ : Odrv4
    port map (
            O => \N__47813\,
            I => n14_adj_1552
        );

    \I__11113\ : Odrv4
    port map (
            O => \N__47810\,
            I => n14_adj_1552
        );

    \I__11112\ : CascadeMux
    port map (
            O => \N__47805\,
            I => \N__47802\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47798\
        );

    \I__11110\ : CascadeMux
    port map (
            O => \N__47801\,
            I => \N__47795\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__47798\,
            I => \N__47791\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47795\,
            I => \N__47788\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47794\,
            I => \N__47785\
        );

    \I__11106\ : Span4Mux_h
    port map (
            O => \N__47791\,
            I => \N__47778\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__47788\,
            I => \N__47778\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47785\,
            I => \N__47775\
        );

    \I__11103\ : CascadeMux
    port map (
            O => \N__47784\,
            I => \N__47772\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47769\
        );

    \I__11101\ : Span4Mux_v
    port map (
            O => \N__47778\,
            I => \N__47764\
        );

    \I__11100\ : Span4Mux_h
    port map (
            O => \N__47775\,
            I => \N__47764\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47772\,
            I => \N__47760\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__47769\,
            I => \N__47757\
        );

    \I__11097\ : Span4Mux_h
    port map (
            O => \N__47764\,
            I => \N__47754\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47763\,
            I => \N__47751\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__47760\,
            I => \N__47748\
        );

    \I__11094\ : Span4Mux_h
    port map (
            O => \N__47757\,
            I => \N__47745\
        );

    \I__11093\ : Span4Mux_h
    port map (
            O => \N__47754\,
            I => \N__47740\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__47751\,
            I => \N__47740\
        );

    \I__11091\ : Span4Mux_h
    port map (
            O => \N__47748\,
            I => \N__47737\
        );

    \I__11090\ : Span4Mux_v
    port map (
            O => \N__47745\,
            I => \N__47732\
        );

    \I__11089\ : Span4Mux_v
    port map (
            O => \N__47740\,
            I => \N__47732\
        );

    \I__11088\ : Odrv4
    port map (
            O => \N__47737\,
            I => comm_buf_1_4
        );

    \I__11087\ : Odrv4
    port map (
            O => \N__47732\,
            I => comm_buf_1_4
        );

    \I__11086\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47724\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47724\,
            I => \N__47719\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47716\
        );

    \I__11083\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47713\
        );

    \I__11082\ : Span12Mux_s10_h
    port map (
            O => \N__47719\,
            I => \N__47706\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__47716\,
            I => \N__47706\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__47713\,
            I => \N__47706\
        );

    \I__11079\ : Odrv12
    port map (
            O => \N__47706\,
            I => data_index_4
        );

    \I__11078\ : InMux
    port map (
            O => \N__47703\,
            I => \N__47698\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47702\,
            I => \N__47695\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47692\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__47698\,
            I => \N__47684\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47695\,
            I => \N__47684\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__47692\,
            I => \N__47677\
        );

    \I__11072\ : InMux
    port map (
            O => \N__47691\,
            I => \N__47674\
        );

    \I__11071\ : InMux
    port map (
            O => \N__47690\,
            I => \N__47669\
        );

    \I__11070\ : InMux
    port map (
            O => \N__47689\,
            I => \N__47669\
        );

    \I__11069\ : Span4Mux_h
    port map (
            O => \N__47684\,
            I => \N__47666\
        );

    \I__11068\ : InMux
    port map (
            O => \N__47683\,
            I => \N__47663\
        );

    \I__11067\ : InMux
    port map (
            O => \N__47682\,
            I => \N__47656\
        );

    \I__11066\ : InMux
    port map (
            O => \N__47681\,
            I => \N__47656\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47680\,
            I => \N__47656\
        );

    \I__11064\ : Span4Mux_v
    port map (
            O => \N__47677\,
            I => \N__47651\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__47674\,
            I => \N__47651\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__47669\,
            I => n8813
        );

    \I__11061\ : Odrv4
    port map (
            O => \N__47666\,
            I => n8813
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__47663\,
            I => n8813
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__47656\,
            I => n8813
        );

    \I__11058\ : Odrv4
    port map (
            O => \N__47651\,
            I => n8813
        );

    \I__11057\ : InMux
    port map (
            O => \N__47640\,
            I => \N__47637\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__47637\,
            I => \N__47634\
        );

    \I__11055\ : Span12Mux_h
    port map (
            O => \N__47634\,
            I => \N__47630\
        );

    \I__11054\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47627\
        );

    \I__11053\ : Odrv12
    port map (
            O => \N__47630\,
            I => n8_adj_1567
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__47627\,
            I => n8_adj_1567
        );

    \I__11051\ : InMux
    port map (
            O => \N__47622\,
            I => \N__47618\
        );

    \I__11050\ : InMux
    port map (
            O => \N__47621\,
            I => \N__47615\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__47618\,
            I => \N__47612\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47615\,
            I => \N__47609\
        );

    \I__11047\ : Span4Mux_h
    port map (
            O => \N__47612\,
            I => \N__47604\
        );

    \I__11046\ : Span4Mux_v
    port map (
            O => \N__47609\,
            I => \N__47604\
        );

    \I__11045\ : Odrv4
    port map (
            O => \N__47604\,
            I => n7_adj_1566
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__47601\,
            I => \N__47598\
        );

    \I__11043\ : CascadeBuf
    port map (
            O => \N__47598\,
            I => \N__47595\
        );

    \I__11042\ : CascadeMux
    port map (
            O => \N__47595\,
            I => \N__47592\
        );

    \I__11041\ : CascadeBuf
    port map (
            O => \N__47592\,
            I => \N__47589\
        );

    \I__11040\ : CascadeMux
    port map (
            O => \N__47589\,
            I => \N__47586\
        );

    \I__11039\ : CascadeBuf
    port map (
            O => \N__47586\,
            I => \N__47583\
        );

    \I__11038\ : CascadeMux
    port map (
            O => \N__47583\,
            I => \N__47580\
        );

    \I__11037\ : CascadeBuf
    port map (
            O => \N__47580\,
            I => \N__47577\
        );

    \I__11036\ : CascadeMux
    port map (
            O => \N__47577\,
            I => \N__47574\
        );

    \I__11035\ : CascadeBuf
    port map (
            O => \N__47574\,
            I => \N__47571\
        );

    \I__11034\ : CascadeMux
    port map (
            O => \N__47571\,
            I => \N__47568\
        );

    \I__11033\ : CascadeBuf
    port map (
            O => \N__47568\,
            I => \N__47565\
        );

    \I__11032\ : CascadeMux
    port map (
            O => \N__47565\,
            I => \N__47561\
        );

    \I__11031\ : CascadeMux
    port map (
            O => \N__47564\,
            I => \N__47558\
        );

    \I__11030\ : CascadeBuf
    port map (
            O => \N__47561\,
            I => \N__47555\
        );

    \I__11029\ : CascadeBuf
    port map (
            O => \N__47558\,
            I => \N__47552\
        );

    \I__11028\ : CascadeMux
    port map (
            O => \N__47555\,
            I => \N__47549\
        );

    \I__11027\ : CascadeMux
    port map (
            O => \N__47552\,
            I => \N__47546\
        );

    \I__11026\ : CascadeBuf
    port map (
            O => \N__47549\,
            I => \N__47543\
        );

    \I__11025\ : InMux
    port map (
            O => \N__47546\,
            I => \N__47540\
        );

    \I__11024\ : CascadeMux
    port map (
            O => \N__47543\,
            I => \N__47537\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__47540\,
            I => \N__47534\
        );

    \I__11022\ : CascadeBuf
    port map (
            O => \N__47537\,
            I => \N__47531\
        );

    \I__11021\ : Sp12to4
    port map (
            O => \N__47534\,
            I => \N__47528\
        );

    \I__11020\ : CascadeMux
    port map (
            O => \N__47531\,
            I => \N__47525\
        );

    \I__11019\ : Span12Mux_v
    port map (
            O => \N__47528\,
            I => \N__47522\
        );

    \I__11018\ : InMux
    port map (
            O => \N__47525\,
            I => \N__47519\
        );

    \I__11017\ : Span12Mux_h
    port map (
            O => \N__47522\,
            I => \N__47516\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__47519\,
            I => \N__47513\
        );

    \I__11015\ : Odrv12
    port map (
            O => \N__47516\,
            I => \data_index_9_N_216_4\
        );

    \I__11014\ : Odrv4
    port map (
            O => \N__47513\,
            I => \data_index_9_N_216_4\
        );

    \I__11013\ : CEMux
    port map (
            O => \N__47508\,
            I => \N__47505\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__47505\,
            I => \N__47502\
        );

    \I__11011\ : Span4Mux_h
    port map (
            O => \N__47502\,
            I => \N__47499\
        );

    \I__11010\ : Span4Mux_h
    port map (
            O => \N__47499\,
            I => \N__47496\
        );

    \I__11009\ : Odrv4
    port map (
            O => \N__47496\,
            I => \ADC_VDC.n11750\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47493\,
            I => \N__47486\
        );

    \I__11007\ : CascadeMux
    port map (
            O => \N__47492\,
            I => \N__47483\
        );

    \I__11006\ : CascadeMux
    port map (
            O => \N__47491\,
            I => \N__47477\
        );

    \I__11005\ : CascadeMux
    port map (
            O => \N__47490\,
            I => \N__47474\
        );

    \I__11004\ : CascadeMux
    port map (
            O => \N__47489\,
            I => \N__47470\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__47486\,
            I => \N__47467\
        );

    \I__11002\ : InMux
    port map (
            O => \N__47483\,
            I => \N__47464\
        );

    \I__11001\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47461\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47481\,
            I => \N__47456\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47480\,
            I => \N__47456\
        );

    \I__10998\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47453\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47474\,
            I => \N__47448\
        );

    \I__10996\ : InMux
    port map (
            O => \N__47473\,
            I => \N__47448\
        );

    \I__10995\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47445\
        );

    \I__10994\ : Span4Mux_v
    port map (
            O => \N__47467\,
            I => \N__47442\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__47464\,
            I => \N__47439\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__47461\,
            I => \N__47436\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__47456\,
            I => \N__47427\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__47453\,
            I => \N__47427\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__47448\,
            I => \N__47427\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__47445\,
            I => \N__47427\
        );

    \I__10987\ : Span4Mux_h
    port map (
            O => \N__47442\,
            I => \N__47419\
        );

    \I__10986\ : Span4Mux_v
    port map (
            O => \N__47439\,
            I => \N__47419\
        );

    \I__10985\ : Span4Mux_v
    port map (
            O => \N__47436\,
            I => \N__47419\
        );

    \I__10984\ : Span4Mux_v
    port map (
            O => \N__47427\,
            I => \N__47416\
        );

    \I__10983\ : CascadeMux
    port map (
            O => \N__47426\,
            I => \N__47413\
        );

    \I__10982\ : Span4Mux_v
    port map (
            O => \N__47419\,
            I => \N__47410\
        );

    \I__10981\ : Span4Mux_v
    port map (
            O => \N__47416\,
            I => \N__47407\
        );

    \I__10980\ : InMux
    port map (
            O => \N__47413\,
            I => \N__47404\
        );

    \I__10979\ : Sp12to4
    port map (
            O => \N__47410\,
            I => \N__47401\
        );

    \I__10978\ : Span4Mux_h
    port map (
            O => \N__47407\,
            I => \N__47398\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__47404\,
            I => \N__47395\
        );

    \I__10976\ : Span12Mux_h
    port map (
            O => \N__47401\,
            I => \N__47388\
        );

    \I__10975\ : Sp12to4
    port map (
            O => \N__47398\,
            I => \N__47388\
        );

    \I__10974\ : Span12Mux_v
    port map (
            O => \N__47395\,
            I => \N__47388\
        );

    \I__10973\ : Odrv12
    port map (
            O => \N__47388\,
            I => \VDC_SDO\
        );

    \I__10972\ : InMux
    port map (
            O => \N__47385\,
            I => \N__47378\
        );

    \I__10971\ : InMux
    port map (
            O => \N__47384\,
            I => \N__47378\
        );

    \I__10970\ : InMux
    port map (
            O => \N__47383\,
            I => \N__47374\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__47378\,
            I => \N__47371\
        );

    \I__10968\ : InMux
    port map (
            O => \N__47377\,
            I => \N__47368\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__47374\,
            I => \N__47352\
        );

    \I__10966\ : Span4Mux_v
    port map (
            O => \N__47371\,
            I => \N__47352\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47349\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47367\,
            I => \N__47344\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47366\,
            I => \N__47341\
        );

    \I__10962\ : InMux
    port map (
            O => \N__47365\,
            I => \N__47336\
        );

    \I__10961\ : InMux
    port map (
            O => \N__47364\,
            I => \N__47336\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47363\,
            I => \N__47329\
        );

    \I__10959\ : InMux
    port map (
            O => \N__47362\,
            I => \N__47322\
        );

    \I__10958\ : InMux
    port map (
            O => \N__47361\,
            I => \N__47322\
        );

    \I__10957\ : InMux
    port map (
            O => \N__47360\,
            I => \N__47322\
        );

    \I__10956\ : InMux
    port map (
            O => \N__47359\,
            I => \N__47317\
        );

    \I__10955\ : InMux
    port map (
            O => \N__47358\,
            I => \N__47317\
        );

    \I__10954\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47314\
        );

    \I__10953\ : Span4Mux_h
    port map (
            O => \N__47352\,
            I => \N__47309\
        );

    \I__10952\ : Span4Mux_h
    port map (
            O => \N__47349\,
            I => \N__47309\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47348\,
            I => \N__47304\
        );

    \I__10950\ : InMux
    port map (
            O => \N__47347\,
            I => \N__47304\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__47344\,
            I => \N__47297\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__47341\,
            I => \N__47297\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__47336\,
            I => \N__47297\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47335\,
            I => \N__47290\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47334\,
            I => \N__47290\
        );

    \I__10944\ : InMux
    port map (
            O => \N__47333\,
            I => \N__47290\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47332\,
            I => \N__47287\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__47329\,
            I => \N__47284\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__47322\,
            I => \N__47279\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__47317\,
            I => \N__47279\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__47314\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10938\ : Odrv4
    port map (
            O => \N__47309\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__47304\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10936\ : Odrv12
    port map (
            O => \N__47297\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__47290\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__47287\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10933\ : Odrv12
    port map (
            O => \N__47284\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10932\ : Odrv4
    port map (
            O => \N__47279\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__10931\ : CascadeMux
    port map (
            O => \N__47262\,
            I => \N__47259\
        );

    \I__10930\ : InMux
    port map (
            O => \N__47259\,
            I => \N__47256\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__47256\,
            I => \ADC_VDC.n62\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47250\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__47250\,
            I => n22210
        );

    \I__10926\ : CascadeMux
    port map (
            O => \N__47247\,
            I => \n22432_cascade_\
        );

    \I__10925\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47240\
        );

    \I__10924\ : InMux
    port map (
            O => \N__47243\,
            I => \N__47237\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__47240\,
            I => \N__47233\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__47237\,
            I => \N__47228\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47236\,
            I => \N__47225\
        );

    \I__10920\ : Span4Mux_v
    port map (
            O => \N__47233\,
            I => \N__47220\
        );

    \I__10919\ : InMux
    port map (
            O => \N__47232\,
            I => \N__47217\
        );

    \I__10918\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47214\
        );

    \I__10917\ : Span4Mux_v
    port map (
            O => \N__47228\,
            I => \N__47209\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__47225\,
            I => \N__47209\
        );

    \I__10915\ : CascadeMux
    port map (
            O => \N__47224\,
            I => \N__47206\
        );

    \I__10914\ : CascadeMux
    port map (
            O => \N__47223\,
            I => \N__47203\
        );

    \I__10913\ : Span4Mux_h
    port map (
            O => \N__47220\,
            I => \N__47196\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__47217\,
            I => \N__47196\
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__47214\,
            I => \N__47196\
        );

    \I__10910\ : Span4Mux_v
    port map (
            O => \N__47209\,
            I => \N__47193\
        );

    \I__10909\ : InMux
    port map (
            O => \N__47206\,
            I => \N__47190\
        );

    \I__10908\ : InMux
    port map (
            O => \N__47203\,
            I => \N__47187\
        );

    \I__10907\ : Span4Mux_v
    port map (
            O => \N__47196\,
            I => \N__47184\
        );

    \I__10906\ : Span4Mux_h
    port map (
            O => \N__47193\,
            I => \N__47179\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__47190\,
            I => \N__47179\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__47187\,
            I => \N__47176\
        );

    \I__10903\ : Sp12to4
    port map (
            O => \N__47184\,
            I => \N__47171\
        );

    \I__10902\ : Span4Mux_v
    port map (
            O => \N__47179\,
            I => \N__47166\
        );

    \I__10901\ : Span4Mux_v
    port map (
            O => \N__47176\,
            I => \N__47166\
        );

    \I__10900\ : InMux
    port map (
            O => \N__47175\,
            I => \N__47163\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47160\
        );

    \I__10898\ : Odrv12
    port map (
            O => \N__47171\,
            I => comm_rx_buf_2
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__47166\,
            I => comm_rx_buf_2
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47163\,
            I => comm_rx_buf_2
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__47160\,
            I => comm_rx_buf_2
        );

    \I__10894\ : CascadeMux
    port map (
            O => \N__47151\,
            I => \n30_adj_1520_cascade_\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47148\,
            I => \N__47144\
        );

    \I__10892\ : CascadeMux
    port map (
            O => \N__47147\,
            I => \N__47141\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__47144\,
            I => \N__47138\
        );

    \I__10890\ : InMux
    port map (
            O => \N__47141\,
            I => \N__47135\
        );

    \I__10889\ : Span4Mux_h
    port map (
            O => \N__47138\,
            I => \N__47132\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__47135\,
            I => data_idxvec_2
        );

    \I__10887\ : Odrv4
    port map (
            O => \N__47132\,
            I => data_idxvec_2
        );

    \I__10886\ : InMux
    port map (
            O => \N__47127\,
            I => \N__47124\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__47124\,
            I => \N__47119\
        );

    \I__10884\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47116\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47113\
        );

    \I__10882\ : Span4Mux_h
    port map (
            O => \N__47119\,
            I => \N__47110\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__47116\,
            I => data_cntvec_2
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__47113\,
            I => data_cntvec_2
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__47110\,
            I => data_cntvec_2
        );

    \I__10878\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47100\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__47100\,
            I => n26_adj_1519
        );

    \I__10876\ : InMux
    port map (
            O => \N__47097\,
            I => \N__47093\
        );

    \I__10875\ : InMux
    port map (
            O => \N__47096\,
            I => \N__47089\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__47093\,
            I => \N__47086\
        );

    \I__10873\ : InMux
    port map (
            O => \N__47092\,
            I => \N__47083\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__47089\,
            I => \N__47080\
        );

    \I__10871\ : Span4Mux_v
    port map (
            O => \N__47086\,
            I => \N__47077\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__47083\,
            I => \N__47074\
        );

    \I__10869\ : Span4Mux_h
    port map (
            O => \N__47080\,
            I => \N__47071\
        );

    \I__10868\ : Span4Mux_h
    port map (
            O => \N__47077\,
            I => \N__47068\
        );

    \I__10867\ : Span4Mux_v
    port map (
            O => \N__47074\,
            I => \N__47063\
        );

    \I__10866\ : Span4Mux_h
    port map (
            O => \N__47071\,
            I => \N__47063\
        );

    \I__10865\ : Odrv4
    port map (
            O => \N__47068\,
            I => n14_adj_1585
        );

    \I__10864\ : Odrv4
    port map (
            O => \N__47063\,
            I => n14_adj_1585
        );

    \I__10863\ : InMux
    port map (
            O => \N__47058\,
            I => \N__47055\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__47055\,
            I => \N__47052\
        );

    \I__10861\ : Span4Mux_h
    port map (
            O => \N__47052\,
            I => \N__47049\
        );

    \I__10860\ : Odrv4
    port map (
            O => \N__47049\,
            I => n8
        );

    \I__10859\ : InMux
    port map (
            O => \N__47046\,
            I => \N__47043\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__47043\,
            I => \N__47040\
        );

    \I__10857\ : Span4Mux_v
    port map (
            O => \N__47040\,
            I => \N__47036\
        );

    \I__10856\ : InMux
    port map (
            O => \N__47039\,
            I => \N__47033\
        );

    \I__10855\ : Sp12to4
    port map (
            O => \N__47036\,
            I => \N__47027\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__47033\,
            I => \N__47027\
        );

    \I__10853\ : InMux
    port map (
            O => \N__47032\,
            I => \N__47024\
        );

    \I__10852\ : Span12Mux_h
    port map (
            O => \N__47027\,
            I => \N__47021\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__47024\,
            I => buf_adcdata_iac_14
        );

    \I__10850\ : Odrv12
    port map (
            O => \N__47021\,
            I => buf_adcdata_iac_14
        );

    \I__10849\ : InMux
    port map (
            O => \N__47016\,
            I => \N__47013\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__47013\,
            I => \N__47010\
        );

    \I__10847\ : Odrv4
    port map (
            O => \N__47010\,
            I => n16
        );

    \I__10846\ : InMux
    port map (
            O => \N__47007\,
            I => \N__47004\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__47004\,
            I => \N__47001\
        );

    \I__10844\ : Odrv4
    port map (
            O => \N__47001\,
            I => n21045
        );

    \I__10843\ : InMux
    port map (
            O => \N__46998\,
            I => \N__46994\
        );

    \I__10842\ : CascadeMux
    port map (
            O => \N__46997\,
            I => \N__46990\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46994\,
            I => \N__46987\
        );

    \I__10840\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46982\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46990\,
            I => \N__46982\
        );

    \I__10838\ : Odrv12
    port map (
            O => \N__46987\,
            I => req_data_cnt_7
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__46982\,
            I => req_data_cnt_7
        );

    \I__10836\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46973\
        );

    \I__10835\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46969\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__46973\,
            I => \N__46966\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46972\,
            I => \N__46963\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46969\,
            I => \acadc_skipCount_7\
        );

    \I__10831\ : Odrv4
    port map (
            O => \N__46966\,
            I => \acadc_skipCount_7\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__46963\,
            I => \acadc_skipCount_7\
        );

    \I__10829\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46953\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__46953\,
            I => \N__46949\
        );

    \I__10827\ : CascadeMux
    port map (
            O => \N__46952\,
            I => \N__46946\
        );

    \I__10826\ : Sp12to4
    port map (
            O => \N__46949\,
            I => \N__46942\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46939\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46945\,
            I => \N__46936\
        );

    \I__10823\ : Span12Mux_v
    port map (
            O => \N__46942\,
            I => \N__46933\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__46939\,
            I => \N__46930\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__46936\,
            I => buf_dds1_3
        );

    \I__10820\ : Odrv12
    port map (
            O => \N__46933\,
            I => buf_dds1_3
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__46930\,
            I => buf_dds1_3
        );

    \I__10818\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46920\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__46920\,
            I => \N__46917\
        );

    \I__10816\ : Span4Mux_h
    port map (
            O => \N__46917\,
            I => \N__46912\
        );

    \I__10815\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46909\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46906\
        );

    \I__10813\ : Span4Mux_h
    port map (
            O => \N__46912\,
            I => \N__46903\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46909\,
            I => \N__46900\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__46906\,
            I => buf_dds0_3
        );

    \I__10810\ : Odrv4
    port map (
            O => \N__46903\,
            I => buf_dds0_3
        );

    \I__10809\ : Odrv4
    port map (
            O => \N__46900\,
            I => buf_dds0_3
        );

    \I__10808\ : InMux
    port map (
            O => \N__46893\,
            I => \N__46888\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46885\
        );

    \I__10806\ : CascadeMux
    port map (
            O => \N__46891\,
            I => \N__46882\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46888\,
            I => \N__46879\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__46885\,
            I => \N__46876\
        );

    \I__10803\ : InMux
    port map (
            O => \N__46882\,
            I => \N__46873\
        );

    \I__10802\ : Span4Mux_h
    port map (
            O => \N__46879\,
            I => \N__46868\
        );

    \I__10801\ : Span4Mux_v
    port map (
            O => \N__46876\,
            I => \N__46868\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__46873\,
            I => buf_dds1_2
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__46868\,
            I => buf_dds1_2
        );

    \I__10798\ : InMux
    port map (
            O => \N__46863\,
            I => \N__46860\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__46860\,
            I => \N__46857\
        );

    \I__10796\ : Odrv4
    port map (
            O => \N__46857\,
            I => n16_adj_1517
        );

    \I__10795\ : CascadeMux
    port map (
            O => \N__46854\,
            I => \n26_adj_1512_cascade_\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46848\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__46848\,
            I => \N__46845\
        );

    \I__10792\ : Span4Mux_h
    port map (
            O => \N__46845\,
            I => \N__46842\
        );

    \I__10791\ : Span4Mux_v
    port map (
            O => \N__46842\,
            I => \N__46839\
        );

    \I__10790\ : Span4Mux_h
    port map (
            O => \N__46839\,
            I => \N__46834\
        );

    \I__10789\ : InMux
    port map (
            O => \N__46838\,
            I => \N__46829\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46837\,
            I => \N__46829\
        );

    \I__10787\ : Odrv4
    port map (
            O => \N__46834\,
            I => \acadc_skipCount_4\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__46829\,
            I => \acadc_skipCount_4\
        );

    \I__10785\ : CascadeMux
    port map (
            O => \N__46824\,
            I => \n22351_cascade_\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46821\,
            I => \N__46818\
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__46818\,
            I => \N__46814\
        );

    \I__10782\ : CascadeMux
    port map (
            O => \N__46817\,
            I => \N__46810\
        );

    \I__10781\ : Span4Mux_v
    port map (
            O => \N__46814\,
            I => \N__46807\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46802\
        );

    \I__10779\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46802\
        );

    \I__10778\ : Odrv4
    port map (
            O => \N__46807\,
            I => req_data_cnt_4
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__46802\,
            I => req_data_cnt_4
        );

    \I__10776\ : InMux
    port map (
            O => \N__46797\,
            I => \N__46794\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46794\,
            I => n22234
        );

    \I__10774\ : CascadeMux
    port map (
            O => \N__46791\,
            I => \n22354_cascade_\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46783\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46780\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46786\,
            I => \N__46777\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46783\,
            I => \N__46773\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__46780\,
            I => \N__46769\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__46777\,
            I => \N__46766\
        );

    \I__10767\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46763\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__46773\,
            I => \N__46759\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46756\
        );

    \I__10764\ : Span4Mux_v
    port map (
            O => \N__46769\,
            I => \N__46748\
        );

    \I__10763\ : Span4Mux_h
    port map (
            O => \N__46766\,
            I => \N__46748\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__46763\,
            I => \N__46748\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46762\,
            I => \N__46745\
        );

    \I__10760\ : Span4Mux_v
    port map (
            O => \N__46759\,
            I => \N__46740\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46756\,
            I => \N__46740\
        );

    \I__10758\ : CascadeMux
    port map (
            O => \N__46755\,
            I => \N__46737\
        );

    \I__10757\ : Span4Mux_v
    port map (
            O => \N__46748\,
            I => \N__46734\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__46745\,
            I => \N__46731\
        );

    \I__10755\ : Span4Mux_h
    port map (
            O => \N__46740\,
            I => \N__46727\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46737\,
            I => \N__46724\
        );

    \I__10753\ : Span4Mux_h
    port map (
            O => \N__46734\,
            I => \N__46719\
        );

    \I__10752\ : Span4Mux_h
    port map (
            O => \N__46731\,
            I => \N__46719\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46730\,
            I => \N__46716\
        );

    \I__10750\ : Span4Mux_h
    port map (
            O => \N__46727\,
            I => \N__46712\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__46724\,
            I => \N__46709\
        );

    \I__10748\ : Sp12to4
    port map (
            O => \N__46719\,
            I => \N__46706\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__46716\,
            I => \N__46703\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46700\
        );

    \I__10745\ : Odrv4
    port map (
            O => \N__46712\,
            I => comm_rx_buf_4
        );

    \I__10744\ : Odrv4
    port map (
            O => \N__46709\,
            I => comm_rx_buf_4
        );

    \I__10743\ : Odrv12
    port map (
            O => \N__46706\,
            I => comm_rx_buf_4
        );

    \I__10742\ : Odrv4
    port map (
            O => \N__46703\,
            I => comm_rx_buf_4
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46700\,
            I => comm_rx_buf_4
        );

    \I__10740\ : CascadeMux
    port map (
            O => \N__46689\,
            I => \n30_adj_1513_cascade_\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46686\,
            I => \N__46683\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__46683\,
            I => \N__46680\
        );

    \I__10737\ : Span4Mux_h
    port map (
            O => \N__46680\,
            I => \N__46677\
        );

    \I__10736\ : Odrv4
    port map (
            O => \N__46677\,
            I => n19_adj_1518
        );

    \I__10735\ : CascadeMux
    port map (
            O => \N__46674\,
            I => \N__46671\
        );

    \I__10734\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46668\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__46668\,
            I => \N__46665\
        );

    \I__10732\ : Span12Mux_h
    port map (
            O => \N__46665\,
            I => \N__46661\
        );

    \I__10731\ : CascadeMux
    port map (
            O => \N__46664\,
            I => \N__46658\
        );

    \I__10730\ : Span12Mux_h
    port map (
            O => \N__46661\,
            I => \N__46655\
        );

    \I__10729\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46652\
        );

    \I__10728\ : Odrv12
    port map (
            O => \N__46655\,
            I => \buf_readRTD_2\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__46652\,
            I => \buf_readRTD_2\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46644\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46641\
        );

    \I__10724\ : Span4Mux_v
    port map (
            O => \N__46641\,
            I => \N__46637\
        );

    \I__10723\ : InMux
    port map (
            O => \N__46640\,
            I => \N__46634\
        );

    \I__10722\ : Sp12to4
    port map (
            O => \N__46637\,
            I => \N__46628\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__46634\,
            I => \N__46628\
        );

    \I__10720\ : InMux
    port map (
            O => \N__46633\,
            I => \N__46625\
        );

    \I__10719\ : Span12Mux_h
    port map (
            O => \N__46628\,
            I => \N__46622\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__46625\,
            I => buf_adcdata_iac_10
        );

    \I__10717\ : Odrv12
    port map (
            O => \N__46622\,
            I => buf_adcdata_iac_10
        );

    \I__10716\ : CascadeMux
    port map (
            O => \N__46617\,
            I => \n22207_cascade_\
        );

    \I__10715\ : InMux
    port map (
            O => \N__46614\,
            I => \N__46611\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__46611\,
            I => \N__46608\
        );

    \I__10713\ : Span4Mux_v
    port map (
            O => \N__46608\,
            I => \N__46604\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46607\,
            I => \N__46600\
        );

    \I__10711\ : Span4Mux_h
    port map (
            O => \N__46604\,
            I => \N__46597\
        );

    \I__10710\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46594\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__46600\,
            I => req_data_cnt_2
        );

    \I__10708\ : Odrv4
    port map (
            O => \N__46597\,
            I => req_data_cnt_2
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__46594\,
            I => req_data_cnt_2
        );

    \I__10706\ : CascadeMux
    port map (
            O => \N__46587\,
            I => \n22429_cascade_\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46581\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__46581\,
            I => \N__46576\
        );

    \I__10703\ : CascadeMux
    port map (
            O => \N__46580\,
            I => \N__46573\
        );

    \I__10702\ : InMux
    port map (
            O => \N__46579\,
            I => \N__46570\
        );

    \I__10701\ : Span4Mux_h
    port map (
            O => \N__46576\,
            I => \N__46567\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46573\,
            I => \N__46564\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__46570\,
            I => \acadc_skipCount_2\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__46567\,
            I => \acadc_skipCount_2\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__46564\,
            I => \acadc_skipCount_2\
        );

    \I__10696\ : CascadeMux
    port map (
            O => \N__46557\,
            I => \N__46554\
        );

    \I__10695\ : InMux
    port map (
            O => \N__46554\,
            I => \N__46551\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__46551\,
            I => \N__46548\
        );

    \I__10693\ : Span4Mux_v
    port map (
            O => \N__46548\,
            I => \N__46545\
        );

    \I__10692\ : Span4Mux_h
    port map (
            O => \N__46545\,
            I => \N__46542\
        );

    \I__10691\ : Odrv4
    port map (
            O => \N__46542\,
            I => n21177
        );

    \I__10690\ : CascadeMux
    port map (
            O => \N__46539\,
            I => \n22225_cascade_\
        );

    \I__10689\ : InMux
    port map (
            O => \N__46536\,
            I => \N__46532\
        );

    \I__10688\ : CascadeMux
    port map (
            O => \N__46535\,
            I => \N__46529\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__46532\,
            I => \N__46526\
        );

    \I__10686\ : InMux
    port map (
            O => \N__46529\,
            I => \N__46523\
        );

    \I__10685\ : Span4Mux_h
    port map (
            O => \N__46526\,
            I => \N__46520\
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__46523\,
            I => data_idxvec_6
        );

    \I__10683\ : Odrv4
    port map (
            O => \N__46520\,
            I => data_idxvec_6
        );

    \I__10682\ : InMux
    port map (
            O => \N__46515\,
            I => \N__46512\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__46512\,
            I => \N__46508\
        );

    \I__10680\ : InMux
    port map (
            O => \N__46511\,
            I => \N__46504\
        );

    \I__10679\ : Span4Mux_v
    port map (
            O => \N__46508\,
            I => \N__46501\
        );

    \I__10678\ : InMux
    port map (
            O => \N__46507\,
            I => \N__46498\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__46504\,
            I => \N__46495\
        );

    \I__10676\ : Span4Mux_h
    port map (
            O => \N__46501\,
            I => \N__46492\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__46498\,
            I => data_cntvec_6
        );

    \I__10674\ : Odrv4
    port map (
            O => \N__46495\,
            I => data_cntvec_6
        );

    \I__10673\ : Odrv4
    port map (
            O => \N__46492\,
            I => data_cntvec_6
        );

    \I__10672\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46482\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__46482\,
            I => \N__46479\
        );

    \I__10670\ : Span12Mux_h
    port map (
            O => \N__46479\,
            I => \N__46476\
        );

    \I__10669\ : Odrv12
    port map (
            O => \N__46476\,
            I => buf_data_iac_14
        );

    \I__10668\ : CascadeMux
    port map (
            O => \N__46473\,
            I => \n26_adj_1507_cascade_\
        );

    \I__10667\ : InMux
    port map (
            O => \N__46470\,
            I => \N__46467\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__46467\,
            I => n21178
        );

    \I__10665\ : CascadeMux
    port map (
            O => \N__46464\,
            I => \N__46458\
        );

    \I__10664\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46455\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46452\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46449\
        );

    \I__10661\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46443\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__46455\,
            I => \N__46436\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__46452\,
            I => \N__46436\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__46449\,
            I => \N__46436\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__46448\,
            I => \N__46433\
        );

    \I__10656\ : InMux
    port map (
            O => \N__46447\,
            I => \N__46430\
        );

    \I__10655\ : InMux
    port map (
            O => \N__46446\,
            I => \N__46427\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__46443\,
            I => \N__46424\
        );

    \I__10653\ : Span4Mux_v
    port map (
            O => \N__46436\,
            I => \N__46421\
        );

    \I__10652\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46418\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__46430\,
            I => \N__46413\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__46427\,
            I => \N__46413\
        );

    \I__10649\ : Span4Mux_v
    port map (
            O => \N__46424\,
            I => \N__46406\
        );

    \I__10648\ : Span4Mux_h
    port map (
            O => \N__46421\,
            I => \N__46406\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__46418\,
            I => \N__46406\
        );

    \I__10646\ : Span4Mux_v
    port map (
            O => \N__46413\,
            I => \N__46401\
        );

    \I__10645\ : Span4Mux_v
    port map (
            O => \N__46406\,
            I => \N__46398\
        );

    \I__10644\ : InMux
    port map (
            O => \N__46405\,
            I => \N__46395\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46404\,
            I => \N__46392\
        );

    \I__10642\ : Odrv4
    port map (
            O => \N__46401\,
            I => comm_rx_buf_6
        );

    \I__10641\ : Odrv4
    port map (
            O => \N__46398\,
            I => comm_rx_buf_6
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__46395\,
            I => comm_rx_buf_6
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46392\,
            I => comm_rx_buf_6
        );

    \I__10638\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46380\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46380\,
            I => n22228
        );

    \I__10636\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46374\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__46374\,
            I => \N__46371\
        );

    \I__10634\ : Span4Mux_h
    port map (
            O => \N__46371\,
            I => \N__46368\
        );

    \I__10633\ : Span4Mux_h
    port map (
            O => \N__46368\,
            I => \N__46365\
        );

    \I__10632\ : Span4Mux_v
    port map (
            O => \N__46365\,
            I => \N__46361\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46364\,
            I => \N__46358\
        );

    \I__10630\ : Odrv4
    port map (
            O => \N__46361\,
            I => buf_adcdata_vdc_14
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__46358\,
            I => buf_adcdata_vdc_14
        );

    \I__10628\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46350\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46350\,
            I => \N__46346\
        );

    \I__10626\ : InMux
    port map (
            O => \N__46349\,
            I => \N__46343\
        );

    \I__10625\ : Span12Mux_v
    port map (
            O => \N__46346\,
            I => \N__46339\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__46343\,
            I => \N__46336\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46342\,
            I => \N__46333\
        );

    \I__10622\ : Span12Mux_h
    port map (
            O => \N__46339\,
            I => \N__46330\
        );

    \I__10621\ : Span12Mux_s10_h
    port map (
            O => \N__46336\,
            I => \N__46327\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__46333\,
            I => buf_adcdata_vac_14
        );

    \I__10619\ : Odrv12
    port map (
            O => \N__46330\,
            I => buf_adcdata_vac_14
        );

    \I__10618\ : Odrv12
    port map (
            O => \N__46327\,
            I => buf_adcdata_vac_14
        );

    \I__10617\ : CascadeMux
    port map (
            O => \N__46320\,
            I => \n19_cascade_\
        );

    \I__10616\ : InMux
    port map (
            O => \N__46317\,
            I => \N__46314\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__46314\,
            I => \N__46311\
        );

    \I__10614\ : Span4Mux_v
    port map (
            O => \N__46311\,
            I => \N__46308\
        );

    \I__10613\ : Span4Mux_h
    port map (
            O => \N__46308\,
            I => \N__46305\
        );

    \I__10612\ : Span4Mux_h
    port map (
            O => \N__46305\,
            I => \N__46301\
        );

    \I__10611\ : CascadeMux
    port map (
            O => \N__46304\,
            I => \N__46298\
        );

    \I__10610\ : Span4Mux_h
    port map (
            O => \N__46301\,
            I => \N__46295\
        );

    \I__10609\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46292\
        );

    \I__10608\ : Odrv4
    port map (
            O => \N__46295\,
            I => \buf_readRTD_6\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__46292\,
            I => \buf_readRTD_6\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46284\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46284\,
            I => n21046
        );

    \I__10604\ : InMux
    port map (
            O => \N__46281\,
            I => \N__46278\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__46278\,
            I => \N__46275\
        );

    \I__10602\ : Sp12to4
    port map (
            O => \N__46275\,
            I => \N__46272\
        );

    \I__10601\ : Odrv12
    port map (
            O => \N__46272\,
            I => n16_adj_1510
        );

    \I__10600\ : CascadeMux
    port map (
            O => \N__46269\,
            I => \N__46265\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46268\,
            I => \N__46262\
        );

    \I__10598\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46259\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__46262\,
            I => \N__46256\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__46259\,
            I => \N__46252\
        );

    \I__10595\ : Span12Mux_v
    port map (
            O => \N__46256\,
            I => \N__46249\
        );

    \I__10594\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46246\
        );

    \I__10593\ : Span4Mux_h
    port map (
            O => \N__46252\,
            I => \N__46243\
        );

    \I__10592\ : Span12Mux_h
    port map (
            O => \N__46249\,
            I => \N__46240\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__46246\,
            I => \N__46235\
        );

    \I__10590\ : Span4Mux_h
    port map (
            O => \N__46243\,
            I => \N__46235\
        );

    \I__10589\ : Odrv12
    port map (
            O => \N__46240\,
            I => buf_adcdata_iac_12
        );

    \I__10588\ : Odrv4
    port map (
            O => \N__46235\,
            I => buf_adcdata_iac_12
        );

    \I__10587\ : InMux
    port map (
            O => \N__46230\,
            I => \N__46227\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__46227\,
            I => \N__46224\
        );

    \I__10585\ : Sp12to4
    port map (
            O => \N__46224\,
            I => \N__46221\
        );

    \I__10584\ : Odrv12
    port map (
            O => \N__46221\,
            I => n22231
        );

    \I__10583\ : InMux
    port map (
            O => \N__46218\,
            I => \N__46214\
        );

    \I__10582\ : CascadeMux
    port map (
            O => \N__46217\,
            I => \N__46211\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__46214\,
            I => \N__46208\
        );

    \I__10580\ : InMux
    port map (
            O => \N__46211\,
            I => \N__46205\
        );

    \I__10579\ : Span4Mux_h
    port map (
            O => \N__46208\,
            I => \N__46202\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__46205\,
            I => data_idxvec_4
        );

    \I__10577\ : Odrv4
    port map (
            O => \N__46202\,
            I => data_idxvec_4
        );

    \I__10576\ : InMux
    port map (
            O => \N__46197\,
            I => \N__46194\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__46194\,
            I => \N__46189\
        );

    \I__10574\ : InMux
    port map (
            O => \N__46193\,
            I => \N__46186\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46183\
        );

    \I__10572\ : Span4Mux_v
    port map (
            O => \N__46189\,
            I => \N__46180\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__46186\,
            I => data_cntvec_4
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__46183\,
            I => data_cntvec_4
        );

    \I__10569\ : Odrv4
    port map (
            O => \N__46180\,
            I => data_cntvec_4
        );

    \I__10568\ : CEMux
    port map (
            O => \N__46173\,
            I => \N__46170\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__46170\,
            I => \N__46161\
        );

    \I__10566\ : CEMux
    port map (
            O => \N__46169\,
            I => \N__46158\
        );

    \I__10565\ : CEMux
    port map (
            O => \N__46168\,
            I => \N__46155\
        );

    \I__10564\ : CEMux
    port map (
            O => \N__46167\,
            I => \N__46152\
        );

    \I__10563\ : CEMux
    port map (
            O => \N__46166\,
            I => \N__46149\
        );

    \I__10562\ : CEMux
    port map (
            O => \N__46165\,
            I => \N__46146\
        );

    \I__10561\ : CEMux
    port map (
            O => \N__46164\,
            I => \N__46143\
        );

    \I__10560\ : Span4Mux_v
    port map (
            O => \N__46161\,
            I => \N__46138\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__46158\,
            I => \N__46138\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__46155\,
            I => \N__46135\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__46152\,
            I => \N__46132\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46127\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46146\,
            I => \N__46127\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__46143\,
            I => \N__46124\
        );

    \I__10553\ : Span4Mux_v
    port map (
            O => \N__46138\,
            I => \N__46120\
        );

    \I__10552\ : Span4Mux_h
    port map (
            O => \N__46135\,
            I => \N__46117\
        );

    \I__10551\ : Span4Mux_h
    port map (
            O => \N__46132\,
            I => \N__46114\
        );

    \I__10550\ : Span4Mux_v
    port map (
            O => \N__46127\,
            I => \N__46109\
        );

    \I__10549\ : Span4Mux_h
    port map (
            O => \N__46124\,
            I => \N__46109\
        );

    \I__10548\ : InMux
    port map (
            O => \N__46123\,
            I => \N__46106\
        );

    \I__10547\ : Odrv4
    port map (
            O => \N__46120\,
            I => n11961
        );

    \I__10546\ : Odrv4
    port map (
            O => \N__46117\,
            I => n11961
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__46114\,
            I => n11961
        );

    \I__10544\ : Odrv4
    port map (
            O => \N__46109\,
            I => n11961
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__46106\,
            I => n11961
        );

    \I__10542\ : CascadeMux
    port map (
            O => \N__46095\,
            I => \n18993_cascade_\
        );

    \I__10541\ : InMux
    port map (
            O => \N__46092\,
            I => \N__46089\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__46089\,
            I => n12_adj_1605
        );

    \I__10539\ : CascadeMux
    port map (
            O => \N__46086\,
            I => \n11991_cascade_\
        );

    \I__10538\ : InMux
    port map (
            O => \N__46083\,
            I => \N__46075\
        );

    \I__10537\ : CascadeMux
    port map (
            O => \N__46082\,
            I => \N__46072\
        );

    \I__10536\ : InMux
    port map (
            O => \N__46081\,
            I => \N__46067\
        );

    \I__10535\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46064\
        );

    \I__10534\ : InMux
    port map (
            O => \N__46079\,
            I => \N__46061\
        );

    \I__10533\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46058\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__46075\,
            I => \N__46055\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46072\,
            I => \N__46050\
        );

    \I__10530\ : InMux
    port map (
            O => \N__46071\,
            I => \N__46050\
        );

    \I__10529\ : InMux
    port map (
            O => \N__46070\,
            I => \N__46047\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__46067\,
            I => \N__46040\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__46064\,
            I => \N__46040\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__46061\,
            I => \N__46040\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__46058\,
            I => \N__46037\
        );

    \I__10524\ : Span4Mux_h
    port map (
            O => \N__46055\,
            I => \N__46032\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__46050\,
            I => \N__46032\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__46047\,
            I => \N__46025\
        );

    \I__10521\ : Span4Mux_v
    port map (
            O => \N__46040\,
            I => \N__46025\
        );

    \I__10520\ : Span4Mux_h
    port map (
            O => \N__46037\,
            I => \N__46025\
        );

    \I__10519\ : Span4Mux_h
    port map (
            O => \N__46032\,
            I => \N__46022\
        );

    \I__10518\ : Span4Mux_h
    port map (
            O => \N__46025\,
            I => \N__46019\
        );

    \I__10517\ : Odrv4
    port map (
            O => \N__46022\,
            I => n14506
        );

    \I__10516\ : Odrv4
    port map (
            O => \N__46019\,
            I => n14506
        );

    \I__10515\ : InMux
    port map (
            O => \N__46014\,
            I => \N__46009\
        );

    \I__10514\ : InMux
    port map (
            O => \N__46013\,
            I => \N__46005\
        );

    \I__10513\ : InMux
    port map (
            O => \N__46012\,
            I => \N__46002\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__46009\,
            I => \N__45995\
        );

    \I__10511\ : InMux
    port map (
            O => \N__46008\,
            I => \N__45992\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__46005\,
            I => \N__45987\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__46002\,
            I => \N__45987\
        );

    \I__10508\ : InMux
    port map (
            O => \N__46001\,
            I => \N__45984\
        );

    \I__10507\ : InMux
    port map (
            O => \N__46000\,
            I => \N__45979\
        );

    \I__10506\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45979\
        );

    \I__10505\ : InMux
    port map (
            O => \N__45998\,
            I => \N__45976\
        );

    \I__10504\ : Span4Mux_h
    port map (
            O => \N__45995\,
            I => \N__45973\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45992\,
            I => \N__45970\
        );

    \I__10502\ : Span4Mux_v
    port map (
            O => \N__45987\,
            I => \N__45961\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__45984\,
            I => \N__45961\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__45979\,
            I => \N__45961\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__45976\,
            I => \N__45961\
        );

    \I__10498\ : Odrv4
    port map (
            O => \N__45973\,
            I => n11896
        );

    \I__10497\ : Odrv12
    port map (
            O => \N__45970\,
            I => n11896
        );

    \I__10496\ : Odrv4
    port map (
            O => \N__45961\,
            I => n11896
        );

    \I__10495\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45949\
        );

    \I__10494\ : InMux
    port map (
            O => \N__45953\,
            I => \N__45944\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45952\,
            I => \N__45944\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__45949\,
            I => \N__45939\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__45944\,
            I => \N__45939\
        );

    \I__10490\ : Span12Mux_v
    port map (
            O => \N__45939\,
            I => \N__45936\
        );

    \I__10489\ : Odrv12
    port map (
            O => \N__45936\,
            I => n10697
        );

    \I__10488\ : InMux
    port map (
            O => \N__45933\,
            I => \N__45930\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__45930\,
            I => n18993
        );

    \I__10486\ : InMux
    port map (
            O => \N__45927\,
            I => \N__45924\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45924\,
            I => \N__45921\
        );

    \I__10484\ : Span4Mux_h
    port map (
            O => \N__45921\,
            I => \N__45917\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__45920\,
            I => \N__45911\
        );

    \I__10482\ : Span4Mux_h
    port map (
            O => \N__45917\,
            I => \N__45907\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45916\,
            I => \N__45904\
        );

    \I__10480\ : InMux
    port map (
            O => \N__45915\,
            I => \N__45899\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45914\,
            I => \N__45899\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45894\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45910\,
            I => \N__45894\
        );

    \I__10476\ : Odrv4
    port map (
            O => \N__45907\,
            I => n20843
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__45904\,
            I => n20843
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45899\,
            I => n20843
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45894\,
            I => n20843
        );

    \I__10472\ : CascadeMux
    port map (
            O => \N__45885\,
            I => \n12_adj_1635_cascade_\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45873\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45881\,
            I => \N__45870\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45880\,
            I => \N__45865\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45865\
        );

    \I__10467\ : CascadeMux
    port map (
            O => \N__45878\,
            I => \N__45862\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45877\,
            I => \N__45856\
        );

    \I__10465\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45856\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__45873\,
            I => \N__45853\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__45870\,
            I => \N__45850\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__45865\,
            I => \N__45847\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45862\,
            I => \N__45843\
        );

    \I__10460\ : InMux
    port map (
            O => \N__45861\,
            I => \N__45840\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__45856\,
            I => \N__45837\
        );

    \I__10458\ : Span4Mux_v
    port map (
            O => \N__45853\,
            I => \N__45834\
        );

    \I__10457\ : Span4Mux_h
    port map (
            O => \N__45850\,
            I => \N__45829\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__45847\,
            I => \N__45829\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45846\,
            I => \N__45826\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__45843\,
            I => \N__45819\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__45840\,
            I => \N__45819\
        );

    \I__10452\ : Span4Mux_h
    port map (
            O => \N__45837\,
            I => \N__45819\
        );

    \I__10451\ : Odrv4
    port map (
            O => \N__45834\,
            I => n20917
        );

    \I__10450\ : Odrv4
    port map (
            O => \N__45829\,
            I => n20917
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45826\,
            I => n20917
        );

    \I__10448\ : Odrv4
    port map (
            O => \N__45819\,
            I => n20917
        );

    \I__10447\ : CEMux
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45807\,
            I => \N__45803\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45806\,
            I => \N__45800\
        );

    \I__10444\ : Odrv4
    port map (
            O => \N__45803\,
            I => n12178
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__45800\,
            I => n12178
        );

    \I__10442\ : InMux
    port map (
            O => \N__45795\,
            I => \N__45788\
        );

    \I__10441\ : CascadeMux
    port map (
            O => \N__45794\,
            I => \N__45784\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45793\,
            I => \N__45781\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45792\,
            I => \N__45778\
        );

    \I__10438\ : CascadeMux
    port map (
            O => \N__45791\,
            I => \N__45775\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__45788\,
            I => \N__45772\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45769\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45784\,
            I => \N__45765\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__45781\,
            I => \N__45760\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__45778\,
            I => \N__45760\
        );

    \I__10432\ : InMux
    port map (
            O => \N__45775\,
            I => \N__45757\
        );

    \I__10431\ : Span4Mux_v
    port map (
            O => \N__45772\,
            I => \N__45754\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45769\,
            I => \N__45751\
        );

    \I__10429\ : InMux
    port map (
            O => \N__45768\,
            I => \N__45748\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45745\
        );

    \I__10427\ : Span4Mux_v
    port map (
            O => \N__45760\,
            I => \N__45740\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45757\,
            I => \N__45740\
        );

    \I__10425\ : Span4Mux_h
    port map (
            O => \N__45754\,
            I => \N__45737\
        );

    \I__10424\ : Span4Mux_v
    port map (
            O => \N__45751\,
            I => \N__45732\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__45748\,
            I => \N__45732\
        );

    \I__10422\ : Span4Mux_v
    port map (
            O => \N__45745\,
            I => \N__45729\
        );

    \I__10421\ : Span4Mux_h
    port map (
            O => \N__45740\,
            I => \N__45726\
        );

    \I__10420\ : Sp12to4
    port map (
            O => \N__45737\,
            I => \N__45721\
        );

    \I__10419\ : Span4Mux_h
    port map (
            O => \N__45732\,
            I => \N__45716\
        );

    \I__10418\ : Span4Mux_h
    port map (
            O => \N__45729\,
            I => \N__45716\
        );

    \I__10417\ : Span4Mux_h
    port map (
            O => \N__45726\,
            I => \N__45713\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45725\,
            I => \N__45710\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45707\
        );

    \I__10414\ : Odrv12
    port map (
            O => \N__45721\,
            I => comm_rx_buf_1
        );

    \I__10413\ : Odrv4
    port map (
            O => \N__45716\,
            I => comm_rx_buf_1
        );

    \I__10412\ : Odrv4
    port map (
            O => \N__45713\,
            I => comm_rx_buf_1
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__45710\,
            I => comm_rx_buf_1
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__45707\,
            I => comm_rx_buf_1
        );

    \I__10409\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__45693\,
            I => \N__45690\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__45690\,
            I => \N__45687\
        );

    \I__10406\ : Odrv4
    port map (
            O => \N__45687\,
            I => buf_data_vac_17
        );

    \I__10405\ : CascadeMux
    port map (
            O => \N__45684\,
            I => \N__45681\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45681\,
            I => \N__45678\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45675\
        );

    \I__10402\ : Span4Mux_h
    port map (
            O => \N__45675\,
            I => \N__45672\
        );

    \I__10401\ : Span4Mux_h
    port map (
            O => \N__45672\,
            I => \N__45669\
        );

    \I__10400\ : Odrv4
    port map (
            O => \N__45669\,
            I => comm_buf_3_1
        );

    \I__10399\ : InMux
    port map (
            O => \N__45666\,
            I => \N__45663\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45663\,
            I => \N__45660\
        );

    \I__10397\ : Odrv12
    port map (
            O => \N__45660\,
            I => n20878
        );

    \I__10396\ : CascadeMux
    port map (
            O => \N__45657\,
            I => \n21352_cascade_\
        );

    \I__10395\ : CascadeMux
    port map (
            O => \N__45654\,
            I => \n12_cascade_\
        );

    \I__10394\ : CEMux
    port map (
            O => \N__45651\,
            I => \N__45648\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__45648\,
            I => n12136
        );

    \I__10392\ : CascadeMux
    port map (
            O => \N__45645\,
            I => \n12136_cascade_\
        );

    \I__10391\ : SRMux
    port map (
            O => \N__45642\,
            I => \N__45639\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45639\,
            I => n14771
        );

    \I__10389\ : InMux
    port map (
            O => \N__45636\,
            I => \N__45633\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__45633\,
            I => \N__45628\
        );

    \I__10387\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45623\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45631\,
            I => \N__45623\
        );

    \I__10385\ : Span4Mux_v
    port map (
            O => \N__45628\,
            I => \N__45620\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__45623\,
            I => \N__45617\
        );

    \I__10383\ : Sp12to4
    port map (
            O => \N__45620\,
            I => \N__45614\
        );

    \I__10382\ : Span4Mux_v
    port map (
            O => \N__45617\,
            I => \N__45611\
        );

    \I__10381\ : Odrv12
    port map (
            O => \N__45614\,
            I => n19783
        );

    \I__10380\ : Odrv4
    port map (
            O => \N__45611\,
            I => n19783
        );

    \I__10379\ : CascadeMux
    port map (
            O => \N__45606\,
            I => \n18991_cascade_\
        );

    \I__10378\ : CascadeMux
    port map (
            O => \N__45603\,
            I => \n4_adj_1545_cascade_\
        );

    \I__10377\ : InMux
    port map (
            O => \N__45600\,
            I => \N__45597\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45597\,
            I => \N__45594\
        );

    \I__10375\ : Span4Mux_h
    port map (
            O => \N__45594\,
            I => \N__45590\
        );

    \I__10374\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45587\
        );

    \I__10373\ : Span4Mux_h
    port map (
            O => \N__45590\,
            I => \N__45584\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45587\,
            I => comm_buf_6_6
        );

    \I__10371\ : Odrv4
    port map (
            O => \N__45584\,
            I => comm_buf_6_6
        );

    \I__10370\ : InMux
    port map (
            O => \N__45579\,
            I => \N__45576\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__45576\,
            I => n4_adj_1590
        );

    \I__10368\ : CascadeMux
    port map (
            O => \N__45573\,
            I => \n21539_cascade_\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45567\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__45567\,
            I => n22339
        );

    \I__10365\ : InMux
    port map (
            O => \N__45564\,
            I => \N__45561\
        );

    \I__10364\ : LocalMux
    port map (
            O => \N__45561\,
            I => \N__45558\
        );

    \I__10363\ : Span4Mux_h
    port map (
            O => \N__45558\,
            I => \N__45555\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__45555\,
            I => buf_data_vac_16
        );

    \I__10361\ : InMux
    port map (
            O => \N__45552\,
            I => \N__45549\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__45549\,
            I => comm_buf_3_0
        );

    \I__10359\ : InMux
    port map (
            O => \N__45546\,
            I => \N__45543\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__45543\,
            I => \N__45540\
        );

    \I__10357\ : Span4Mux_v
    port map (
            O => \N__45540\,
            I => \N__45537\
        );

    \I__10356\ : Span4Mux_h
    port map (
            O => \N__45537\,
            I => \N__45534\
        );

    \I__10355\ : Odrv4
    port map (
            O => \N__45534\,
            I => buf_data_vac_20
        );

    \I__10354\ : InMux
    port map (
            O => \N__45531\,
            I => \N__45528\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__45528\,
            I => \N__45525\
        );

    \I__10352\ : Span4Mux_v
    port map (
            O => \N__45525\,
            I => \N__45522\
        );

    \I__10351\ : Odrv4
    port map (
            O => \N__45522\,
            I => comm_buf_3_4
        );

    \I__10350\ : InMux
    port map (
            O => \N__45519\,
            I => \N__45516\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__45516\,
            I => \N__45513\
        );

    \I__10348\ : Span4Mux_v
    port map (
            O => \N__45513\,
            I => \N__45510\
        );

    \I__10347\ : Span4Mux_v
    port map (
            O => \N__45510\,
            I => \N__45507\
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__45507\,
            I => buf_data_vac_23
        );

    \I__10345\ : CascadeMux
    port map (
            O => \N__45504\,
            I => \N__45501\
        );

    \I__10344\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45498\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__45498\,
            I => \N__45495\
        );

    \I__10342\ : Span12Mux_h
    port map (
            O => \N__45495\,
            I => \N__45492\
        );

    \I__10341\ : Odrv12
    port map (
            O => \N__45492\,
            I => comm_buf_3_7
        );

    \I__10340\ : InMux
    port map (
            O => \N__45489\,
            I => \N__45486\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__45486\,
            I => \N__45483\
        );

    \I__10338\ : Span4Mux_h
    port map (
            O => \N__45483\,
            I => \N__45480\
        );

    \I__10337\ : Span4Mux_v
    port map (
            O => \N__45480\,
            I => \N__45477\
        );

    \I__10336\ : Odrv4
    port map (
            O => \N__45477\,
            I => buf_data_vac_22
        );

    \I__10335\ : InMux
    port map (
            O => \N__45474\,
            I => \N__45471\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__45471\,
            I => \N__45468\
        );

    \I__10333\ : Odrv4
    port map (
            O => \N__45468\,
            I => comm_buf_3_6
        );

    \I__10332\ : InMux
    port map (
            O => \N__45465\,
            I => \N__45462\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45462\,
            I => \N__45459\
        );

    \I__10330\ : Span4Mux_h
    port map (
            O => \N__45459\,
            I => \N__45456\
        );

    \I__10329\ : Span4Mux_v
    port map (
            O => \N__45456\,
            I => \N__45453\
        );

    \I__10328\ : Odrv4
    port map (
            O => \N__45453\,
            I => buf_data_vac_21
        );

    \I__10327\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45447\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__45447\,
            I => comm_buf_3_5
        );

    \I__10325\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45441\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__45441\,
            I => \N__45438\
        );

    \I__10323\ : Odrv4
    port map (
            O => \N__45438\,
            I => buf_data_vac_19
        );

    \I__10322\ : CascadeMux
    port map (
            O => \N__45435\,
            I => \N__45432\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45432\,
            I => \N__45429\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__45429\,
            I => \N__45426\
        );

    \I__10319\ : Span4Mux_h
    port map (
            O => \N__45426\,
            I => \N__45423\
        );

    \I__10318\ : Odrv4
    port map (
            O => \N__45423\,
            I => comm_buf_3_3
        );

    \I__10317\ : InMux
    port map (
            O => \N__45420\,
            I => \N__45417\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__45417\,
            I => \N__45414\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__45414\,
            I => \N__45411\
        );

    \I__10314\ : Odrv4
    port map (
            O => \N__45411\,
            I => buf_data_vac_18
        );

    \I__10313\ : CascadeMux
    port map (
            O => \N__45408\,
            I => \N__45405\
        );

    \I__10312\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45402\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45402\,
            I => \N__45399\
        );

    \I__10310\ : Odrv12
    port map (
            O => \N__45399\,
            I => comm_buf_3_2
        );

    \I__10309\ : CascadeMux
    port map (
            O => \N__45396\,
            I => \ADC_VDC.genclk.n21446_cascade_\
        );

    \I__10308\ : InMux
    port map (
            O => \N__45393\,
            I => \N__45390\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__45390\,
            I => \ADC_VDC.genclk.n26\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45387\,
            I => \N__45384\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__45384\,
            I => \ADC_VDC.genclk.n27\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45378\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__45378\,
            I => \ADC_VDC.genclk.n28_adj_1397\
        );

    \I__10302\ : SRMux
    port map (
            O => \N__45375\,
            I => \N__45372\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__45372\,
            I => \N__45369\
        );

    \I__10300\ : Span4Mux_h
    port map (
            O => \N__45369\,
            I => \N__45366\
        );

    \I__10299\ : Odrv4
    port map (
            O => \N__45366\,
            I => \comm_spi.data_tx_7__N_767\
        );

    \I__10298\ : CascadeMux
    port map (
            O => \N__45363\,
            I => \N__45359\
        );

    \I__10297\ : CascadeMux
    port map (
            O => \N__45362\,
            I => \N__45354\
        );

    \I__10296\ : InMux
    port map (
            O => \N__45359\,
            I => \N__45350\
        );

    \I__10295\ : CascadeMux
    port map (
            O => \N__45358\,
            I => \N__45347\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45357\,
            I => \N__45344\
        );

    \I__10293\ : InMux
    port map (
            O => \N__45354\,
            I => \N__45341\
        );

    \I__10292\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45335\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__45350\,
            I => \N__45332\
        );

    \I__10290\ : InMux
    port map (
            O => \N__45347\,
            I => \N__45329\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45344\,
            I => \N__45324\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__45341\,
            I => \N__45324\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45321\
        );

    \I__10286\ : CascadeMux
    port map (
            O => \N__45339\,
            I => \N__45318\
        );

    \I__10285\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45315\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__45335\,
            I => \N__45308\
        );

    \I__10283\ : Span4Mux_h
    port map (
            O => \N__45332\,
            I => \N__45308\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__45329\,
            I => \N__45308\
        );

    \I__10281\ : Span4Mux_v
    port map (
            O => \N__45324\,
            I => \N__45303\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__45321\,
            I => \N__45303\
        );

    \I__10279\ : InMux
    port map (
            O => \N__45318\,
            I => \N__45300\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45315\,
            I => \N__45297\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__45308\,
            I => \N__45294\
        );

    \I__10276\ : Span4Mux_h
    port map (
            O => \N__45303\,
            I => \N__45291\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__45300\,
            I => \N__45288\
        );

    \I__10274\ : Span4Mux_h
    port map (
            O => \N__45297\,
            I => \N__45285\
        );

    \I__10273\ : Span4Mux_h
    port map (
            O => \N__45294\,
            I => \N__45280\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__45291\,
            I => \N__45280\
        );

    \I__10271\ : Odrv12
    port map (
            O => \N__45288\,
            I => comm_buf_0_6
        );

    \I__10270\ : Odrv4
    port map (
            O => \N__45285\,
            I => comm_buf_0_6
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__45280\,
            I => comm_buf_0_6
        );

    \I__10268\ : CascadeMux
    port map (
            O => \N__45273\,
            I => \n1_adj_1588_cascade_\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45270\,
            I => \N__45267\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__45267\,
            I => \N__45264\
        );

    \I__10265\ : Span4Mux_h
    port map (
            O => \N__45264\,
            I => \N__45261\
        );

    \I__10264\ : Span4Mux_v
    port map (
            O => \N__45261\,
            I => \N__45256\
        );

    \I__10263\ : InMux
    port map (
            O => \N__45260\,
            I => \N__45253\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45259\,
            I => \N__45250\
        );

    \I__10261\ : Odrv4
    port map (
            O => \N__45256\,
            I => comm_tx_buf_6
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__45253\,
            I => comm_tx_buf_6
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__45250\,
            I => comm_tx_buf_6
        );

    \I__10258\ : CEMux
    port map (
            O => \N__45243\,
            I => \N__45240\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__45240\,
            I => \N__45237\
        );

    \I__10256\ : Span4Mux_v
    port map (
            O => \N__45237\,
            I => \N__45230\
        );

    \I__10255\ : CEMux
    port map (
            O => \N__45236\,
            I => \N__45227\
        );

    \I__10254\ : CEMux
    port map (
            O => \N__45235\,
            I => \N__45223\
        );

    \I__10253\ : CEMux
    port map (
            O => \N__45234\,
            I => \N__45220\
        );

    \I__10252\ : CEMux
    port map (
            O => \N__45233\,
            I => \N__45217\
        );

    \I__10251\ : Span4Mux_v
    port map (
            O => \N__45230\,
            I => \N__45212\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__45227\,
            I => \N__45212\
        );

    \I__10249\ : CEMux
    port map (
            O => \N__45226\,
            I => \N__45209\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__45223\,
            I => \N__45206\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__45220\,
            I => \N__45203\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__45217\,
            I => \N__45200\
        );

    \I__10245\ : Span4Mux_v
    port map (
            O => \N__45212\,
            I => \N__45197\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__45209\,
            I => \N__45194\
        );

    \I__10243\ : Span4Mux_v
    port map (
            O => \N__45206\,
            I => \N__45187\
        );

    \I__10242\ : Span4Mux_v
    port map (
            O => \N__45203\,
            I => \N__45187\
        );

    \I__10241\ : Span4Mux_v
    port map (
            O => \N__45200\,
            I => \N__45187\
        );

    \I__10240\ : Span4Mux_h
    port map (
            O => \N__45197\,
            I => \N__45184\
        );

    \I__10239\ : Odrv4
    port map (
            O => \N__45194\,
            I => n12336
        );

    \I__10238\ : Odrv4
    port map (
            O => \N__45187\,
            I => n12336
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__45184\,
            I => n12336
        );

    \I__10236\ : SRMux
    port map (
            O => \N__45177\,
            I => \N__45174\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45174\,
            I => \N__45168\
        );

    \I__10234\ : SRMux
    port map (
            O => \N__45173\,
            I => \N__45165\
        );

    \I__10233\ : SRMux
    port map (
            O => \N__45172\,
            I => \N__45161\
        );

    \I__10232\ : SRMux
    port map (
            O => \N__45171\,
            I => \N__45158\
        );

    \I__10231\ : Span4Mux_h
    port map (
            O => \N__45168\,
            I => \N__45152\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__45165\,
            I => \N__45152\
        );

    \I__10229\ : SRMux
    port map (
            O => \N__45164\,
            I => \N__45149\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__45161\,
            I => \N__45146\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__45158\,
            I => \N__45143\
        );

    \I__10226\ : SRMux
    port map (
            O => \N__45157\,
            I => \N__45140\
        );

    \I__10225\ : Span4Mux_v
    port map (
            O => \N__45152\,
            I => \N__45135\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__45149\,
            I => \N__45135\
        );

    \I__10223\ : Span4Mux_h
    port map (
            O => \N__45146\,
            I => \N__45132\
        );

    \I__10222\ : Span4Mux_h
    port map (
            O => \N__45143\,
            I => \N__45129\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__45140\,
            I => \N__45126\
        );

    \I__10220\ : Span4Mux_h
    port map (
            O => \N__45135\,
            I => \N__45123\
        );

    \I__10219\ : Odrv4
    port map (
            O => \N__45132\,
            I => n14799
        );

    \I__10218\ : Odrv4
    port map (
            O => \N__45129\,
            I => n14799
        );

    \I__10217\ : Odrv4
    port map (
            O => \N__45126\,
            I => n14799
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__45123\,
            I => n14799
        );

    \I__10215\ : InMux
    port map (
            O => \N__45114\,
            I => \N__45111\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__45111\,
            I => \N__45108\
        );

    \I__10213\ : Odrv12
    port map (
            O => \N__45108\,
            I => comm_buf_2_6
        );

    \I__10212\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45102\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__45102\,
            I => n2_adj_1589
        );

    \I__10210\ : InMux
    port map (
            O => \N__45099\,
            I => \N__45096\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__45096\,
            I => n8_adj_1571
        );

    \I__10208\ : InMux
    port map (
            O => \N__45093\,
            I => \N__45089\
        );

    \I__10207\ : InMux
    port map (
            O => \N__45092\,
            I => \N__45086\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__45089\,
            I => \N__45081\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__45086\,
            I => \N__45081\
        );

    \I__10204\ : Span4Mux_h
    port map (
            O => \N__45081\,
            I => \N__45078\
        );

    \I__10203\ : Odrv4
    port map (
            O => \N__45078\,
            I => n7_adj_1570
        );

    \I__10202\ : CascadeMux
    port map (
            O => \N__45075\,
            I => \N__45072\
        );

    \I__10201\ : CascadeBuf
    port map (
            O => \N__45072\,
            I => \N__45069\
        );

    \I__10200\ : CascadeMux
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__10199\ : CascadeBuf
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__10198\ : CascadeMux
    port map (
            O => \N__45063\,
            I => \N__45060\
        );

    \I__10197\ : CascadeBuf
    port map (
            O => \N__45060\,
            I => \N__45057\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__45057\,
            I => \N__45054\
        );

    \I__10195\ : CascadeBuf
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__10194\ : CascadeMux
    port map (
            O => \N__45051\,
            I => \N__45048\
        );

    \I__10193\ : CascadeBuf
    port map (
            O => \N__45048\,
            I => \N__45045\
        );

    \I__10192\ : CascadeMux
    port map (
            O => \N__45045\,
            I => \N__45042\
        );

    \I__10191\ : CascadeBuf
    port map (
            O => \N__45042\,
            I => \N__45039\
        );

    \I__10190\ : CascadeMux
    port map (
            O => \N__45039\,
            I => \N__45036\
        );

    \I__10189\ : CascadeBuf
    port map (
            O => \N__45036\,
            I => \N__45032\
        );

    \I__10188\ : CascadeMux
    port map (
            O => \N__45035\,
            I => \N__45029\
        );

    \I__10187\ : CascadeMux
    port map (
            O => \N__45032\,
            I => \N__45026\
        );

    \I__10186\ : CascadeBuf
    port map (
            O => \N__45029\,
            I => \N__45023\
        );

    \I__10185\ : CascadeBuf
    port map (
            O => \N__45026\,
            I => \N__45020\
        );

    \I__10184\ : CascadeMux
    port map (
            O => \N__45023\,
            I => \N__45017\
        );

    \I__10183\ : CascadeMux
    port map (
            O => \N__45020\,
            I => \N__45014\
        );

    \I__10182\ : InMux
    port map (
            O => \N__45017\,
            I => \N__45011\
        );

    \I__10181\ : CascadeBuf
    port map (
            O => \N__45014\,
            I => \N__45008\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__45011\,
            I => \N__45005\
        );

    \I__10179\ : CascadeMux
    port map (
            O => \N__45008\,
            I => \N__45002\
        );

    \I__10178\ : Sp12to4
    port map (
            O => \N__45005\,
            I => \N__44999\
        );

    \I__10177\ : InMux
    port map (
            O => \N__45002\,
            I => \N__44996\
        );

    \I__10176\ : Span12Mux_v
    port map (
            O => \N__44999\,
            I => \N__44993\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__44996\,
            I => \N__44990\
        );

    \I__10174\ : Span12Mux_h
    port map (
            O => \N__44993\,
            I => \N__44987\
        );

    \I__10173\ : Span4Mux_h
    port map (
            O => \N__44990\,
            I => \N__44984\
        );

    \I__10172\ : Odrv12
    port map (
            O => \N__44987\,
            I => \data_index_9_N_216_2\
        );

    \I__10171\ : Odrv4
    port map (
            O => \N__44984\,
            I => \data_index_9_N_216_2\
        );

    \I__10170\ : CascadeMux
    port map (
            O => \N__44979\,
            I => \N__44972\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44967\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44964\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44961\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44975\,
            I => \N__44958\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44972\,
            I => \N__44954\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44971\,
            I => \N__44951\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44970\,
            I => \N__44948\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__44967\,
            I => \N__44942\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44964\,
            I => \N__44942\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44939\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__44958\,
            I => \N__44936\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44928\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__44954\,
            I => \N__44923\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44951\,
            I => \N__44923\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44948\,
            I => \N__44920\
        );

    \I__10154\ : InMux
    port map (
            O => \N__44947\,
            I => \N__44917\
        );

    \I__10153\ : Span4Mux_v
    port map (
            O => \N__44942\,
            I => \N__44910\
        );

    \I__10152\ : Span4Mux_h
    port map (
            O => \N__44939\,
            I => \N__44910\
        );

    \I__10151\ : Span4Mux_v
    port map (
            O => \N__44936\,
            I => \N__44910\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44935\,
            I => \N__44902\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44934\,
            I => \N__44902\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44933\,
            I => \N__44895\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44932\,
            I => \N__44895\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44895\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__44928\,
            I => \N__44890\
        );

    \I__10144\ : Span4Mux_v
    port map (
            O => \N__44923\,
            I => \N__44890\
        );

    \I__10143\ : Span12Mux_v
    port map (
            O => \N__44920\,
            I => \N__44887\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__44917\,
            I => \N__44882\
        );

    \I__10141\ : Span4Mux_h
    port map (
            O => \N__44910\,
            I => \N__44882\
        );

    \I__10140\ : InMux
    port map (
            O => \N__44909\,
            I => \N__44875\
        );

    \I__10139\ : InMux
    port map (
            O => \N__44908\,
            I => \N__44875\
        );

    \I__10138\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44875\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__44902\,
            I => n11819
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44895\,
            I => n11819
        );

    \I__10135\ : Odrv4
    port map (
            O => \N__44890\,
            I => n11819
        );

    \I__10134\ : Odrv12
    port map (
            O => \N__44887\,
            I => n11819
        );

    \I__10133\ : Odrv4
    port map (
            O => \N__44882\,
            I => n11819
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__44875\,
            I => n11819
        );

    \I__10131\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44857\
        );

    \I__10130\ : InMux
    port map (
            O => \N__44861\,
            I => \N__44853\
        );

    \I__10129\ : InMux
    port map (
            O => \N__44860\,
            I => \N__44850\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__44857\,
            I => \N__44846\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44856\,
            I => \N__44843\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__44853\,
            I => \N__44838\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__44850\,
            I => \N__44838\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44835\
        );

    \I__10123\ : Span4Mux_v
    port map (
            O => \N__44846\,
            I => \N__44830\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__44843\,
            I => \N__44830\
        );

    \I__10121\ : Span4Mux_h
    port map (
            O => \N__44838\,
            I => \N__44827\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__44835\,
            I => \N__44824\
        );

    \I__10119\ : Span4Mux_h
    port map (
            O => \N__44830\,
            I => \N__44821\
        );

    \I__10118\ : Span4Mux_h
    port map (
            O => \N__44827\,
            I => \N__44816\
        );

    \I__10117\ : Span12Mux_h
    port map (
            O => \N__44824\,
            I => \N__44813\
        );

    \I__10116\ : Span4Mux_h
    port map (
            O => \N__44821\,
            I => \N__44810\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44820\,
            I => \N__44807\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44804\
        );

    \I__10113\ : Odrv4
    port map (
            O => \N__44816\,
            I => n12381
        );

    \I__10112\ : Odrv12
    port map (
            O => \N__44813\,
            I => n12381
        );

    \I__10111\ : Odrv4
    port map (
            O => \N__44810\,
            I => n12381
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__44807\,
            I => n12381
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44804\,
            I => n12381
        );

    \I__10108\ : CascadeMux
    port map (
            O => \N__44793\,
            I => \N__44789\
        );

    \I__10107\ : CascadeMux
    port map (
            O => \N__44792\,
            I => \N__44783\
        );

    \I__10106\ : InMux
    port map (
            O => \N__44789\,
            I => \N__44780\
        );

    \I__10105\ : CascadeMux
    port map (
            O => \N__44788\,
            I => \N__44776\
        );

    \I__10104\ : InMux
    port map (
            O => \N__44787\,
            I => \N__44773\
        );

    \I__10103\ : CascadeMux
    port map (
            O => \N__44786\,
            I => \N__44770\
        );

    \I__10102\ : InMux
    port map (
            O => \N__44783\,
            I => \N__44766\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__44780\,
            I => \N__44763\
        );

    \I__10100\ : InMux
    port map (
            O => \N__44779\,
            I => \N__44760\
        );

    \I__10099\ : InMux
    port map (
            O => \N__44776\,
            I => \N__44756\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44773\,
            I => \N__44753\
        );

    \I__10097\ : InMux
    port map (
            O => \N__44770\,
            I => \N__44750\
        );

    \I__10096\ : CascadeMux
    port map (
            O => \N__44769\,
            I => \N__44746\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__44766\,
            I => \N__44743\
        );

    \I__10094\ : Span4Mux_v
    port map (
            O => \N__44763\,
            I => \N__44740\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__44760\,
            I => \N__44737\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44759\,
            I => \N__44734\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__44756\,
            I => \N__44729\
        );

    \I__10090\ : Span4Mux_v
    port map (
            O => \N__44753\,
            I => \N__44729\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44750\,
            I => \N__44726\
        );

    \I__10088\ : InMux
    port map (
            O => \N__44749\,
            I => \N__44723\
        );

    \I__10087\ : InMux
    port map (
            O => \N__44746\,
            I => \N__44720\
        );

    \I__10086\ : Span4Mux_v
    port map (
            O => \N__44743\,
            I => \N__44713\
        );

    \I__10085\ : Span4Mux_h
    port map (
            O => \N__44740\,
            I => \N__44713\
        );

    \I__10084\ : Span4Mux_v
    port map (
            O => \N__44737\,
            I => \N__44713\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__44734\,
            I => \N__44710\
        );

    \I__10082\ : Span4Mux_h
    port map (
            O => \N__44729\,
            I => \N__44703\
        );

    \I__10081\ : Span4Mux_h
    port map (
            O => \N__44726\,
            I => \N__44703\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__44723\,
            I => \N__44703\
        );

    \I__10079\ : LocalMux
    port map (
            O => \N__44720\,
            I => \N__44700\
        );

    \I__10078\ : Span4Mux_h
    port map (
            O => \N__44713\,
            I => \N__44695\
        );

    \I__10077\ : Span4Mux_v
    port map (
            O => \N__44710\,
            I => \N__44695\
        );

    \I__10076\ : Span4Mux_v
    port map (
            O => \N__44703\,
            I => \N__44692\
        );

    \I__10075\ : Odrv12
    port map (
            O => \N__44700\,
            I => comm_buf_0_2
        );

    \I__10074\ : Odrv4
    port map (
            O => \N__44695\,
            I => comm_buf_0_2
        );

    \I__10073\ : Odrv4
    port map (
            O => \N__44692\,
            I => comm_buf_0_2
        );

    \I__10072\ : IoInMux
    port map (
            O => \N__44685\,
            I => \N__44682\
        );

    \I__10071\ : LocalMux
    port map (
            O => \N__44682\,
            I => \N__44679\
        );

    \I__10070\ : Span4Mux_s3_v
    port map (
            O => \N__44679\,
            I => \N__44675\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44678\,
            I => \N__44672\
        );

    \I__10068\ : Sp12to4
    port map (
            O => \N__44675\,
            I => \N__44669\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__44672\,
            I => \N__44665\
        );

    \I__10066\ : Span12Mux_h
    port map (
            O => \N__44669\,
            I => \N__44662\
        );

    \I__10065\ : InMux
    port map (
            O => \N__44668\,
            I => \N__44659\
        );

    \I__10064\ : Span4Mux_v
    port map (
            O => \N__44665\,
            I => \N__44656\
        );

    \I__10063\ : Odrv12
    port map (
            O => \N__44662\,
            I => \IAC_FLT0\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__44659\,
            I => \IAC_FLT0\
        );

    \I__10061\ : Odrv4
    port map (
            O => \N__44656\,
            I => \IAC_FLT0\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44646\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__44646\,
            I => \N__44643\
        );

    \I__10058\ : Span4Mux_v
    port map (
            O => \N__44643\,
            I => \N__44640\
        );

    \I__10057\ : Span4Mux_v
    port map (
            O => \N__44640\,
            I => \N__44637\
        );

    \I__10056\ : Span4Mux_v
    port map (
            O => \N__44637\,
            I => \N__44634\
        );

    \I__10055\ : Span4Mux_v
    port map (
            O => \N__44634\,
            I => \N__44629\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44633\,
            I => \N__44626\
        );

    \I__10053\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44623\
        );

    \I__10052\ : Odrv4
    port map (
            O => \N__44629\,
            I => wdtick_flag
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44626\,
            I => wdtick_flag
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__44623\,
            I => wdtick_flag
        );

    \I__10049\ : CascadeMux
    port map (
            O => \N__44616\,
            I => \N__44613\
        );

    \I__10048\ : InMux
    port map (
            O => \N__44613\,
            I => \N__44608\
        );

    \I__10047\ : InMux
    port map (
            O => \N__44612\,
            I => \N__44605\
        );

    \I__10046\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44602\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__44608\,
            I => \N__44599\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__44605\,
            I => buf_control_0
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__44602\,
            I => buf_control_0
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__44599\,
            I => buf_control_0
        );

    \I__10041\ : IoInMux
    port map (
            O => \N__44592\,
            I => \N__44589\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__44589\,
            I => \N__44586\
        );

    \I__10039\ : Span4Mux_s3_v
    port map (
            O => \N__44586\,
            I => \N__44583\
        );

    \I__10038\ : Span4Mux_h
    port map (
            O => \N__44583\,
            I => \N__44580\
        );

    \I__10037\ : Odrv4
    port map (
            O => \N__44580\,
            I => \CONT_SD\
        );

    \I__10036\ : SRMux
    port map (
            O => \N__44577\,
            I => \N__44574\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__44574\,
            I => \N__44571\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__44571\,
            I => \N__44568\
        );

    \I__10033\ : Span4Mux_h
    port map (
            O => \N__44568\,
            I => \N__44565\
        );

    \I__10032\ : Odrv4
    port map (
            O => \N__44565\,
            I => \comm_spi.imosi_N_753\
        );

    \I__10031\ : InMux
    port map (
            O => \N__44562\,
            I => \N__44558\
        );

    \I__10030\ : InMux
    port map (
            O => \N__44561\,
            I => \N__44555\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__44558\,
            I => \N__44550\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__44555\,
            I => \N__44550\
        );

    \I__10027\ : Span4Mux_h
    port map (
            O => \N__44550\,
            I => \N__44547\
        );

    \I__10026\ : Sp12to4
    port map (
            O => \N__44547\,
            I => \N__44543\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44540\
        );

    \I__10024\ : Odrv12
    port map (
            O => \N__44543\,
            I => \comm_spi.n22872\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__44540\,
            I => \comm_spi.n22872\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44532\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44532\,
            I => \N__44529\
        );

    \I__10020\ : Span4Mux_v
    port map (
            O => \N__44529\,
            I => \N__44525\
        );

    \I__10019\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44522\
        );

    \I__10018\ : Odrv4
    port map (
            O => \N__44525\,
            I => \comm_spi.n14630\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__44522\,
            I => \comm_spi.n14630\
        );

    \I__10016\ : InMux
    port map (
            O => \N__44517\,
            I => \N__44513\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44510\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__44513\,
            I => \N__44505\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__44510\,
            I => \N__44505\
        );

    \I__10012\ : Span4Mux_v
    port map (
            O => \N__44505\,
            I => \N__44502\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__44502\,
            I => \comm_spi.n14631\
        );

    \I__10010\ : SRMux
    port map (
            O => \N__44499\,
            I => \N__44496\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__44496\,
            I => \N__44493\
        );

    \I__10008\ : Span4Mux_v
    port map (
            O => \N__44493\,
            I => \N__44490\
        );

    \I__10007\ : Odrv4
    port map (
            O => \N__44490\,
            I => \comm_spi.data_tx_7__N_768\
        );

    \I__10006\ : InMux
    port map (
            O => \N__44487\,
            I => \N__44482\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44479\
        );

    \I__10004\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44476\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__44482\,
            I => \comm_spi.n22869\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__44479\,
            I => \comm_spi.n22869\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__44476\,
            I => \comm_spi.n22869\
        );

    \I__10000\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44465\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44468\,
            I => \N__44462\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__44465\,
            I => \comm_spi.n14634\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__44462\,
            I => \comm_spi.n14634\
        );

    \I__9996\ : InMux
    port map (
            O => \N__44457\,
            I => \N__44453\
        );

    \I__9995\ : InMux
    port map (
            O => \N__44456\,
            I => \N__44450\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44453\,
            I => \comm_spi.n14635\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__44450\,
            I => \comm_spi.n14635\
        );

    \I__9992\ : InMux
    port map (
            O => \N__44445\,
            I => \N__44442\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__44442\,
            I => \N__44438\
        );

    \I__9990\ : InMux
    port map (
            O => \N__44441\,
            I => \N__44435\
        );

    \I__9989\ : Sp12to4
    port map (
            O => \N__44438\,
            I => \N__44430\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__44435\,
            I => \N__44430\
        );

    \I__9987\ : Odrv12
    port map (
            O => \N__44430\,
            I => \comm_spi.n14638\
        );

    \I__9986\ : InMux
    port map (
            O => \N__44427\,
            I => \N__44423\
        );

    \I__9985\ : InMux
    port map (
            O => \N__44426\,
            I => \N__44420\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44423\,
            I => \N__44415\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__44420\,
            I => \N__44415\
        );

    \I__9982\ : Span4Mux_v
    port map (
            O => \N__44415\,
            I => \N__44412\
        );

    \I__9981\ : Odrv4
    port map (
            O => \N__44412\,
            I => n14_adj_1578
        );

    \I__9980\ : CascadeMux
    port map (
            O => \N__44409\,
            I => \N__44406\
        );

    \I__9979\ : InMux
    port map (
            O => \N__44406\,
            I => \N__44403\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__44403\,
            I => \N__44400\
        );

    \I__9977\ : Span4Mux_v
    port map (
            O => \N__44400\,
            I => \N__44397\
        );

    \I__9976\ : Odrv4
    port map (
            O => \N__44397\,
            I => n9_adj_1415
        );

    \I__9975\ : CascadeMux
    port map (
            O => \N__44394\,
            I => \N__44391\
        );

    \I__9974\ : InMux
    port map (
            O => \N__44391\,
            I => \N__44388\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__44388\,
            I => \N__44385\
        );

    \I__9972\ : Span4Mux_h
    port map (
            O => \N__44385\,
            I => \N__44382\
        );

    \I__9971\ : Span4Mux_v
    port map (
            O => \N__44382\,
            I => \N__44379\
        );

    \I__9970\ : Odrv4
    port map (
            O => \N__44379\,
            I => buf_data_iac_16
        );

    \I__9969\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44373\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__44373\,
            I => n21165
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__44370\,
            I => \n21167_cascade_\
        );

    \I__9966\ : InMux
    port map (
            O => \N__44367\,
            I => \N__44364\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__44364\,
            I => n22222
        );

    \I__9964\ : CascadeMux
    port map (
            O => \N__44361\,
            I => \N__44358\
        );

    \I__9963\ : InMux
    port map (
            O => \N__44358\,
            I => \N__44355\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__44355\,
            I => n21070
        );

    \I__9961\ : InMux
    port map (
            O => \N__44352\,
            I => \N__44349\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__44349\,
            I => n21084
        );

    \I__9959\ : InMux
    port map (
            O => \N__44346\,
            I => \N__44343\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__44343\,
            I => n21085
        );

    \I__9957\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44337\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__44337\,
            I => \N__44334\
        );

    \I__9955\ : Odrv4
    port map (
            O => \N__44334\,
            I => n22309
        );

    \I__9954\ : CascadeMux
    port map (
            O => \N__44331\,
            I => \N__44318\
        );

    \I__9953\ : InMux
    port map (
            O => \N__44330\,
            I => \N__44311\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44311\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44308\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44303\
        );

    \I__9949\ : InMux
    port map (
            O => \N__44326\,
            I => \N__44303\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44300\
        );

    \I__9947\ : InMux
    port map (
            O => \N__44324\,
            I => \N__44288\
        );

    \I__9946\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44288\
        );

    \I__9945\ : InMux
    port map (
            O => \N__44322\,
            I => \N__44288\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44288\
        );

    \I__9943\ : InMux
    port map (
            O => \N__44318\,
            I => \N__44285\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44317\,
            I => \N__44282\
        );

    \I__9941\ : InMux
    port map (
            O => \N__44316\,
            I => \N__44279\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__44311\,
            I => \N__44276\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__44308\,
            I => \N__44271\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__44303\,
            I => \N__44271\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__44300\,
            I => \N__44268\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44299\,
            I => \N__44261\
        );

    \I__9935\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44261\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44297\,
            I => \N__44261\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44258\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__44285\,
            I => \N__44253\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__44282\,
            I => \N__44253\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__44279\,
            I => \N__44248\
        );

    \I__9929\ : Span4Mux_v
    port map (
            O => \N__44276\,
            I => \N__44248\
        );

    \I__9928\ : Span4Mux_v
    port map (
            O => \N__44271\,
            I => \N__44245\
        );

    \I__9927\ : Span4Mux_v
    port map (
            O => \N__44268\,
            I => \N__44242\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__44261\,
            I => n12399
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__44258\,
            I => n12399
        );

    \I__9924\ : Odrv12
    port map (
            O => \N__44253\,
            I => n12399
        );

    \I__9923\ : Odrv4
    port map (
            O => \N__44248\,
            I => n12399
        );

    \I__9922\ : Odrv4
    port map (
            O => \N__44245\,
            I => n12399
        );

    \I__9921\ : Odrv4
    port map (
            O => \N__44242\,
            I => n12399
        );

    \I__9920\ : CascadeMux
    port map (
            O => \N__44229\,
            I => \N__44223\
        );

    \I__9919\ : CascadeMux
    port map (
            O => \N__44228\,
            I => \N__44219\
        );

    \I__9918\ : CascadeMux
    port map (
            O => \N__44227\,
            I => \N__44216\
        );

    \I__9917\ : CascadeMux
    port map (
            O => \N__44226\,
            I => \N__44213\
        );

    \I__9916\ : InMux
    port map (
            O => \N__44223\,
            I => \N__44210\
        );

    \I__9915\ : InMux
    port map (
            O => \N__44222\,
            I => \N__44207\
        );

    \I__9914\ : InMux
    port map (
            O => \N__44219\,
            I => \N__44204\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44201\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44198\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__44210\,
            I => \N__44194\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44207\,
            I => \N__44191\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__44204\,
            I => \N__44188\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__44201\,
            I => \N__44184\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__44198\,
            I => \N__44181\
        );

    \I__9906\ : CascadeMux
    port map (
            O => \N__44197\,
            I => \N__44178\
        );

    \I__9905\ : Span4Mux_h
    port map (
            O => \N__44194\,
            I => \N__44174\
        );

    \I__9904\ : Span4Mux_v
    port map (
            O => \N__44191\,
            I => \N__44171\
        );

    \I__9903\ : Span4Mux_h
    port map (
            O => \N__44188\,
            I => \N__44168\
        );

    \I__9902\ : InMux
    port map (
            O => \N__44187\,
            I => \N__44165\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__44184\,
            I => \N__44160\
        );

    \I__9900\ : Span4Mux_v
    port map (
            O => \N__44181\,
            I => \N__44160\
        );

    \I__9899\ : InMux
    port map (
            O => \N__44178\,
            I => \N__44157\
        );

    \I__9898\ : InMux
    port map (
            O => \N__44177\,
            I => \N__44154\
        );

    \I__9897\ : Span4Mux_h
    port map (
            O => \N__44174\,
            I => \N__44151\
        );

    \I__9896\ : Span4Mux_h
    port map (
            O => \N__44171\,
            I => \N__44148\
        );

    \I__9895\ : Span4Mux_h
    port map (
            O => \N__44168\,
            I => \N__44143\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__44165\,
            I => \N__44143\
        );

    \I__9893\ : Span4Mux_h
    port map (
            O => \N__44160\,
            I => \N__44140\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__44157\,
            I => \N__44133\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__44154\,
            I => \N__44133\
        );

    \I__9890\ : Span4Mux_h
    port map (
            O => \N__44151\,
            I => \N__44133\
        );

    \I__9889\ : Span4Mux_v
    port map (
            O => \N__44148\,
            I => \N__44128\
        );

    \I__9888\ : Span4Mux_v
    port map (
            O => \N__44143\,
            I => \N__44128\
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__44140\,
            I => comm_buf_0_3
        );

    \I__9886\ : Odrv4
    port map (
            O => \N__44133\,
            I => comm_buf_0_3
        );

    \I__9885\ : Odrv4
    port map (
            O => \N__44128\,
            I => comm_buf_0_3
        );

    \I__9884\ : IoInMux
    port map (
            O => \N__44121\,
            I => \N__44118\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__44118\,
            I => \N__44115\
        );

    \I__9882\ : Span4Mux_s3_v
    port map (
            O => \N__44115\,
            I => \N__44112\
        );

    \I__9881\ : Span4Mux_v
    port map (
            O => \N__44112\,
            I => \N__44109\
        );

    \I__9880\ : Sp12to4
    port map (
            O => \N__44109\,
            I => \N__44105\
        );

    \I__9879\ : InMux
    port map (
            O => \N__44108\,
            I => \N__44101\
        );

    \I__9878\ : Span12Mux_h
    port map (
            O => \N__44105\,
            I => \N__44098\
        );

    \I__9877\ : InMux
    port map (
            O => \N__44104\,
            I => \N__44095\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__44101\,
            I => \N__44092\
        );

    \I__9875\ : Odrv12
    port map (
            O => \N__44098\,
            I => \IAC_FLT1\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__44095\,
            I => \IAC_FLT1\
        );

    \I__9873\ : Odrv4
    port map (
            O => \N__44092\,
            I => \IAC_FLT1\
        );

    \I__9872\ : InMux
    port map (
            O => \N__44085\,
            I => \N__44082\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__44082\,
            I => \N__44079\
        );

    \I__9870\ : Span12Mux_h
    port map (
            O => \N__44079\,
            I => \N__44076\
        );

    \I__9869\ : Odrv12
    port map (
            O => \N__44076\,
            I => n20914
        );

    \I__9868\ : CascadeMux
    port map (
            O => \N__44073\,
            I => \N__44070\
        );

    \I__9867\ : InMux
    port map (
            O => \N__44070\,
            I => \N__44066\
        );

    \I__9866\ : CascadeMux
    port map (
            O => \N__44069\,
            I => \N__44063\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__44066\,
            I => \N__44060\
        );

    \I__9864\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44056\
        );

    \I__9863\ : Span4Mux_v
    port map (
            O => \N__44060\,
            I => \N__44053\
        );

    \I__9862\ : CascadeMux
    port map (
            O => \N__44059\,
            I => \N__44050\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__44056\,
            I => \N__44047\
        );

    \I__9860\ : Span4Mux_h
    port map (
            O => \N__44053\,
            I => \N__44044\
        );

    \I__9859\ : InMux
    port map (
            O => \N__44050\,
            I => \N__44041\
        );

    \I__9858\ : Span4Mux_h
    port map (
            O => \N__44047\,
            I => \N__44038\
        );

    \I__9857\ : Span4Mux_h
    port map (
            O => \N__44044\,
            I => \N__44033\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__44041\,
            I => \N__44033\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__44038\,
            I => \N__44029\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__44033\,
            I => \N__44026\
        );

    \I__9853\ : CascadeMux
    port map (
            O => \N__44032\,
            I => \N__44023\
        );

    \I__9852\ : Span4Mux_h
    port map (
            O => \N__44029\,
            I => \N__44020\
        );

    \I__9851\ : Span4Mux_v
    port map (
            O => \N__44026\,
            I => \N__44017\
        );

    \I__9850\ : InMux
    port map (
            O => \N__44023\,
            I => \N__44014\
        );

    \I__9849\ : Span4Mux_h
    port map (
            O => \N__44020\,
            I => \N__44011\
        );

    \I__9848\ : Span4Mux_v
    port map (
            O => \N__44017\,
            I => \N__44008\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__44014\,
            I => trig_dds1
        );

    \I__9846\ : Odrv4
    port map (
            O => \N__44011\,
            I => trig_dds1
        );

    \I__9845\ : Odrv4
    port map (
            O => \N__44008\,
            I => trig_dds1
        );

    \I__9844\ : InMux
    port map (
            O => \N__44001\,
            I => \N__43997\
        );

    \I__9843\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43994\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__43997\,
            I => \N__43990\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43994\,
            I => \N__43987\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43993\,
            I => \N__43984\
        );

    \I__9839\ : Span4Mux_h
    port map (
            O => \N__43990\,
            I => \N__43981\
        );

    \I__9838\ : Odrv4
    port map (
            O => \N__43987\,
            I => buf_dds0_11
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__43984\,
            I => buf_dds0_11
        );

    \I__9836\ : Odrv4
    port map (
            O => \N__43981\,
            I => buf_dds0_11
        );

    \I__9835\ : CascadeMux
    port map (
            O => \N__43974\,
            I => \n22297_cascade_\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43971\,
            I => \N__43967\
        );

    \I__9833\ : InMux
    port map (
            O => \N__43970\,
            I => \N__43963\
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__43967\,
            I => \N__43960\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43966\,
            I => \N__43957\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__43963\,
            I => \N__43954\
        );

    \I__9829\ : Span12Mux_h
    port map (
            O => \N__43960\,
            I => \N__43951\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43957\,
            I => \N__43946\
        );

    \I__9827\ : Span4Mux_h
    port map (
            O => \N__43954\,
            I => \N__43946\
        );

    \I__9826\ : Odrv12
    port map (
            O => \N__43951\,
            I => buf_dds1_11
        );

    \I__9825\ : Odrv4
    port map (
            O => \N__43946\,
            I => buf_dds1_11
        );

    \I__9824\ : InMux
    port map (
            O => \N__43941\,
            I => \N__43938\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43938\,
            I => \N__43935\
        );

    \I__9822\ : Odrv12
    port map (
            O => \N__43935\,
            I => n21076
        );

    \I__9821\ : CascadeMux
    port map (
            O => \N__43932\,
            I => \N__43929\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43926\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__43926\,
            I => n22300
        );

    \I__9818\ : CascadeMux
    port map (
            O => \N__43923\,
            I => \n22312_cascade_\
        );

    \I__9817\ : CascadeMux
    port map (
            O => \N__43920\,
            I => \N__43917\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43914\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43914\,
            I => \N__43911\
        );

    \I__9814\ : Span4Mux_h
    port map (
            O => \N__43911\,
            I => \N__43907\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43910\,
            I => \N__43901\
        );

    \I__9812\ : Span4Mux_h
    port map (
            O => \N__43907\,
            I => \N__43898\
        );

    \I__9811\ : InMux
    port map (
            O => \N__43906\,
            I => \N__43895\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43905\,
            I => \N__43890\
        );

    \I__9809\ : InMux
    port map (
            O => \N__43904\,
            I => \N__43890\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__43901\,
            I => eis_start
        );

    \I__9807\ : Odrv4
    port map (
            O => \N__43898\,
            I => eis_start
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__43895\,
            I => eis_start
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__43890\,
            I => eis_start
        );

    \I__9804\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43878\,
            I => \N__43873\
        );

    \I__9802\ : CascadeMux
    port map (
            O => \N__43877\,
            I => \N__43870\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43876\,
            I => \N__43867\
        );

    \I__9800\ : Span4Mux_h
    port map (
            O => \N__43873\,
            I => \N__43864\
        );

    \I__9799\ : InMux
    port map (
            O => \N__43870\,
            I => \N__43861\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43867\,
            I => req_data_cnt_8
        );

    \I__9797\ : Odrv4
    port map (
            O => \N__43864\,
            I => req_data_cnt_8
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__43861\,
            I => req_data_cnt_8
        );

    \I__9795\ : InMux
    port map (
            O => \N__43854\,
            I => \N__43851\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__43851\,
            I => \N__43848\
        );

    \I__9793\ : Span4Mux_h
    port map (
            O => \N__43848\,
            I => \N__43845\
        );

    \I__9792\ : Span4Mux_h
    port map (
            O => \N__43845\,
            I => \N__43842\
        );

    \I__9791\ : Odrv4
    port map (
            O => \N__43842\,
            I => n22294
        );

    \I__9790\ : CascadeMux
    port map (
            O => \N__43839\,
            I => \n21071_cascade_\
        );

    \I__9789\ : CascadeMux
    port map (
            O => \N__43836\,
            I => \N__43832\
        );

    \I__9788\ : CascadeMux
    port map (
            O => \N__43835\,
            I => \N__43826\
        );

    \I__9787\ : InMux
    port map (
            O => \N__43832\,
            I => \N__43819\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43831\,
            I => \N__43819\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43830\,
            I => \N__43816\
        );

    \I__9784\ : CascadeMux
    port map (
            O => \N__43829\,
            I => \N__43812\
        );

    \I__9783\ : InMux
    port map (
            O => \N__43826\,
            I => \N__43809\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43805\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43802\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__43819\,
            I => \N__43799\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43816\,
            I => \N__43796\
        );

    \I__9778\ : InMux
    port map (
            O => \N__43815\,
            I => \N__43793\
        );

    \I__9777\ : InMux
    port map (
            O => \N__43812\,
            I => \N__43790\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43809\,
            I => \N__43787\
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__43808\,
            I => \N__43784\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__43805\,
            I => \N__43780\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__43802\,
            I => \N__43775\
        );

    \I__9772\ : Span4Mux_v
    port map (
            O => \N__43799\,
            I => \N__43775\
        );

    \I__9771\ : Span4Mux_v
    port map (
            O => \N__43796\,
            I => \N__43770\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__43793\,
            I => \N__43770\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43790\,
            I => \N__43767\
        );

    \I__9768\ : Span4Mux_h
    port map (
            O => \N__43787\,
            I => \N__43764\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43784\,
            I => \N__43761\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43783\,
            I => \N__43758\
        );

    \I__9765\ : Span4Mux_v
    port map (
            O => \N__43780\,
            I => \N__43755\
        );

    \I__9764\ : Span4Mux_h
    port map (
            O => \N__43775\,
            I => \N__43750\
        );

    \I__9763\ : Span4Mux_h
    port map (
            O => \N__43770\,
            I => \N__43750\
        );

    \I__9762\ : Span4Mux_h
    port map (
            O => \N__43767\,
            I => \N__43745\
        );

    \I__9761\ : Span4Mux_v
    port map (
            O => \N__43764\,
            I => \N__43745\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__43761\,
            I => \N__43740\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__43758\,
            I => \N__43740\
        );

    \I__9758\ : Span4Mux_v
    port map (
            O => \N__43755\,
            I => \N__43735\
        );

    \I__9757\ : Span4Mux_h
    port map (
            O => \N__43750\,
            I => \N__43735\
        );

    \I__9756\ : Span4Mux_h
    port map (
            O => \N__43745\,
            I => \N__43730\
        );

    \I__9755\ : Span4Mux_v
    port map (
            O => \N__43740\,
            I => \N__43730\
        );

    \I__9754\ : Odrv4
    port map (
            O => \N__43735\,
            I => comm_buf_0_0
        );

    \I__9753\ : Odrv4
    port map (
            O => \N__43730\,
            I => comm_buf_0_0
        );

    \I__9752\ : SRMux
    port map (
            O => \N__43725\,
            I => \N__43720\
        );

    \I__9751\ : SRMux
    port map (
            O => \N__43724\,
            I => \N__43717\
        );

    \I__9750\ : SRMux
    port map (
            O => \N__43723\,
            I => \N__43714\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__43720\,
            I => \N__43711\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43717\,
            I => \N__43707\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43714\,
            I => \N__43704\
        );

    \I__9746\ : Span4Mux_h
    port map (
            O => \N__43711\,
            I => \N__43701\
        );

    \I__9745\ : SRMux
    port map (
            O => \N__43710\,
            I => \N__43695\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__43707\,
            I => \N__43690\
        );

    \I__9743\ : Span4Mux_v
    port map (
            O => \N__43704\,
            I => \N__43690\
        );

    \I__9742\ : Span4Mux_h
    port map (
            O => \N__43701\,
            I => \N__43687\
        );

    \I__9741\ : SRMux
    port map (
            O => \N__43700\,
            I => \N__43684\
        );

    \I__9740\ : SRMux
    port map (
            O => \N__43699\,
            I => \N__43681\
        );

    \I__9739\ : SRMux
    port map (
            O => \N__43698\,
            I => \N__43678\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__43695\,
            I => \N__43675\
        );

    \I__9737\ : Sp12to4
    port map (
            O => \N__43690\,
            I => \N__43672\
        );

    \I__9736\ : Span4Mux_v
    port map (
            O => \N__43687\,
            I => \N__43669\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__43684\,
            I => n14750
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43681\,
            I => n14750
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__43678\,
            I => n14750
        );

    \I__9732\ : Odrv12
    port map (
            O => \N__43675\,
            I => n14750
        );

    \I__9731\ : Odrv12
    port map (
            O => \N__43672\,
            I => n14750
        );

    \I__9730\ : Odrv4
    port map (
            O => \N__43669\,
            I => n14750
        );

    \I__9729\ : InMux
    port map (
            O => \N__43656\,
            I => \N__43653\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__43653\,
            I => n22219
        );

    \I__9727\ : InMux
    port map (
            O => \N__43650\,
            I => \N__43646\
        );

    \I__9726\ : InMux
    port map (
            O => \N__43649\,
            I => \N__43643\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__43646\,
            I => \N__43640\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__43643\,
            I => \N__43636\
        );

    \I__9723\ : Span12Mux_h
    port map (
            O => \N__43640\,
            I => \N__43633\
        );

    \I__9722\ : InMux
    port map (
            O => \N__43639\,
            I => \N__43630\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__43636\,
            I => \acadc_skipCount_8\
        );

    \I__9720\ : Odrv12
    port map (
            O => \N__43633\,
            I => \acadc_skipCount_8\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__43630\,
            I => \acadc_skipCount_8\
        );

    \I__9718\ : InMux
    port map (
            O => \N__43623\,
            I => \N__43620\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43620\,
            I => \N__43617\
        );

    \I__9716\ : Span4Mux_v
    port map (
            O => \N__43617\,
            I => \N__43614\
        );

    \I__9715\ : Span4Mux_h
    port map (
            O => \N__43614\,
            I => \N__43611\
        );

    \I__9714\ : Span4Mux_h
    port map (
            O => \N__43611\,
            I => \N__43608\
        );

    \I__9713\ : Odrv4
    port map (
            O => \N__43608\,
            I => n22324
        );

    \I__9712\ : CascadeMux
    port map (
            O => \N__43605\,
            I => \N__43602\
        );

    \I__9711\ : InMux
    port map (
            O => \N__43602\,
            I => \N__43597\
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__43601\,
            I => \N__43594\
        );

    \I__9709\ : CascadeMux
    port map (
            O => \N__43600\,
            I => \N__43590\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43586\
        );

    \I__9707\ : InMux
    port map (
            O => \N__43594\,
            I => \N__43583\
        );

    \I__9706\ : InMux
    port map (
            O => \N__43593\,
            I => \N__43580\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43590\,
            I => \N__43577\
        );

    \I__9704\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43574\
        );

    \I__9703\ : Span4Mux_v
    port map (
            O => \N__43586\,
            I => \N__43569\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__43583\,
            I => \N__43569\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__43580\,
            I => \N__43564\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__43577\,
            I => \N__43561\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__43574\,
            I => \N__43556\
        );

    \I__9698\ : Span4Mux_h
    port map (
            O => \N__43569\,
            I => \N__43556\
        );

    \I__9697\ : InMux
    port map (
            O => \N__43568\,
            I => \N__43553\
        );

    \I__9696\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43550\
        );

    \I__9695\ : Span4Mux_v
    port map (
            O => \N__43564\,
            I => \N__43547\
        );

    \I__9694\ : Span12Mux_v
    port map (
            O => \N__43561\,
            I => \N__43544\
        );

    \I__9693\ : Sp12to4
    port map (
            O => \N__43556\,
            I => \N__43539\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__43553\,
            I => \N__43539\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__43550\,
            I => \N__43536\
        );

    \I__9690\ : Sp12to4
    port map (
            O => \N__43547\,
            I => \N__43531\
        );

    \I__9689\ : Span12Mux_h
    port map (
            O => \N__43544\,
            I => \N__43531\
        );

    \I__9688\ : Span12Mux_v
    port map (
            O => \N__43539\,
            I => \N__43528\
        );

    \I__9687\ : Odrv4
    port map (
            O => \N__43536\,
            I => comm_buf_0_5
        );

    \I__9686\ : Odrv12
    port map (
            O => \N__43531\,
            I => comm_buf_0_5
        );

    \I__9685\ : Odrv12
    port map (
            O => \N__43528\,
            I => comm_buf_0_5
        );

    \I__9684\ : CascadeMux
    port map (
            O => \N__43521\,
            I => \N__43518\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43514\
        );

    \I__9682\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43511\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__43514\,
            I => \N__43508\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__43511\,
            I => \N__43505\
        );

    \I__9679\ : Span4Mux_v
    port map (
            O => \N__43508\,
            I => \N__43499\
        );

    \I__9678\ : Span4Mux_v
    port map (
            O => \N__43505\,
            I => \N__43499\
        );

    \I__9677\ : CascadeMux
    port map (
            O => \N__43504\,
            I => \N__43496\
        );

    \I__9676\ : Sp12to4
    port map (
            O => \N__43499\,
            I => \N__43493\
        );

    \I__9675\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43490\
        );

    \I__9674\ : Span12Mux_h
    port map (
            O => \N__43493\,
            I => \N__43487\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__43490\,
            I => buf_adcdata_iac_8
        );

    \I__9672\ : Odrv12
    port map (
            O => \N__43487\,
            I => buf_adcdata_iac_8
        );

    \I__9671\ : InMux
    port map (
            O => \N__43482\,
            I => \N__43479\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43479\,
            I => \N__43476\
        );

    \I__9669\ : Span4Mux_v
    port map (
            O => \N__43476\,
            I => \N__43473\
        );

    \I__9668\ : Span4Mux_h
    port map (
            O => \N__43473\,
            I => \N__43470\
        );

    \I__9667\ : Odrv4
    port map (
            O => \N__43470\,
            I => n16_adj_1487
        );

    \I__9666\ : InMux
    port map (
            O => \N__43467\,
            I => \N__43464\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__43464\,
            I => \N__43461\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__43461\,
            I => \N__43458\
        );

    \I__9663\ : Span4Mux_h
    port map (
            O => \N__43458\,
            I => \N__43455\
        );

    \I__9662\ : Span4Mux_h
    port map (
            O => \N__43455\,
            I => \N__43452\
        );

    \I__9661\ : Odrv4
    port map (
            O => \N__43452\,
            I => n19_adj_1486
        );

    \I__9660\ : CascadeMux
    port map (
            O => \N__43449\,
            I => \N__43446\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43446\,
            I => \N__43443\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__43443\,
            I => \N__43440\
        );

    \I__9657\ : Span12Mux_v
    port map (
            O => \N__43440\,
            I => \N__43436\
        );

    \I__9656\ : CascadeMux
    port map (
            O => \N__43439\,
            I => \N__43433\
        );

    \I__9655\ : Span12Mux_h
    port map (
            O => \N__43436\,
            I => \N__43430\
        );

    \I__9654\ : InMux
    port map (
            O => \N__43433\,
            I => \N__43427\
        );

    \I__9653\ : Odrv12
    port map (
            O => \N__43430\,
            I => \buf_readRTD_0\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__43427\,
            I => \buf_readRTD_0\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43422\,
            I => \N__43419\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__43419\,
            I => n22213
        );

    \I__9649\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43413\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__43413\,
            I => \N__43409\
        );

    \I__9647\ : CascadeMux
    port map (
            O => \N__43412\,
            I => \N__43406\
        );

    \I__9646\ : Span4Mux_v
    port map (
            O => \N__43409\,
            I => \N__43403\
        );

    \I__9645\ : InMux
    port map (
            O => \N__43406\,
            I => \N__43400\
        );

    \I__9644\ : Span4Mux_h
    port map (
            O => \N__43403\,
            I => \N__43397\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__43400\,
            I => data_idxvec_0
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__43397\,
            I => data_idxvec_0
        );

    \I__9641\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43388\
        );

    \I__9640\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43384\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__43388\,
            I => \N__43381\
        );

    \I__9638\ : InMux
    port map (
            O => \N__43387\,
            I => \N__43378\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43373\
        );

    \I__9636\ : Span4Mux_h
    port map (
            O => \N__43381\,
            I => \N__43373\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__43378\,
            I => data_cntvec_0
        );

    \I__9634\ : Odrv4
    port map (
            O => \N__43373\,
            I => data_cntvec_0
        );

    \I__9633\ : CascadeMux
    port map (
            O => \N__43368\,
            I => \n26_cascade_\
        );

    \I__9632\ : InMux
    port map (
            O => \N__43365\,
            I => \N__43362\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__43362\,
            I => \N__43358\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43361\,
            I => \N__43354\
        );

    \I__9629\ : Span4Mux_v
    port map (
            O => \N__43358\,
            I => \N__43351\
        );

    \I__9628\ : InMux
    port map (
            O => \N__43357\,
            I => \N__43348\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43354\,
            I => \acadc_skipCount_0\
        );

    \I__9626\ : Odrv4
    port map (
            O => \N__43351\,
            I => \acadc_skipCount_0\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__43348\,
            I => \acadc_skipCount_0\
        );

    \I__9624\ : CascadeMux
    port map (
            O => \N__43341\,
            I => \n22201_cascade_\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43338\,
            I => \N__43335\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__43335\,
            I => \N__43330\
        );

    \I__9621\ : CascadeMux
    port map (
            O => \N__43334\,
            I => \N__43327\
        );

    \I__9620\ : CascadeMux
    port map (
            O => \N__43333\,
            I => \N__43324\
        );

    \I__9619\ : Span4Mux_v
    port map (
            O => \N__43330\,
            I => \N__43321\
        );

    \I__9618\ : InMux
    port map (
            O => \N__43327\,
            I => \N__43316\
        );

    \I__9617\ : InMux
    port map (
            O => \N__43324\,
            I => \N__43316\
        );

    \I__9616\ : Odrv4
    port map (
            O => \N__43321\,
            I => req_data_cnt_0
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__43316\,
            I => req_data_cnt_0
        );

    \I__9614\ : InMux
    port map (
            O => \N__43311\,
            I => \N__43308\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__43308\,
            I => n22216
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__43305\,
            I => \n22204_cascade_\
        );

    \I__9611\ : CascadeMux
    port map (
            O => \N__43302\,
            I => \n30_adj_1485_cascade_\
        );

    \I__9610\ : CascadeMux
    port map (
            O => \N__43299\,
            I => \N__43296\
        );

    \I__9609\ : InMux
    port map (
            O => \N__43296\,
            I => \N__43293\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__43293\,
            I => \N__43287\
        );

    \I__9607\ : InMux
    port map (
            O => \N__43292\,
            I => \N__43284\
        );

    \I__9606\ : InMux
    port map (
            O => \N__43291\,
            I => \N__43279\
        );

    \I__9605\ : InMux
    port map (
            O => \N__43290\,
            I => \N__43276\
        );

    \I__9604\ : Span4Mux_v
    port map (
            O => \N__43287\,
            I => \N__43271\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__43284\,
            I => \N__43271\
        );

    \I__9602\ : InMux
    port map (
            O => \N__43283\,
            I => \N__43268\
        );

    \I__9601\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43265\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__43279\,
            I => \N__43262\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__43276\,
            I => \N__43259\
        );

    \I__9598\ : Span4Mux_v
    port map (
            O => \N__43271\,
            I => \N__43254\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__43268\,
            I => \N__43254\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__43265\,
            I => \N__43251\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__43262\,
            I => \N__43248\
        );

    \I__9594\ : Span4Mux_v
    port map (
            O => \N__43259\,
            I => \N__43243\
        );

    \I__9593\ : Span4Mux_v
    port map (
            O => \N__43254\,
            I => \N__43243\
        );

    \I__9592\ : Span4Mux_v
    port map (
            O => \N__43251\,
            I => \N__43240\
        );

    \I__9591\ : Span4Mux_v
    port map (
            O => \N__43248\,
            I => \N__43235\
        );

    \I__9590\ : Span4Mux_h
    port map (
            O => \N__43243\,
            I => \N__43235\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__43240\,
            I => comm_buf_1_0
        );

    \I__9588\ : Odrv4
    port map (
            O => \N__43235\,
            I => comm_buf_1_0
        );

    \I__9587\ : InMux
    port map (
            O => \N__43230\,
            I => \N__43226\
        );

    \I__9586\ : CascadeMux
    port map (
            O => \N__43229\,
            I => \N__43223\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__43226\,
            I => \N__43220\
        );

    \I__9584\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43217\
        );

    \I__9583\ : Span12Mux_v
    port map (
            O => \N__43220\,
            I => \N__43213\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43217\,
            I => \N__43210\
        );

    \I__9581\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43207\
        );

    \I__9580\ : Span12Mux_h
    port map (
            O => \N__43213\,
            I => \N__43204\
        );

    \I__9579\ : Span12Mux_v
    port map (
            O => \N__43210\,
            I => \N__43201\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__43207\,
            I => buf_adcdata_iac_19
        );

    \I__9577\ : Odrv12
    port map (
            O => \N__43204\,
            I => buf_adcdata_iac_19
        );

    \I__9576\ : Odrv12
    port map (
            O => \N__43201\,
            I => buf_adcdata_iac_19
        );

    \I__9575\ : InMux
    port map (
            O => \N__43194\,
            I => \N__43191\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__43191\,
            I => comm_buf_4_1
        );

    \I__9573\ : InMux
    port map (
            O => \N__43188\,
            I => \N__43185\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__43185\,
            I => \N__43181\
        );

    \I__9571\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43178\
        );

    \I__9570\ : Span4Mux_h
    port map (
            O => \N__43181\,
            I => \N__43175\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__43178\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__9568\ : Odrv4
    port map (
            O => \N__43175\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__9567\ : InMux
    port map (
            O => \N__43170\,
            I => \N__43161\
        );

    \I__9566\ : InMux
    port map (
            O => \N__43169\,
            I => \N__43161\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43168\,
            I => \N__43161\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__43161\,
            I => \N__43158\
        );

    \I__9563\ : Span4Mux_v
    port map (
            O => \N__43158\,
            I => \N__43154\
        );

    \I__9562\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43151\
        );

    \I__9561\ : Span4Mux_h
    port map (
            O => \N__43154\,
            I => \N__43147\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__43151\,
            I => \N__43144\
        );

    \I__9559\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43141\
        );

    \I__9558\ : Odrv4
    port map (
            O => \N__43147\,
            I => bit_cnt_0
        );

    \I__9557\ : Odrv4
    port map (
            O => \N__43144\,
            I => bit_cnt_0
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__43141\,
            I => bit_cnt_0
        );

    \I__9555\ : InMux
    port map (
            O => \N__43134\,
            I => \N__43131\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__43131\,
            I => \N__43128\
        );

    \I__9553\ : Span4Mux_v
    port map (
            O => \N__43128\,
            I => \N__43123\
        );

    \I__9552\ : CascadeMux
    port map (
            O => \N__43127\,
            I => \N__43120\
        );

    \I__9551\ : CascadeMux
    port map (
            O => \N__43126\,
            I => \N__43117\
        );

    \I__9550\ : Sp12to4
    port map (
            O => \N__43123\,
            I => \N__43113\
        );

    \I__9549\ : InMux
    port map (
            O => \N__43120\,
            I => \N__43106\
        );

    \I__9548\ : InMux
    port map (
            O => \N__43117\,
            I => \N__43106\
        );

    \I__9547\ : InMux
    port map (
            O => \N__43116\,
            I => \N__43106\
        );

    \I__9546\ : Span12Mux_v
    port map (
            O => \N__43113\,
            I => \N__43103\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__43106\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__9544\ : Odrv12
    port map (
            O => \N__43103\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__9543\ : CascadeMux
    port map (
            O => \N__43098\,
            I => \N__43095\
        );

    \I__9542\ : InMux
    port map (
            O => \N__43095\,
            I => \N__43092\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__43092\,
            I => \N__43087\
        );

    \I__9540\ : InMux
    port map (
            O => \N__43091\,
            I => \N__43082\
        );

    \I__9539\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43082\
        );

    \I__9538\ : Span12Mux_h
    port map (
            O => \N__43087\,
            I => \N__43079\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__43082\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__9536\ : Odrv12
    port map (
            O => \N__43079\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__9535\ : CEMux
    port map (
            O => \N__43074\,
            I => \N__43071\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__43071\,
            I => \N__43056\
        );

    \I__9533\ : InMux
    port map (
            O => \N__43070\,
            I => \N__43053\
        );

    \I__9532\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43027\
        );

    \I__9531\ : InMux
    port map (
            O => \N__43068\,
            I => \N__43027\
        );

    \I__9530\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43027\
        );

    \I__9529\ : InMux
    port map (
            O => \N__43066\,
            I => \N__43027\
        );

    \I__9528\ : InMux
    port map (
            O => \N__43065\,
            I => \N__43027\
        );

    \I__9527\ : InMux
    port map (
            O => \N__43064\,
            I => \N__43027\
        );

    \I__9526\ : InMux
    port map (
            O => \N__43063\,
            I => \N__43027\
        );

    \I__9525\ : InMux
    port map (
            O => \N__43062\,
            I => \N__43027\
        );

    \I__9524\ : InMux
    port map (
            O => \N__43061\,
            I => \N__43024\
        );

    \I__9523\ : SRMux
    port map (
            O => \N__43060\,
            I => \N__43021\
        );

    \I__9522\ : CascadeMux
    port map (
            O => \N__43059\,
            I => \N__43017\
        );

    \I__9521\ : Span4Mux_v
    port map (
            O => \N__43056\,
            I => \N__43014\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__43053\,
            I => \N__43011\
        );

    \I__9519\ : InMux
    port map (
            O => \N__43052\,
            I => \N__43006\
        );

    \I__9518\ : InMux
    port map (
            O => \N__43051\,
            I => \N__43006\
        );

    \I__9517\ : InMux
    port map (
            O => \N__43050\,
            I => \N__42993\
        );

    \I__9516\ : InMux
    port map (
            O => \N__43049\,
            I => \N__42993\
        );

    \I__9515\ : InMux
    port map (
            O => \N__43048\,
            I => \N__42993\
        );

    \I__9514\ : InMux
    port map (
            O => \N__43047\,
            I => \N__42993\
        );

    \I__9513\ : InMux
    port map (
            O => \N__43046\,
            I => \N__42993\
        );

    \I__9512\ : InMux
    port map (
            O => \N__43045\,
            I => \N__42993\
        );

    \I__9511\ : InMux
    port map (
            O => \N__43044\,
            I => \N__42990\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__43027\,
            I => \N__42987\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__43024\,
            I => \N__42984\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__43021\,
            I => \N__42980\
        );

    \I__9507\ : InMux
    port map (
            O => \N__43020\,
            I => \N__42977\
        );

    \I__9506\ : InMux
    port map (
            O => \N__43017\,
            I => \N__42973\
        );

    \I__9505\ : Span4Mux_h
    port map (
            O => \N__43014\,
            I => \N__42968\
        );

    \I__9504\ : Span4Mux_h
    port map (
            O => \N__43011\,
            I => \N__42968\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__43006\,
            I => \N__42965\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__42993\,
            I => \N__42962\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42990\,
            I => \N__42959\
        );

    \I__9500\ : Span4Mux_v
    port map (
            O => \N__42987\,
            I => \N__42953\
        );

    \I__9499\ : Span4Mux_h
    port map (
            O => \N__42984\,
            I => \N__42950\
        );

    \I__9498\ : InMux
    port map (
            O => \N__42983\,
            I => \N__42947\
        );

    \I__9497\ : Span4Mux_h
    port map (
            O => \N__42980\,
            I => \N__42944\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__42977\,
            I => \N__42941\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42938\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42973\,
            I => \N__42933\
        );

    \I__9493\ : Span4Mux_v
    port map (
            O => \N__42968\,
            I => \N__42933\
        );

    \I__9492\ : Span4Mux_v
    port map (
            O => \N__42965\,
            I => \N__42930\
        );

    \I__9491\ : Span4Mux_v
    port map (
            O => \N__42962\,
            I => \N__42925\
        );

    \I__9490\ : Span4Mux_v
    port map (
            O => \N__42959\,
            I => \N__42925\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42918\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42918\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42956\,
            I => \N__42918\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__42953\,
            I => \N__42915\
        );

    \I__9485\ : Sp12to4
    port map (
            O => \N__42950\,
            I => \N__42912\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__42947\,
            I => \N__42905\
        );

    \I__9483\ : Span4Mux_h
    port map (
            O => \N__42944\,
            I => \N__42905\
        );

    \I__9482\ : Span4Mux_v
    port map (
            O => \N__42941\,
            I => \N__42905\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__42938\,
            I => \N__42900\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__42933\,
            I => \N__42900\
        );

    \I__9479\ : Odrv4
    port map (
            O => \N__42930\,
            I => dds_state_1
        );

    \I__9478\ : Odrv4
    port map (
            O => \N__42925\,
            I => dds_state_1
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__42918\,
            I => dds_state_1
        );

    \I__9476\ : Odrv4
    port map (
            O => \N__42915\,
            I => dds_state_1
        );

    \I__9475\ : Odrv12
    port map (
            O => \N__42912\,
            I => dds_state_1
        );

    \I__9474\ : Odrv4
    port map (
            O => \N__42905\,
            I => dds_state_1
        );

    \I__9473\ : Odrv4
    port map (
            O => \N__42900\,
            I => dds_state_1
        );

    \I__9472\ : SRMux
    port map (
            O => \N__42885\,
            I => \N__42882\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42882\,
            I => \N__42878\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42881\,
            I => \N__42875\
        );

    \I__9469\ : Span4Mux_v
    port map (
            O => \N__42878\,
            I => \N__42872\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__42875\,
            I => \N__42869\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__42872\,
            I => \N__42866\
        );

    \I__9466\ : Span4Mux_v
    port map (
            O => \N__42869\,
            I => \N__42863\
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__42866\,
            I => n14884
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__42863\,
            I => n14884
        );

    \I__9463\ : CEMux
    port map (
            O => \N__42858\,
            I => \N__42855\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42855\,
            I => n12220
        );

    \I__9461\ : CascadeMux
    port map (
            O => \N__42852\,
            I => \n12220_cascade_\
        );

    \I__9460\ : SRMux
    port map (
            O => \N__42849\,
            I => \N__42846\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__42846\,
            I => n14785
        );

    \I__9458\ : SRMux
    port map (
            O => \N__42843\,
            I => \N__42840\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__42840\,
            I => \N__42837\
        );

    \I__9456\ : Span4Mux_h
    port map (
            O => \N__42837\,
            I => \N__42834\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__42834\,
            I => n14778
        );

    \I__9454\ : InMux
    port map (
            O => \N__42831\,
            I => \N__42828\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__42828\,
            I => \N__42825\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__42825\,
            I => \N__42822\
        );

    \I__9451\ : Span4Mux_h
    port map (
            O => \N__42822\,
            I => \N__42819\
        );

    \I__9450\ : Odrv4
    port map (
            O => \N__42819\,
            I => n30_adj_1531
        );

    \I__9449\ : CascadeMux
    port map (
            O => \N__42816\,
            I => \N__42811\
        );

    \I__9448\ : CascadeMux
    port map (
            O => \N__42815\,
            I => \N__42807\
        );

    \I__9447\ : CascadeMux
    port map (
            O => \N__42814\,
            I => \N__42804\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42811\,
            I => \N__42799\
        );

    \I__9445\ : InMux
    port map (
            O => \N__42810\,
            I => \N__42794\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42807\,
            I => \N__42794\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42791\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42803\,
            I => \N__42788\
        );

    \I__9441\ : InMux
    port map (
            O => \N__42802\,
            I => \N__42785\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__42799\,
            I => \N__42782\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__42794\,
            I => \N__42777\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__42791\,
            I => \N__42777\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__42788\,
            I => \N__42774\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__42785\,
            I => \N__42771\
        );

    \I__9435\ : Span4Mux_h
    port map (
            O => \N__42782\,
            I => \N__42767\
        );

    \I__9434\ : Span4Mux_v
    port map (
            O => \N__42777\,
            I => \N__42762\
        );

    \I__9433\ : Span4Mux_v
    port map (
            O => \N__42774\,
            I => \N__42762\
        );

    \I__9432\ : Span4Mux_h
    port map (
            O => \N__42771\,
            I => \N__42759\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42770\,
            I => \N__42756\
        );

    \I__9430\ : Span4Mux_h
    port map (
            O => \N__42767\,
            I => \N__42753\
        );

    \I__9429\ : Span4Mux_h
    port map (
            O => \N__42762\,
            I => \N__42746\
        );

    \I__9428\ : Span4Mux_v
    port map (
            O => \N__42759\,
            I => \N__42746\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__42756\,
            I => \N__42746\
        );

    \I__9426\ : Span4Mux_v
    port map (
            O => \N__42753\,
            I => \N__42743\
        );

    \I__9425\ : Span4Mux_h
    port map (
            O => \N__42746\,
            I => \N__42740\
        );

    \I__9424\ : Odrv4
    port map (
            O => \N__42743\,
            I => comm_buf_0_7
        );

    \I__9423\ : Odrv4
    port map (
            O => \N__42740\,
            I => comm_buf_0_7
        );

    \I__9422\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42729\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42734\,
            I => \N__42729\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__42729\,
            I => \N__42725\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42728\,
            I => \N__42722\
        );

    \I__9418\ : Odrv12
    port map (
            O => \N__42725\,
            I => comm_tx_buf_5
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__42722\,
            I => comm_tx_buf_5
        );

    \I__9416\ : InMux
    port map (
            O => \N__42717\,
            I => \N__42714\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__42714\,
            I => \N__42711\
        );

    \I__9414\ : Span4Mux_h
    port map (
            O => \N__42711\,
            I => \N__42708\
        );

    \I__9413\ : Span4Mux_v
    port map (
            O => \N__42708\,
            I => \N__42705\
        );

    \I__9412\ : Span4Mux_v
    port map (
            O => \N__42705\,
            I => \N__42702\
        );

    \I__9411\ : Odrv4
    port map (
            O => \N__42702\,
            I => buf_data_vac_8
        );

    \I__9410\ : InMux
    port map (
            O => \N__42699\,
            I => \N__42696\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__42696\,
            I => \N__42693\
        );

    \I__9408\ : Odrv4
    port map (
            O => \N__42693\,
            I => comm_buf_4_0
        );

    \I__9407\ : InMux
    port map (
            O => \N__42690\,
            I => \N__42687\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__42687\,
            I => \N__42684\
        );

    \I__9405\ : Span4Mux_h
    port map (
            O => \N__42684\,
            I => \N__42681\
        );

    \I__9404\ : Span4Mux_h
    port map (
            O => \N__42681\,
            I => \N__42678\
        );

    \I__9403\ : Odrv4
    port map (
            O => \N__42678\,
            I => buf_data_vac_15
        );

    \I__9402\ : InMux
    port map (
            O => \N__42675\,
            I => \N__42672\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__42672\,
            I => \N__42669\
        );

    \I__9400\ : Span4Mux_v
    port map (
            O => \N__42669\,
            I => \N__42666\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__42663\,
            I => comm_buf_4_7
        );

    \I__9397\ : InMux
    port map (
            O => \N__42660\,
            I => \N__42657\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__42657\,
            I => \N__42654\
        );

    \I__9395\ : Span4Mux_v
    port map (
            O => \N__42654\,
            I => \N__42651\
        );

    \I__9394\ : Span4Mux_v
    port map (
            O => \N__42651\,
            I => \N__42648\
        );

    \I__9393\ : Odrv4
    port map (
            O => \N__42648\,
            I => buf_data_vac_14
        );

    \I__9392\ : InMux
    port map (
            O => \N__42645\,
            I => \N__42642\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42642\,
            I => \N__42639\
        );

    \I__9390\ : Odrv4
    port map (
            O => \N__42639\,
            I => comm_buf_4_6
        );

    \I__9389\ : InMux
    port map (
            O => \N__42636\,
            I => \N__42633\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__42633\,
            I => \N__42630\
        );

    \I__9387\ : Span4Mux_h
    port map (
            O => \N__42630\,
            I => \N__42627\
        );

    \I__9386\ : Span4Mux_v
    port map (
            O => \N__42627\,
            I => \N__42624\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__42624\,
            I => buf_data_vac_13
        );

    \I__9384\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42618\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42618\,
            I => comm_buf_4_5
        );

    \I__9382\ : InMux
    port map (
            O => \N__42615\,
            I => \N__42612\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__42612\,
            I => \N__42609\
        );

    \I__9380\ : Span12Mux_h
    port map (
            O => \N__42609\,
            I => \N__42606\
        );

    \I__9379\ : Odrv12
    port map (
            O => \N__42606\,
            I => buf_data_vac_12
        );

    \I__9378\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42600\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__42600\,
            I => \N__42597\
        );

    \I__9376\ : Span4Mux_h
    port map (
            O => \N__42597\,
            I => \N__42594\
        );

    \I__9375\ : Odrv4
    port map (
            O => \N__42594\,
            I => comm_buf_4_4
        );

    \I__9374\ : InMux
    port map (
            O => \N__42591\,
            I => \N__42588\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__42588\,
            I => \N__42585\
        );

    \I__9372\ : Span4Mux_h
    port map (
            O => \N__42585\,
            I => \N__42582\
        );

    \I__9371\ : Span4Mux_v
    port map (
            O => \N__42582\,
            I => \N__42579\
        );

    \I__9370\ : Odrv4
    port map (
            O => \N__42579\,
            I => buf_data_vac_11
        );

    \I__9369\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42573\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__42573\,
            I => \N__42570\
        );

    \I__9367\ : Span4Mux_h
    port map (
            O => \N__42570\,
            I => \N__42567\
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__42567\,
            I => comm_buf_4_3
        );

    \I__9365\ : InMux
    port map (
            O => \N__42564\,
            I => \N__42561\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__42561\,
            I => \N__42558\
        );

    \I__9363\ : Span4Mux_h
    port map (
            O => \N__42558\,
            I => \N__42555\
        );

    \I__9362\ : Span4Mux_v
    port map (
            O => \N__42555\,
            I => \N__42552\
        );

    \I__9361\ : Span4Mux_v
    port map (
            O => \N__42552\,
            I => \N__42549\
        );

    \I__9360\ : Odrv4
    port map (
            O => \N__42549\,
            I => buf_data_vac_10
        );

    \I__9359\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__42543\,
            I => comm_buf_4_2
        );

    \I__9357\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42537\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__42537\,
            I => \N__42534\
        );

    \I__9355\ : Span4Mux_v
    port map (
            O => \N__42534\,
            I => \N__42531\
        );

    \I__9354\ : Span4Mux_h
    port map (
            O => \N__42531\,
            I => \N__42528\
        );

    \I__9353\ : Span4Mux_v
    port map (
            O => \N__42528\,
            I => \N__42525\
        );

    \I__9352\ : Odrv4
    port map (
            O => \N__42525\,
            I => buf_data_vac_9
        );

    \I__9351\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42519\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__42519\,
            I => \N__42516\
        );

    \I__9349\ : Odrv4
    port map (
            O => \N__42516\,
            I => n1
        );

    \I__9348\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42510\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__42510\,
            I => \N__42507\
        );

    \I__9346\ : Span4Mux_h
    port map (
            O => \N__42507\,
            I => \N__42504\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__42504\,
            I => comm_buf_2_0
        );

    \I__9344\ : InMux
    port map (
            O => \N__42501\,
            I => \N__42498\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__42498\,
            I => n2
        );

    \I__9342\ : InMux
    port map (
            O => \N__42495\,
            I => \N__42491\
        );

    \I__9341\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42488\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__42491\,
            I => \N__42485\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__42488\,
            I => \N__42482\
        );

    \I__9338\ : Span4Mux_h
    port map (
            O => \N__42485\,
            I => \N__42478\
        );

    \I__9337\ : Span4Mux_v
    port map (
            O => \N__42482\,
            I => \N__42475\
        );

    \I__9336\ : InMux
    port map (
            O => \N__42481\,
            I => \N__42472\
        );

    \I__9335\ : Odrv4
    port map (
            O => \N__42478\,
            I => comm_tx_buf_0
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__42475\,
            I => comm_tx_buf_0
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__42472\,
            I => comm_tx_buf_0
        );

    \I__9332\ : SRMux
    port map (
            O => \N__42465\,
            I => \N__42462\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__42462\,
            I => \N__42459\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__42459\,
            I => \N__42456\
        );

    \I__9329\ : Span4Mux_v
    port map (
            O => \N__42456\,
            I => \N__42453\
        );

    \I__9328\ : Odrv4
    port map (
            O => \N__42453\,
            I => \comm_spi.data_tx_7__N_773\
        );

    \I__9327\ : CascadeMux
    port map (
            O => \N__42450\,
            I => \n17479_cascade_\
        );

    \I__9326\ : InMux
    port map (
            O => \N__42447\,
            I => \N__42443\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42446\,
            I => \N__42440\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__42443\,
            I => \N__42437\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__42440\,
            I => \N__42432\
        );

    \I__9322\ : Span4Mux_v
    port map (
            O => \N__42437\,
            I => \N__42432\
        );

    \I__9321\ : Odrv4
    port map (
            O => \N__42432\,
            I => comm_buf_6_5
        );

    \I__9320\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42426\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__42426\,
            I => \N__42423\
        );

    \I__9318\ : Span4Mux_h
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__9317\ : Odrv4
    port map (
            O => \N__42420\,
            I => comm_buf_2_5
        );

    \I__9316\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42414\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__42414\,
            I => \N__42411\
        );

    \I__9314\ : Odrv4
    port map (
            O => \N__42411\,
            I => n17480
        );

    \I__9313\ : InMux
    port map (
            O => \N__42408\,
            I => \N__42405\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42405\,
            I => comm_buf_5_5
        );

    \I__9311\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42399\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__42399\,
            I => n21212
        );

    \I__9309\ : CascadeMux
    port map (
            O => \N__42396\,
            I => \n17482_cascade_\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42393\,
            I => \N__42390\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__42390\,
            I => n22189
        );

    \I__9306\ : InMux
    port map (
            O => \N__42387\,
            I => \N__42383\
        );

    \I__9305\ : InMux
    port map (
            O => \N__42386\,
            I => \N__42380\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__42383\,
            I => \N__42375\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__42380\,
            I => \N__42375\
        );

    \I__9302\ : Odrv12
    port map (
            O => \N__42375\,
            I => \comm_spi.n14639\
        );

    \I__9301\ : SRMux
    port map (
            O => \N__42372\,
            I => \N__42369\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__42369\,
            I => \N__42366\
        );

    \I__9299\ : Span4Mux_h
    port map (
            O => \N__42366\,
            I => \N__42363\
        );

    \I__9298\ : Odrv4
    port map (
            O => \N__42363\,
            I => \comm_spi.data_tx_7__N_777\
        );

    \I__9297\ : SRMux
    port map (
            O => \N__42360\,
            I => \N__42357\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__42357\,
            I => \N__42354\
        );

    \I__9295\ : Span4Mux_v
    port map (
            O => \N__42354\,
            I => \N__42351\
        );

    \I__9294\ : Odrv4
    port map (
            O => \N__42351\,
            I => \comm_spi.data_tx_7__N_780\
        );

    \I__9293\ : InMux
    port map (
            O => \N__42348\,
            I => \N__42345\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9291\ : Odrv4
    port map (
            O => \N__42342\,
            I => comm_buf_5_6
        );

    \I__9290\ : CascadeMux
    port map (
            O => \N__42339\,
            I => \n22183_cascade_\
        );

    \I__9289\ : InMux
    port map (
            O => \N__42336\,
            I => \N__42333\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__42333\,
            I => \N__42330\
        );

    \I__9287\ : Span4Mux_h
    port map (
            O => \N__42330\,
            I => \N__42327\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__42327\,
            I => comm_buf_5_0
        );

    \I__9285\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42321\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__42321\,
            I => n4
        );

    \I__9283\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42314\
        );

    \I__9282\ : CascadeMux
    port map (
            O => \N__42317\,
            I => \N__42311\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42314\,
            I => \N__42308\
        );

    \I__9280\ : InMux
    port map (
            O => \N__42311\,
            I => \N__42305\
        );

    \I__9279\ : Span4Mux_v
    port map (
            O => \N__42308\,
            I => \N__42302\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__42305\,
            I => comm_buf_6_0
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__42302\,
            I => comm_buf_6_0
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__9275\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42291\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__42291\,
            I => n21211
        );

    \I__9273\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42279\
        );

    \I__9272\ : CascadeMux
    port map (
            O => \N__42287\,
            I => \N__42276\
        );

    \I__9271\ : InMux
    port map (
            O => \N__42286\,
            I => \N__42263\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__42285\,
            I => \N__42259\
        );

    \I__9269\ : CascadeMux
    port map (
            O => \N__42284\,
            I => \N__42256\
        );

    \I__9268\ : CascadeMux
    port map (
            O => \N__42283\,
            I => \N__42253\
        );

    \I__9267\ : CascadeMux
    port map (
            O => \N__42282\,
            I => \N__42250\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__42279\,
            I => \N__42245\
        );

    \I__9265\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42242\
        );

    \I__9264\ : InMux
    port map (
            O => \N__42275\,
            I => \N__42225\
        );

    \I__9263\ : InMux
    port map (
            O => \N__42274\,
            I => \N__42225\
        );

    \I__9262\ : InMux
    port map (
            O => \N__42273\,
            I => \N__42225\
        );

    \I__9261\ : InMux
    port map (
            O => \N__42272\,
            I => \N__42225\
        );

    \I__9260\ : InMux
    port map (
            O => \N__42271\,
            I => \N__42225\
        );

    \I__9259\ : InMux
    port map (
            O => \N__42270\,
            I => \N__42225\
        );

    \I__9258\ : InMux
    port map (
            O => \N__42269\,
            I => \N__42225\
        );

    \I__9257\ : InMux
    port map (
            O => \N__42268\,
            I => \N__42225\
        );

    \I__9256\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42222\
        );

    \I__9255\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42219\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__42263\,
            I => \N__42216\
        );

    \I__9253\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42201\
        );

    \I__9252\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42201\
        );

    \I__9251\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42201\
        );

    \I__9250\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42201\
        );

    \I__9249\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42201\
        );

    \I__9248\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42201\
        );

    \I__9247\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42201\
        );

    \I__9246\ : Span4Mux_h
    port map (
            O => \N__42245\,
            I => \N__42198\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__42242\,
            I => \N__42191\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__42225\,
            I => \N__42191\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__42222\,
            I => \N__42185\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__42219\,
            I => \N__42182\
        );

    \I__9241\ : Span4Mux_v
    port map (
            O => \N__42216\,
            I => \N__42179\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__42201\,
            I => \N__42174\
        );

    \I__9239\ : Span4Mux_v
    port map (
            O => \N__42198\,
            I => \N__42174\
        );

    \I__9238\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42171\
        );

    \I__9237\ : InMux
    port map (
            O => \N__42196\,
            I => \N__42168\
        );

    \I__9236\ : Span4Mux_h
    port map (
            O => \N__42191\,
            I => \N__42165\
        );

    \I__9235\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42158\
        );

    \I__9234\ : InMux
    port map (
            O => \N__42189\,
            I => \N__42158\
        );

    \I__9233\ : InMux
    port map (
            O => \N__42188\,
            I => \N__42158\
        );

    \I__9232\ : Span4Mux_h
    port map (
            O => \N__42185\,
            I => \N__42153\
        );

    \I__9231\ : Span4Mux_v
    port map (
            O => \N__42182\,
            I => \N__42153\
        );

    \I__9230\ : Span4Mux_v
    port map (
            O => \N__42179\,
            I => \N__42150\
        );

    \I__9229\ : Span4Mux_v
    port map (
            O => \N__42174\,
            I => \N__42147\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__42171\,
            I => dds_state_2
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__42168\,
            I => dds_state_2
        );

    \I__9226\ : Odrv4
    port map (
            O => \N__42165\,
            I => dds_state_2
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__42158\,
            I => dds_state_2
        );

    \I__9224\ : Odrv4
    port map (
            O => \N__42153\,
            I => dds_state_2
        );

    \I__9223\ : Odrv4
    port map (
            O => \N__42150\,
            I => dds_state_2
        );

    \I__9222\ : Odrv4
    port map (
            O => \N__42147\,
            I => dds_state_2
        );

    \I__9221\ : CascadeMux
    port map (
            O => \N__42132\,
            I => \N__42128\
        );

    \I__9220\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42125\
        );

    \I__9219\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42121\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__42125\,
            I => \N__42117\
        );

    \I__9217\ : InMux
    port map (
            O => \N__42124\,
            I => \N__42114\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__42121\,
            I => \N__42111\
        );

    \I__9215\ : CascadeMux
    port map (
            O => \N__42120\,
            I => \N__42108\
        );

    \I__9214\ : Span4Mux_v
    port map (
            O => \N__42117\,
            I => \N__42105\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__42114\,
            I => \N__42100\
        );

    \I__9212\ : Span4Mux_h
    port map (
            O => \N__42111\,
            I => \N__42100\
        );

    \I__9211\ : InMux
    port map (
            O => \N__42108\,
            I => \N__42097\
        );

    \I__9210\ : Odrv4
    port map (
            O => \N__42105\,
            I => trig_dds0
        );

    \I__9209\ : Odrv4
    port map (
            O => \N__42100\,
            I => trig_dds0
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__42097\,
            I => trig_dds0
        );

    \I__9207\ : CEMux
    port map (
            O => \N__42090\,
            I => \N__42086\
        );

    \I__9206\ : CEMux
    port map (
            O => \N__42089\,
            I => \N__42083\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__42086\,
            I => \N__42080\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__42083\,
            I => \N__42077\
        );

    \I__9203\ : Span4Mux_h
    port map (
            O => \N__42080\,
            I => \N__42074\
        );

    \I__9202\ : Span4Mux_h
    port map (
            O => \N__42077\,
            I => \N__42071\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__42074\,
            I => \N__42068\
        );

    \I__9200\ : Odrv4
    port map (
            O => \N__42071\,
            I => \SIG_DDS.n12722\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__42068\,
            I => \SIG_DDS.n12722\
        );

    \I__9198\ : InMux
    port map (
            O => \N__42063\,
            I => \N__42059\
        );

    \I__9197\ : InMux
    port map (
            O => \N__42062\,
            I => \N__42055\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__42059\,
            I => \N__42052\
        );

    \I__9195\ : InMux
    port map (
            O => \N__42058\,
            I => \N__42049\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__42055\,
            I => data_index_8
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__42052\,
            I => data_index_8
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__42049\,
            I => data_index_8
        );

    \I__9191\ : InMux
    port map (
            O => \N__42042\,
            I => \N__42039\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__42036\
        );

    \I__9189\ : Span4Mux_h
    port map (
            O => \N__42036\,
            I => \N__42032\
        );

    \I__9188\ : InMux
    port map (
            O => \N__42035\,
            I => \N__42029\
        );

    \I__9187\ : Odrv4
    port map (
            O => \N__42032\,
            I => n8_adj_1561
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__42029\,
            I => n8_adj_1561
        );

    \I__9185\ : InMux
    port map (
            O => \N__42024\,
            I => \N__42020\
        );

    \I__9184\ : InMux
    port map (
            O => \N__42023\,
            I => \N__42017\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__42020\,
            I => n8_adj_1563
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__42017\,
            I => n8_adj_1563
        );

    \I__9181\ : CascadeMux
    port map (
            O => \N__42012\,
            I => \N__42009\
        );

    \I__9180\ : InMux
    port map (
            O => \N__42009\,
            I => \N__42006\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__42006\,
            I => \N__42003\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__42003\,
            I => \N__41999\
        );

    \I__9177\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41996\
        );

    \I__9176\ : Odrv4
    port map (
            O => \N__41999\,
            I => n7_adj_1562
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__41996\,
            I => n7_adj_1562
        );

    \I__9174\ : InMux
    port map (
            O => \N__41991\,
            I => \N__41987\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41984\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__41987\,
            I => \N__41979\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__41984\,
            I => \N__41979\
        );

    \I__9170\ : Span4Mux_h
    port map (
            O => \N__41979\,
            I => \N__41975\
        );

    \I__9169\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41972\
        );

    \I__9168\ : Span4Mux_h
    port map (
            O => \N__41975\,
            I => \N__41969\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__41972\,
            I => data_index_7
        );

    \I__9166\ : Odrv4
    port map (
            O => \N__41969\,
            I => data_index_7
        );

    \I__9165\ : IoInMux
    port map (
            O => \N__41964\,
            I => \N__41961\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__9163\ : IoSpan4Mux
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__9162\ : Span4Mux_s3_v
    port map (
            O => \N__41955\,
            I => \N__41950\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41954\,
            I => \N__41947\
        );

    \I__9160\ : InMux
    port map (
            O => \N__41953\,
            I => \N__41944\
        );

    \I__9159\ : Span4Mux_v
    port map (
            O => \N__41950\,
            I => \N__41939\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41947\,
            I => \N__41939\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41944\,
            I => \SELIRNG1\
        );

    \I__9156\ : Odrv4
    port map (
            O => \N__41939\,
            I => \SELIRNG1\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41934\,
            I => \N__41931\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41931\,
            I => \N__41928\
        );

    \I__9153\ : Span4Mux_h
    port map (
            O => \N__41928\,
            I => \N__41923\
        );

    \I__9152\ : CascadeMux
    port map (
            O => \N__41927\,
            I => \N__41920\
        );

    \I__9151\ : InMux
    port map (
            O => \N__41926\,
            I => \N__41917\
        );

    \I__9150\ : Span4Mux_h
    port map (
            O => \N__41923\,
            I => \N__41914\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41920\,
            I => \N__41911\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__41917\,
            I => \acadc_skipCount_11\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__41914\,
            I => \acadc_skipCount_11\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41911\,
            I => \acadc_skipCount_11\
        );

    \I__9145\ : CascadeMux
    port map (
            O => \N__41904\,
            I => \N__41901\
        );

    \I__9144\ : InMux
    port map (
            O => \N__41901\,
            I => \N__41898\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__41898\,
            I => \N__41895\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__41895\,
            I => n23_adj_1543
        );

    \I__9141\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41888\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41883\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__41888\,
            I => \N__41880\
        );

    \I__9138\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41875\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41875\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41871\
        );

    \I__9135\ : Span4Mux_h
    port map (
            O => \N__41880\,
            I => \N__41866\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__41875\,
            I => \N__41866\
        );

    \I__9133\ : InMux
    port map (
            O => \N__41874\,
            I => \N__41863\
        );

    \I__9132\ : Span12Mux_h
    port map (
            O => \N__41871\,
            I => \N__41858\
        );

    \I__9131\ : Span4Mux_h
    port map (
            O => \N__41866\,
            I => \N__41853\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__41863\,
            I => \N__41853\
        );

    \I__9129\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41850\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41847\
        );

    \I__9127\ : Odrv12
    port map (
            O => \N__41858\,
            I => n11915
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__41853\,
            I => n11915
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__41850\,
            I => n11915
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__41847\,
            I => n11915
        );

    \I__9123\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41835\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41835\,
            I => \N__41832\
        );

    \I__9121\ : Odrv12
    port map (
            O => \N__41832\,
            I => buf_data_iac_22
        );

    \I__9120\ : InMux
    port map (
            O => \N__41829\,
            I => \N__41826\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__41826\,
            I => \N__41823\
        );

    \I__9118\ : Span12Mux_h
    port map (
            O => \N__41823\,
            I => \N__41820\
        );

    \I__9117\ : Odrv12
    port map (
            O => \N__41820\,
            I => n21273
        );

    \I__9116\ : InMux
    port map (
            O => \N__41817\,
            I => \N__41814\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__41814\,
            I => \N__41811\
        );

    \I__9114\ : Span4Mux_h
    port map (
            O => \N__41811\,
            I => \N__41808\
        );

    \I__9113\ : Odrv4
    port map (
            O => \N__41808\,
            I => buf_data_iac_20
        );

    \I__9112\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41802\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__41802\,
            I => \N__41799\
        );

    \I__9110\ : Span4Mux_v
    port map (
            O => \N__41799\,
            I => \N__41796\
        );

    \I__9109\ : Span4Mux_v
    port map (
            O => \N__41796\,
            I => \N__41793\
        );

    \I__9108\ : Odrv4
    port map (
            O => \N__41793\,
            I => n21569
        );

    \I__9107\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41786\
        );

    \I__9106\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41783\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__41786\,
            I => \comm_spi.n14592\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__41783\,
            I => \comm_spi.n14592\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41778\,
            I => \N__41774\
        );

    \I__9102\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41771\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__41774\,
            I => \N__41768\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__41771\,
            I => \N__41765\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__41768\,
            I => \N__41757\
        );

    \I__9098\ : Span4Mux_v
    port map (
            O => \N__41765\,
            I => \N__41757\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41754\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41749\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41762\,
            I => \N__41749\
        );

    \I__9094\ : Odrv4
    port map (
            O => \N__41757\,
            I => n20907
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__41754\,
            I => n20907
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__41749\,
            I => n20907
        );

    \I__9091\ : InMux
    port map (
            O => \N__41742\,
            I => \N__41736\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41741\,
            I => \N__41731\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41740\,
            I => \N__41731\
        );

    \I__9088\ : CascadeMux
    port map (
            O => \N__41739\,
            I => \N__41726\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__41736\,
            I => \N__41718\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__41731\,
            I => \N__41718\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41730\,
            I => \N__41713\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41729\,
            I => \N__41713\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41726\,
            I => \N__41708\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41725\,
            I => \N__41708\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__41724\,
            I => \N__41705\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41695\
        );

    \I__9079\ : Span4Mux_v
    port map (
            O => \N__41718\,
            I => \N__41688\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41713\,
            I => \N__41688\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__41708\,
            I => \N__41688\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41679\
        );

    \I__9075\ : InMux
    port map (
            O => \N__41704\,
            I => \N__41679\
        );

    \I__9074\ : InMux
    port map (
            O => \N__41703\,
            I => \N__41679\
        );

    \I__9073\ : InMux
    port map (
            O => \N__41702\,
            I => \N__41679\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41701\,
            I => \N__41672\
        );

    \I__9071\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41672\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41699\,
            I => \N__41672\
        );

    \I__9069\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41669\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__41695\,
            I => \N__41666\
        );

    \I__9067\ : Span4Mux_h
    port map (
            O => \N__41688\,
            I => \N__41663\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__41679\,
            I => \N__41660\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__41672\,
            I => \N__41655\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__41669\,
            I => \N__41655\
        );

    \I__9063\ : Span4Mux_v
    port map (
            O => \N__41666\,
            I => \N__41652\
        );

    \I__9062\ : Span4Mux_h
    port map (
            O => \N__41663\,
            I => \N__41649\
        );

    \I__9061\ : Span4Mux_h
    port map (
            O => \N__41660\,
            I => \N__41646\
        );

    \I__9060\ : Span4Mux_h
    port map (
            O => \N__41655\,
            I => \N__41643\
        );

    \I__9059\ : Odrv4
    port map (
            O => \N__41652\,
            I => n12429
        );

    \I__9058\ : Odrv4
    port map (
            O => \N__41649\,
            I => n12429
        );

    \I__9057\ : Odrv4
    port map (
            O => \N__41646\,
            I => n12429
        );

    \I__9056\ : Odrv4
    port map (
            O => \N__41643\,
            I => n12429
        );

    \I__9055\ : CascadeMux
    port map (
            O => \N__41634\,
            I => \n9306_cascade_\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41631\,
            I => \N__41627\
        );

    \I__9053\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41624\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41627\,
            I => \N__41621\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__41624\,
            I => \N__41618\
        );

    \I__9050\ : Span4Mux_v
    port map (
            O => \N__41621\,
            I => \N__41612\
        );

    \I__9049\ : Span4Mux_h
    port map (
            O => \N__41618\,
            I => \N__41612\
        );

    \I__9048\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41609\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__41612\,
            I => \N__41606\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__41609\,
            I => buf_dds0_13
        );

    \I__9045\ : Odrv4
    port map (
            O => \N__41606\,
            I => buf_dds0_13
        );

    \I__9044\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41598\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__41598\,
            I => \N__41594\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41591\
        );

    \I__9041\ : Span4Mux_h
    port map (
            O => \N__41594\,
            I => \N__41588\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__41591\,
            I => acadc_skipcnt_7
        );

    \I__9039\ : Odrv4
    port map (
            O => \N__41588\,
            I => acadc_skipcnt_7
        );

    \I__9038\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41580\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41580\,
            I => \N__41576\
        );

    \I__9036\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41573\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__41576\,
            I => \N__41570\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__41573\,
            I => acadc_skipcnt_2
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__41570\,
            I => acadc_skipcnt_2
        );

    \I__9032\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41562\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41562\,
            I => \N__41559\
        );

    \I__9030\ : Span4Mux_h
    port map (
            O => \N__41559\,
            I => \N__41556\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__41556\,
            I => n22
        );

    \I__9028\ : InMux
    port map (
            O => \N__41553\,
            I => \N__41549\
        );

    \I__9027\ : InMux
    port map (
            O => \N__41552\,
            I => \N__41546\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__41549\,
            I => n9
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__41546\,
            I => n9
        );

    \I__9024\ : CascadeMux
    port map (
            O => \N__41541\,
            I => \N__41537\
        );

    \I__9023\ : CascadeMux
    port map (
            O => \N__41540\,
            I => \N__41534\
        );

    \I__9022\ : InMux
    port map (
            O => \N__41537\,
            I => \N__41529\
        );

    \I__9021\ : InMux
    port map (
            O => \N__41534\,
            I => \N__41526\
        );

    \I__9020\ : InMux
    port map (
            O => \N__41533\,
            I => \N__41523\
        );

    \I__9019\ : CascadeMux
    port map (
            O => \N__41532\,
            I => \N__41520\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__41529\,
            I => \N__41517\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__41526\,
            I => \N__41514\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__41523\,
            I => \N__41511\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41508\
        );

    \I__9014\ : Span4Mux_v
    port map (
            O => \N__41517\,
            I => \N__41503\
        );

    \I__9013\ : Span4Mux_v
    port map (
            O => \N__41514\,
            I => \N__41503\
        );

    \I__9012\ : Odrv12
    port map (
            O => \N__41511\,
            I => n20912
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__41508\,
            I => n20912
        );

    \I__9010\ : Odrv4
    port map (
            O => \N__41503\,
            I => n20912
        );

    \I__9009\ : CascadeMux
    port map (
            O => \N__41496\,
            I => \N__41488\
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__41495\,
            I => \N__41485\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41481\
        );

    \I__9006\ : CascadeMux
    port map (
            O => \N__41493\,
            I => \N__41478\
        );

    \I__9005\ : CascadeMux
    port map (
            O => \N__41492\,
            I => \N__41475\
        );

    \I__9004\ : CascadeMux
    port map (
            O => \N__41491\,
            I => \N__41472\
        );

    \I__9003\ : InMux
    port map (
            O => \N__41488\,
            I => \N__41469\
        );

    \I__9002\ : InMux
    port map (
            O => \N__41485\,
            I => \N__41466\
        );

    \I__9001\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41462\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41481\,
            I => \N__41459\
        );

    \I__8999\ : InMux
    port map (
            O => \N__41478\,
            I => \N__41456\
        );

    \I__8998\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41453\
        );

    \I__8997\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41450\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__41469\,
            I => \N__41447\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__41466\,
            I => \N__41444\
        );

    \I__8994\ : InMux
    port map (
            O => \N__41465\,
            I => \N__41441\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__41462\,
            I => \N__41438\
        );

    \I__8992\ : Span4Mux_v
    port map (
            O => \N__41459\,
            I => \N__41433\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__41456\,
            I => \N__41433\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__41453\,
            I => \N__41428\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__41450\,
            I => \N__41428\
        );

    \I__8988\ : Span12Mux_h
    port map (
            O => \N__41447\,
            I => \N__41425\
        );

    \I__8987\ : Span4Mux_v
    port map (
            O => \N__41444\,
            I => \N__41422\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__41441\,
            I => \N__41417\
        );

    \I__8985\ : Sp12to4
    port map (
            O => \N__41438\,
            I => \N__41417\
        );

    \I__8984\ : Span4Mux_h
    port map (
            O => \N__41433\,
            I => \N__41412\
        );

    \I__8983\ : Span4Mux_v
    port map (
            O => \N__41428\,
            I => \N__41412\
        );

    \I__8982\ : Odrv12
    port map (
            O => \N__41425\,
            I => comm_buf_0_4
        );

    \I__8981\ : Odrv4
    port map (
            O => \N__41422\,
            I => comm_buf_0_4
        );

    \I__8980\ : Odrv12
    port map (
            O => \N__41417\,
            I => comm_buf_0_4
        );

    \I__8979\ : Odrv4
    port map (
            O => \N__41412\,
            I => comm_buf_0_4
        );

    \I__8978\ : CascadeMux
    port map (
            O => \N__41403\,
            I => \n12381_cascade_\
        );

    \I__8977\ : IoInMux
    port map (
            O => \N__41400\,
            I => \N__41397\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__41397\,
            I => \N__41394\
        );

    \I__8975\ : Span4Mux_s3_h
    port map (
            O => \N__41394\,
            I => \N__41391\
        );

    \I__8974\ : Span4Mux_h
    port map (
            O => \N__41391\,
            I => \N__41388\
        );

    \I__8973\ : Sp12to4
    port map (
            O => \N__41388\,
            I => \N__41384\
        );

    \I__8972\ : InMux
    port map (
            O => \N__41387\,
            I => \N__41381\
        );

    \I__8971\ : Span12Mux_s11_v
    port map (
            O => \N__41384\,
            I => \N__41378\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__41381\,
            I => \N__41374\
        );

    \I__8969\ : Span12Mux_h
    port map (
            O => \N__41378\,
            I => \N__41371\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41377\,
            I => \N__41368\
        );

    \I__8967\ : Span4Mux_v
    port map (
            O => \N__41374\,
            I => \N__41365\
        );

    \I__8966\ : Odrv12
    port map (
            O => \N__41371\,
            I => \VAC_OSR0\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__41368\,
            I => \VAC_OSR0\
        );

    \I__8964\ : Odrv4
    port map (
            O => \N__41365\,
            I => \VAC_OSR0\
        );

    \I__8963\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41354\
        );

    \I__8962\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41351\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__41354\,
            I => \N__41345\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__41351\,
            I => \N__41345\
        );

    \I__8959\ : InMux
    port map (
            O => \N__41350\,
            I => \N__41342\
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__41345\,
            I => \acadc_skipCount_6\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__41342\,
            I => \acadc_skipCount_6\
        );

    \I__8956\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41331\
        );

    \I__8955\ : CascadeMux
    port map (
            O => \N__41336\,
            I => \N__41328\
        );

    \I__8954\ : InMux
    port map (
            O => \N__41335\,
            I => \N__41324\
        );

    \I__8953\ : InMux
    port map (
            O => \N__41334\,
            I => \N__41320\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__41331\,
            I => \N__41317\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41328\,
            I => \N__41312\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41327\,
            I => \N__41312\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__41324\,
            I => \N__41308\
        );

    \I__8948\ : InMux
    port map (
            O => \N__41323\,
            I => \N__41305\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__41320\,
            I => \N__41302\
        );

    \I__8946\ : Span4Mux_v
    port map (
            O => \N__41317\,
            I => \N__41296\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__41312\,
            I => \N__41296\
        );

    \I__8944\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41293\
        );

    \I__8943\ : Span4Mux_h
    port map (
            O => \N__41308\,
            I => \N__41288\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__41305\,
            I => \N__41288\
        );

    \I__8941\ : Span4Mux_v
    port map (
            O => \N__41302\,
            I => \N__41285\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41301\,
            I => \N__41281\
        );

    \I__8939\ : Span4Mux_v
    port map (
            O => \N__41296\,
            I => \N__41276\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__41293\,
            I => \N__41276\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__41288\,
            I => \N__41273\
        );

    \I__8936\ : Sp12to4
    port map (
            O => \N__41285\,
            I => \N__41270\
        );

    \I__8935\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41267\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41264\
        );

    \I__8933\ : Span4Mux_h
    port map (
            O => \N__41276\,
            I => \N__41261\
        );

    \I__8932\ : Span4Mux_h
    port map (
            O => \N__41273\,
            I => \N__41258\
        );

    \I__8931\ : Span12Mux_h
    port map (
            O => \N__41270\,
            I => \N__41255\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__41267\,
            I => dds_state_0
        );

    \I__8929\ : Odrv12
    port map (
            O => \N__41264\,
            I => dds_state_0
        );

    \I__8928\ : Odrv4
    port map (
            O => \N__41261\,
            I => dds_state_0
        );

    \I__8927\ : Odrv4
    port map (
            O => \N__41258\,
            I => dds_state_0
        );

    \I__8926\ : Odrv12
    port map (
            O => \N__41255\,
            I => dds_state_0
        );

    \I__8925\ : CascadeMux
    port map (
            O => \N__41244\,
            I => \N__41241\
        );

    \I__8924\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41237\
        );

    \I__8923\ : InMux
    port map (
            O => \N__41240\,
            I => \N__41234\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__41237\,
            I => data_idxvec_10
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__41234\,
            I => data_idxvec_10
        );

    \I__8920\ : InMux
    port map (
            O => \N__41229\,
            I => \N__41226\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__41226\,
            I => \N__41222\
        );

    \I__8918\ : InMux
    port map (
            O => \N__41225\,
            I => \N__41218\
        );

    \I__8917\ : Span4Mux_h
    port map (
            O => \N__41222\,
            I => \N__41215\
        );

    \I__8916\ : InMux
    port map (
            O => \N__41221\,
            I => \N__41212\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__41218\,
            I => data_cntvec_10
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__41215\,
            I => data_cntvec_10
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__41212\,
            I => data_cntvec_10
        );

    \I__8912\ : InMux
    port map (
            O => \N__41205\,
            I => \N__41202\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__41202\,
            I => \N__41199\
        );

    \I__8910\ : Odrv4
    port map (
            O => \N__41199\,
            I => n21150
        );

    \I__8909\ : CascadeMux
    port map (
            O => \N__41196\,
            I => \N__41192\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__41195\,
            I => \N__41189\
        );

    \I__8907\ : InMux
    port map (
            O => \N__41192\,
            I => \N__41186\
        );

    \I__8906\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41183\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__41186\,
            I => \N__41180\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__41183\,
            I => data_idxvec_9
        );

    \I__8903\ : Odrv4
    port map (
            O => \N__41180\,
            I => data_idxvec_9
        );

    \I__8902\ : InMux
    port map (
            O => \N__41175\,
            I => \N__41172\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__41172\,
            I => \N__41168\
        );

    \I__8900\ : InMux
    port map (
            O => \N__41171\,
            I => \N__41164\
        );

    \I__8899\ : Span4Mux_v
    port map (
            O => \N__41168\,
            I => \N__41161\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41158\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__41164\,
            I => data_cntvec_9
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__41161\,
            I => data_cntvec_9
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__41158\,
            I => data_cntvec_9
        );

    \I__8894\ : InMux
    port map (
            O => \N__41151\,
            I => \N__41148\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41148\,
            I => \N__41145\
        );

    \I__8892\ : Odrv12
    port map (
            O => \N__41145\,
            I => n21060
        );

    \I__8891\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41139\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__41139\,
            I => \N__41136\
        );

    \I__8889\ : Span4Mux_h
    port map (
            O => \N__41136\,
            I => \N__41132\
        );

    \I__8888\ : InMux
    port map (
            O => \N__41135\,
            I => \N__41129\
        );

    \I__8887\ : Odrv4
    port map (
            O => \N__41132\,
            I => n8_adj_1569
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__41129\,
            I => n8_adj_1569
        );

    \I__8885\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41120\
        );

    \I__8884\ : CascadeMux
    port map (
            O => \N__41123\,
            I => \N__41117\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__41120\,
            I => \N__41114\
        );

    \I__8882\ : InMux
    port map (
            O => \N__41117\,
            I => \N__41111\
        );

    \I__8881\ : Span4Mux_v
    port map (
            O => \N__41114\,
            I => \N__41108\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__41111\,
            I => \N__41105\
        );

    \I__8879\ : Odrv4
    port map (
            O => \N__41108\,
            I => n7_adj_1568
        );

    \I__8878\ : Odrv4
    port map (
            O => \N__41105\,
            I => n7_adj_1568
        );

    \I__8877\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41095\
        );

    \I__8876\ : InMux
    port map (
            O => \N__41099\,
            I => \N__41092\
        );

    \I__8875\ : InMux
    port map (
            O => \N__41098\,
            I => \N__41089\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__41095\,
            I => \N__41084\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__41092\,
            I => \N__41084\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__41089\,
            I => \N__41081\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__41084\,
            I => \N__41078\
        );

    \I__8870\ : Span4Mux_h
    port map (
            O => \N__41081\,
            I => \N__41075\
        );

    \I__8869\ : Odrv4
    port map (
            O => \N__41078\,
            I => data_index_3
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__41075\,
            I => data_index_3
        );

    \I__8867\ : InMux
    port map (
            O => \N__41070\,
            I => \N__41066\
        );

    \I__8866\ : CascadeMux
    port map (
            O => \N__41069\,
            I => \N__41063\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__41066\,
            I => \N__41060\
        );

    \I__8864\ : InMux
    port map (
            O => \N__41063\,
            I => \N__41057\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__41060\,
            I => \N__41054\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__41057\,
            I => data_idxvec_8
        );

    \I__8861\ : Odrv4
    port map (
            O => \N__41054\,
            I => data_idxvec_8
        );

    \I__8860\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41046\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__41046\,
            I => \N__41042\
        );

    \I__8858\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41038\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__41042\,
            I => \N__41035\
        );

    \I__8856\ : InMux
    port map (
            O => \N__41041\,
            I => \N__41032\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__41038\,
            I => data_cntvec_8
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__41035\,
            I => data_cntvec_8
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__41032\,
            I => data_cntvec_8
        );

    \I__8852\ : InMux
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__41022\,
            I => \N__41017\
        );

    \I__8850\ : InMux
    port map (
            O => \N__41021\,
            I => \N__41012\
        );

    \I__8849\ : InMux
    port map (
            O => \N__41020\,
            I => \N__41012\
        );

    \I__8848\ : Odrv4
    port map (
            O => \N__41017\,
            I => req_data_cnt_11
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__41012\,
            I => req_data_cnt_11
        );

    \I__8846\ : CascadeMux
    port map (
            O => \N__41007\,
            I => \n8_adj_1571_cascade_\
        );

    \I__8845\ : InMux
    port map (
            O => \N__41004\,
            I => \N__41000\
        );

    \I__8844\ : InMux
    port map (
            O => \N__41003\,
            I => \N__40997\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__41000\,
            I => \N__40991\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__40997\,
            I => \N__40991\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40988\
        );

    \I__8840\ : Span4Mux_h
    port map (
            O => \N__40991\,
            I => \N__40985\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__40988\,
            I => data_index_2
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__40985\,
            I => data_index_2
        );

    \I__8837\ : InMux
    port map (
            O => \N__40980\,
            I => \N__40977\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40977\,
            I => \N__40973\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40976\,
            I => \N__40970\
        );

    \I__8834\ : Span4Mux_v
    port map (
            O => \N__40973\,
            I => \N__40964\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40970\,
            I => \N__40964\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40961\
        );

    \I__8831\ : Span4Mux_h
    port map (
            O => \N__40964\,
            I => \N__40958\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__40961\,
            I => buf_dds0_10
        );

    \I__8829\ : Odrv4
    port map (
            O => \N__40958\,
            I => buf_dds0_10
        );

    \I__8828\ : CascadeMux
    port map (
            O => \N__40953\,
            I => \N__40950\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40950\,
            I => \N__40946\
        );

    \I__8826\ : InMux
    port map (
            O => \N__40949\,
            I => \N__40943\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__40946\,
            I => data_idxvec_11
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40943\,
            I => data_idxvec_11
        );

    \I__8823\ : InMux
    port map (
            O => \N__40938\,
            I => \N__40933\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40937\,
            I => \N__40930\
        );

    \I__8821\ : InMux
    port map (
            O => \N__40936\,
            I => \N__40927\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__40933\,
            I => \N__40924\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__40930\,
            I => data_cntvec_11
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40927\,
            I => data_cntvec_11
        );

    \I__8817\ : Odrv4
    port map (
            O => \N__40924\,
            I => data_cntvec_11
        );

    \I__8816\ : InMux
    port map (
            O => \N__40917\,
            I => \N__40914\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__40914\,
            I => \N__40911\
        );

    \I__8814\ : Span4Mux_v
    port map (
            O => \N__40911\,
            I => \N__40908\
        );

    \I__8813\ : Span4Mux_h
    port map (
            O => \N__40908\,
            I => \N__40905\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__40905\,
            I => buf_data_iac_19
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__40902\,
            I => \n26_adj_1544_cascade_\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40899\,
            I => \N__40895\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40898\,
            I => \N__40892\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__40895\,
            I => \N__40886\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__40892\,
            I => \N__40881\
        );

    \I__8806\ : SRMux
    port map (
            O => \N__40891\,
            I => \N__40878\
        );

    \I__8805\ : InMux
    port map (
            O => \N__40890\,
            I => \N__40874\
        );

    \I__8804\ : SRMux
    port map (
            O => \N__40889\,
            I => \N__40871\
        );

    \I__8803\ : Span4Mux_h
    port map (
            O => \N__40886\,
            I => \N__40868\
        );

    \I__8802\ : InMux
    port map (
            O => \N__40885\,
            I => \N__40865\
        );

    \I__8801\ : InMux
    port map (
            O => \N__40884\,
            I => \N__40859\
        );

    \I__8800\ : Span4Mux_h
    port map (
            O => \N__40881\,
            I => \N__40854\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__40878\,
            I => \N__40854\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40877\,
            I => \N__40851\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__40874\,
            I => \N__40848\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__40871\,
            I => \N__40841\
        );

    \I__8795\ : Span4Mux_h
    port map (
            O => \N__40868\,
            I => \N__40841\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40865\,
            I => \N__40841\
        );

    \I__8793\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40834\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40834\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40834\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__40859\,
            I => acadc_rst
        );

    \I__8789\ : Odrv4
    port map (
            O => \N__40854\,
            I => acadc_rst
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__40851\,
            I => acadc_rst
        );

    \I__8787\ : Odrv12
    port map (
            O => \N__40848\,
            I => acadc_rst
        );

    \I__8786\ : Odrv4
    port map (
            O => \N__40841\,
            I => acadc_rst
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__40834\,
            I => acadc_rst
        );

    \I__8784\ : InMux
    port map (
            O => \N__40821\,
            I => \N__40817\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__40820\,
            I => \N__40814\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__40817\,
            I => \N__40810\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40814\,
            I => \N__40807\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40813\,
            I => \N__40804\
        );

    \I__8779\ : Span4Mux_h
    port map (
            O => \N__40810\,
            I => \N__40801\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40807\,
            I => \N__40798\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40804\,
            I => req_data_cnt_10
        );

    \I__8776\ : Odrv4
    port map (
            O => \N__40801\,
            I => req_data_cnt_10
        );

    \I__8775\ : Odrv4
    port map (
            O => \N__40798\,
            I => req_data_cnt_10
        );

    \I__8774\ : InMux
    port map (
            O => \N__40791\,
            I => \N__40788\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__40788\,
            I => n21088
        );

    \I__8772\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40782\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40782\,
            I => \N__40778\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40781\,
            I => \N__40774\
        );

    \I__8769\ : Span4Mux_v
    port map (
            O => \N__40778\,
            I => \N__40771\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40777\,
            I => \N__40768\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40774\,
            I => req_data_cnt_6
        );

    \I__8766\ : Odrv4
    port map (
            O => \N__40771\,
            I => req_data_cnt_6
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__40768\,
            I => req_data_cnt_6
        );

    \I__8764\ : InMux
    port map (
            O => \N__40761\,
            I => \N__40758\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__40758\,
            I => \N__40755\
        );

    \I__8762\ : Span4Mux_v
    port map (
            O => \N__40755\,
            I => \N__40751\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40754\,
            I => \N__40747\
        );

    \I__8760\ : Span4Mux_h
    port map (
            O => \N__40751\,
            I => \N__40744\
        );

    \I__8759\ : InMux
    port map (
            O => \N__40750\,
            I => \N__40741\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__40747\,
            I => buf_dds1_6
        );

    \I__8757\ : Odrv4
    port map (
            O => \N__40744\,
            I => buf_dds1_6
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__40741\,
            I => buf_dds1_6
        );

    \I__8755\ : InMux
    port map (
            O => \N__40734\,
            I => \N__40731\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40731\,
            I => \N__40726\
        );

    \I__8753\ : InMux
    port map (
            O => \N__40730\,
            I => \N__40721\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40721\
        );

    \I__8751\ : Odrv12
    port map (
            O => \N__40726\,
            I => buf_dds0_6
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__40721\,
            I => buf_dds0_6
        );

    \I__8749\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40712\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40715\,
            I => \N__40709\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__40712\,
            I => \N__40706\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__40709\,
            I => \N__40703\
        );

    \I__8745\ : Span4Mux_v
    port map (
            O => \N__40706\,
            I => \N__40700\
        );

    \I__8744\ : Span4Mux_v
    port map (
            O => \N__40703\,
            I => \N__40697\
        );

    \I__8743\ : Sp12to4
    port map (
            O => \N__40700\,
            I => \N__40691\
        );

    \I__8742\ : Sp12to4
    port map (
            O => \N__40697\,
            I => \N__40691\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40688\
        );

    \I__8740\ : Span12Mux_h
    port map (
            O => \N__40691\,
            I => \N__40685\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__40688\,
            I => buf_adcdata_iac_18
        );

    \I__8738\ : Odrv12
    port map (
            O => \N__40685\,
            I => buf_adcdata_iac_18
        );

    \I__8737\ : InMux
    port map (
            O => \N__40680\,
            I => \N__40677\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__40677\,
            I => n21073
        );

    \I__8735\ : CascadeMux
    port map (
            O => \N__40674\,
            I => \N__40671\
        );

    \I__8734\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40663\
        );

    \I__8733\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40660\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40669\,
            I => \N__40657\
        );

    \I__8731\ : InMux
    port map (
            O => \N__40668\,
            I => \N__40652\
        );

    \I__8730\ : InMux
    port map (
            O => \N__40667\,
            I => \N__40649\
        );

    \I__8729\ : InMux
    port map (
            O => \N__40666\,
            I => \N__40646\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__40663\,
            I => \N__40643\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40660\,
            I => \N__40638\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__40657\,
            I => \N__40638\
        );

    \I__8725\ : CascadeMux
    port map (
            O => \N__40656\,
            I => \N__40632\
        );

    \I__8724\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40628\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__40652\,
            I => \N__40625\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__40649\,
            I => \N__40622\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__40646\,
            I => \N__40619\
        );

    \I__8720\ : Span4Mux_v
    port map (
            O => \N__40643\,
            I => \N__40614\
        );

    \I__8719\ : Span4Mux_v
    port map (
            O => \N__40638\,
            I => \N__40614\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40611\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40608\
        );

    \I__8716\ : InMux
    port map (
            O => \N__40635\,
            I => \N__40605\
        );

    \I__8715\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40600\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40631\,
            I => \N__40600\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__40628\,
            I => \N__40597\
        );

    \I__8712\ : Span4Mux_h
    port map (
            O => \N__40625\,
            I => \N__40594\
        );

    \I__8711\ : Span4Mux_h
    port map (
            O => \N__40622\,
            I => \N__40591\
        );

    \I__8710\ : Span4Mux_v
    port map (
            O => \N__40619\,
            I => \N__40586\
        );

    \I__8709\ : Span4Mux_h
    port map (
            O => \N__40614\,
            I => \N__40586\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__40611\,
            I => n16891
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__40608\,
            I => n16891
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__40605\,
            I => n16891
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__40600\,
            I => n16891
        );

    \I__8704\ : Odrv12
    port map (
            O => \N__40597\,
            I => n16891
        );

    \I__8703\ : Odrv4
    port map (
            O => \N__40594\,
            I => n16891
        );

    \I__8702\ : Odrv4
    port map (
            O => \N__40591\,
            I => n16891
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__40586\,
            I => n16891
        );

    \I__8700\ : InMux
    port map (
            O => \N__40569\,
            I => \N__40564\
        );

    \I__8699\ : InMux
    port map (
            O => \N__40568\,
            I => \N__40561\
        );

    \I__8698\ : InMux
    port map (
            O => \N__40567\,
            I => \N__40558\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__40564\,
            I => \N__40551\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__40561\,
            I => \N__40551\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__40558\,
            I => \N__40551\
        );

    \I__8694\ : Span4Mux_h
    port map (
            O => \N__40551\,
            I => \N__40548\
        );

    \I__8693\ : Odrv4
    port map (
            O => \N__40548\,
            I => data_index_5
        );

    \I__8692\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40542\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__40542\,
            I => n22306
        );

    \I__8690\ : InMux
    port map (
            O => \N__40539\,
            I => \N__40536\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__40536\,
            I => \N__40533\
        );

    \I__8688\ : Odrv12
    port map (
            O => \N__40533\,
            I => n22420
        );

    \I__8687\ : InMux
    port map (
            O => \N__40530\,
            I => \N__40527\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__40527\,
            I => n22246
        );

    \I__8685\ : CascadeMux
    port map (
            O => \N__40524\,
            I => \n21092_cascade_\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__40521\,
            I => \n30_adj_1542_cascade_\
        );

    \I__8683\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40515\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__40515\,
            I => \N__40512\
        );

    \I__8681\ : Odrv12
    port map (
            O => \N__40512\,
            I => n21087
        );

    \I__8680\ : CascadeMux
    port map (
            O => \N__40509\,
            I => \n22357_cascade_\
        );

    \I__8679\ : CascadeMux
    port map (
            O => \N__40506\,
            I => \n22360_cascade_\
        );

    \I__8678\ : CascadeMux
    port map (
            O => \N__40503\,
            I => \n21137_cascade_\
        );

    \I__8677\ : CascadeMux
    port map (
            O => \N__40500\,
            I => \N__40497\
        );

    \I__8676\ : InMux
    port map (
            O => \N__40497\,
            I => \N__40494\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__40494\,
            I => \N__40491\
        );

    \I__8674\ : Odrv12
    port map (
            O => \N__40491\,
            I => n21072
        );

    \I__8673\ : InMux
    port map (
            O => \N__40488\,
            I => \N__40485\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__40485\,
            I => \N__40482\
        );

    \I__8671\ : Odrv12
    port map (
            O => \N__40482\,
            I => n22327
        );

    \I__8670\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40476\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__40476\,
            I => n22330
        );

    \I__8668\ : CascadeMux
    port map (
            O => \N__40473\,
            I => \n22288_cascade_\
        );

    \I__8667\ : InMux
    port map (
            O => \N__40470\,
            I => \N__40467\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__40467\,
            I => n22276
        );

    \I__8665\ : CascadeMux
    port map (
            O => \N__40464\,
            I => \n30_adj_1539_cascade_\
        );

    \I__8664\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40458\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__40458\,
            I => \N__40455\
        );

    \I__8662\ : Span4Mux_v
    port map (
            O => \N__40455\,
            I => \N__40452\
        );

    \I__8661\ : Span4Mux_v
    port map (
            O => \N__40452\,
            I => \N__40448\
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__40451\,
            I => \N__40445\
        );

    \I__8659\ : Span4Mux_h
    port map (
            O => \N__40448\,
            I => \N__40442\
        );

    \I__8658\ : InMux
    port map (
            O => \N__40445\,
            I => \N__40439\
        );

    \I__8657\ : Odrv4
    port map (
            O => \N__40442\,
            I => buf_adcdata_vdc_22
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__40439\,
            I => buf_adcdata_vdc_22
        );

    \I__8655\ : InMux
    port map (
            O => \N__40434\,
            I => \N__40430\
        );

    \I__8654\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40426\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__40430\,
            I => \N__40423\
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__40429\,
            I => \N__40420\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__40426\,
            I => \N__40415\
        );

    \I__8650\ : Span12Mux_v
    port map (
            O => \N__40423\,
            I => \N__40415\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40412\
        );

    \I__8648\ : Span12Mux_h
    port map (
            O => \N__40415\,
            I => \N__40409\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__40412\,
            I => buf_adcdata_vac_22
        );

    \I__8646\ : Odrv12
    port map (
            O => \N__40409\,
            I => buf_adcdata_vac_22
        );

    \I__8645\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40401\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40401\,
            I => \N__40398\
        );

    \I__8643\ : Odrv12
    port map (
            O => \N__40398\,
            I => n20_adj_1537
        );

    \I__8642\ : CascadeMux
    port map (
            O => \N__40395\,
            I => \n19_adj_1536_cascade_\
        );

    \I__8641\ : InMux
    port map (
            O => \N__40392\,
            I => \N__40389\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__40389\,
            I => n22285
        );

    \I__8639\ : InMux
    port map (
            O => \N__40386\,
            I => \N__40382\
        );

    \I__8638\ : CascadeMux
    port map (
            O => \N__40385\,
            I => \N__40379\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__40382\,
            I => \N__40376\
        );

    \I__8636\ : InMux
    port map (
            O => \N__40379\,
            I => \N__40373\
        );

    \I__8635\ : Sp12to4
    port map (
            O => \N__40376\,
            I => \N__40370\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__40373\,
            I => \N__40366\
        );

    \I__8633\ : Span12Mux_v
    port map (
            O => \N__40370\,
            I => \N__40363\
        );

    \I__8632\ : InMux
    port map (
            O => \N__40369\,
            I => \N__40360\
        );

    \I__8631\ : Span12Mux_h
    port map (
            O => \N__40366\,
            I => \N__40357\
        );

    \I__8630\ : Span12Mux_h
    port map (
            O => \N__40363\,
            I => \N__40354\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__40360\,
            I => buf_adcdata_iac_20
        );

    \I__8628\ : Odrv12
    port map (
            O => \N__40357\,
            I => buf_adcdata_iac_20
        );

    \I__8627\ : Odrv12
    port map (
            O => \N__40354\,
            I => buf_adcdata_iac_20
        );

    \I__8626\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40343\
        );

    \I__8625\ : InMux
    port map (
            O => \N__40346\,
            I => \N__40340\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__40343\,
            I => \N__40336\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__40340\,
            I => \N__40333\
        );

    \I__8622\ : InMux
    port map (
            O => \N__40339\,
            I => \N__40330\
        );

    \I__8621\ : Span12Mux_h
    port map (
            O => \N__40336\,
            I => \N__40327\
        );

    \I__8620\ : Odrv4
    port map (
            O => \N__40333\,
            I => buf_dds0_12
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__40330\,
            I => buf_dds0_12
        );

    \I__8618\ : Odrv12
    port map (
            O => \N__40327\,
            I => buf_dds0_12
        );

    \I__8617\ : CascadeMux
    port map (
            O => \N__40320\,
            I => \n22303_cascade_\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40317\,
            I => \N__40313\
        );

    \I__8615\ : InMux
    port map (
            O => \N__40316\,
            I => \N__40310\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__40313\,
            I => \N__40306\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__40310\,
            I => \N__40303\
        );

    \I__8612\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40300\
        );

    \I__8611\ : Span4Mux_h
    port map (
            O => \N__40306\,
            I => \N__40297\
        );

    \I__8610\ : Span4Mux_v
    port map (
            O => \N__40303\,
            I => \N__40294\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__40300\,
            I => buf_dds1_12
        );

    \I__8608\ : Odrv4
    port map (
            O => \N__40297\,
            I => buf_dds1_12
        );

    \I__8607\ : Odrv4
    port map (
            O => \N__40294\,
            I => buf_dds1_12
        );

    \I__8606\ : InMux
    port map (
            O => \N__40287\,
            I => \N__40284\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__40284\,
            I => \N__40281\
        );

    \I__8604\ : Span12Mux_v
    port map (
            O => \N__40281\,
            I => \N__40278\
        );

    \I__8603\ : Odrv12
    port map (
            O => \N__40278\,
            I => n21309
        );

    \I__8602\ : CascadeMux
    port map (
            O => \N__40275\,
            I => \N__40272\
        );

    \I__8601\ : InMux
    port map (
            O => \N__40272\,
            I => \N__40269\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__40269\,
            I => \N__40266\
        );

    \I__8599\ : Span4Mux_h
    port map (
            O => \N__40266\,
            I => \N__40263\
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__40263\,
            I => n23_adj_1541
        );

    \I__8597\ : CascadeMux
    port map (
            O => \N__40260\,
            I => \N__40257\
        );

    \I__8596\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40254\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__40254\,
            I => n21568
        );

    \I__8594\ : InMux
    port map (
            O => \N__40251\,
            I => \N__40248\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__40248\,
            I => n22243
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__40245\,
            I => \n22237_cascade_\
        );

    \I__8591\ : InMux
    port map (
            O => \N__40242\,
            I => \N__40238\
        );

    \I__8590\ : InMux
    port map (
            O => \N__40241\,
            I => \N__40234\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__40238\,
            I => \N__40231\
        );

    \I__8588\ : InMux
    port map (
            O => \N__40237\,
            I => \N__40228\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__40234\,
            I => \N__40225\
        );

    \I__8586\ : Span4Mux_h
    port map (
            O => \N__40231\,
            I => \N__40222\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__40228\,
            I => buf_dds1_9
        );

    \I__8584\ : Odrv4
    port map (
            O => \N__40225\,
            I => buf_dds1_9
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__40222\,
            I => buf_dds1_9
        );

    \I__8582\ : InMux
    port map (
            O => \N__40215\,
            I => \N__40212\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__8580\ : Odrv12
    port map (
            O => \N__40209\,
            I => buf_data_iac_17
        );

    \I__8579\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40203\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__40203\,
            I => \N__40200\
        );

    \I__8577\ : Span4Mux_h
    port map (
            O => \N__40200\,
            I => \N__40197\
        );

    \I__8576\ : Span4Mux_v
    port map (
            O => \N__40197\,
            I => \N__40194\
        );

    \I__8575\ : Odrv4
    port map (
            O => \N__40194\,
            I => n22378
        );

    \I__8574\ : CascadeMux
    port map (
            O => \N__40191\,
            I => \n21062_cascade_\
        );

    \I__8573\ : InMux
    port map (
            O => \N__40188\,
            I => \N__40185\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__40185\,
            I => n22240
        );

    \I__8571\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40179\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__40179\,
            I => \N__40176\
        );

    \I__8569\ : Span4Mux_h
    port map (
            O => \N__40176\,
            I => \N__40173\
        );

    \I__8568\ : Span4Mux_h
    port map (
            O => \N__40173\,
            I => \N__40170\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__40170\,
            I => n22444
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__40167\,
            I => \n22447_cascade_\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__40164\,
            I => \n22450_cascade_\
        );

    \I__8564\ : CascadeMux
    port map (
            O => \N__40161\,
            I => \N__40157\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__40160\,
            I => \N__40152\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40149\
        );

    \I__8561\ : CascadeMux
    port map (
            O => \N__40156\,
            I => \N__40146\
        );

    \I__8560\ : CascadeMux
    port map (
            O => \N__40155\,
            I => \N__40142\
        );

    \I__8559\ : InMux
    port map (
            O => \N__40152\,
            I => \N__40139\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__40149\,
            I => \N__40136\
        );

    \I__8557\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40132\
        );

    \I__8556\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40129\
        );

    \I__8555\ : InMux
    port map (
            O => \N__40142\,
            I => \N__40126\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__40139\,
            I => \N__40123\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__40136\,
            I => \N__40116\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40135\,
            I => \N__40113\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__40132\,
            I => \N__40110\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__40129\,
            I => \N__40107\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__40126\,
            I => \N__40104\
        );

    \I__8548\ : Span4Mux_v
    port map (
            O => \N__40123\,
            I => \N__40101\
        );

    \I__8547\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40098\
        );

    \I__8546\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40095\
        );

    \I__8545\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40092\
        );

    \I__8544\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40089\
        );

    \I__8543\ : Span4Mux_h
    port map (
            O => \N__40116\,
            I => \N__40084\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__40113\,
            I => \N__40084\
        );

    \I__8541\ : Span4Mux_v
    port map (
            O => \N__40110\,
            I => \N__40081\
        );

    \I__8540\ : Span4Mux_h
    port map (
            O => \N__40107\,
            I => \N__40078\
        );

    \I__8539\ : Span4Mux_h
    port map (
            O => \N__40104\,
            I => \N__40071\
        );

    \I__8538\ : Span4Mux_h
    port map (
            O => \N__40101\,
            I => \N__40071\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__40098\,
            I => \N__40071\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__40095\,
            I => \N__40068\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__40092\,
            I => \N__40065\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__40089\,
            I => \N__40054\
        );

    \I__8533\ : Span4Mux_h
    port map (
            O => \N__40084\,
            I => \N__40054\
        );

    \I__8532\ : Span4Mux_h
    port map (
            O => \N__40081\,
            I => \N__40054\
        );

    \I__8531\ : Span4Mux_v
    port map (
            O => \N__40078\,
            I => \N__40054\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__40071\,
            I => \N__40054\
        );

    \I__8529\ : Span12Mux_h
    port map (
            O => \N__40068\,
            I => \N__40051\
        );

    \I__8528\ : Span12Mux_v
    port map (
            O => \N__40065\,
            I => \N__40048\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__40054\,
            I => \N__40045\
        );

    \I__8526\ : Odrv12
    port map (
            O => \N__40051\,
            I => comm_buf_0_1
        );

    \I__8525\ : Odrv12
    port map (
            O => \N__40048\,
            I => comm_buf_0_1
        );

    \I__8524\ : Odrv4
    port map (
            O => \N__40045\,
            I => comm_buf_0_1
        );

    \I__8523\ : CascadeMux
    port map (
            O => \N__40038\,
            I => \N__40035\
        );

    \I__8522\ : InMux
    port map (
            O => \N__40035\,
            I => \N__40032\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__40032\,
            I => n30
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__40029\,
            I => \N__40026\
        );

    \I__8519\ : InMux
    port map (
            O => \N__40026\,
            I => \N__40023\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__40023\,
            I => n21272
        );

    \I__8517\ : InMux
    port map (
            O => \N__40020\,
            I => \N__40017\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__40017\,
            I => \N__40014\
        );

    \I__8515\ : Span4Mux_h
    port map (
            O => \N__40014\,
            I => \N__40011\
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__40011\,
            I => n23_adj_1538
        );

    \I__8513\ : CascadeMux
    port map (
            O => \N__40008\,
            I => \n22273_cascade_\
        );

    \I__8512\ : InMux
    port map (
            O => \N__40005\,
            I => \N__40002\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__40002\,
            I => \N__39999\
        );

    \I__8510\ : Span4Mux_h
    port map (
            O => \N__39999\,
            I => \N__39996\
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__39996\,
            I => n21286
        );

    \I__8508\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39990\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__39990\,
            I => \N__39987\
        );

    \I__8506\ : Span4Mux_h
    port map (
            O => \N__39987\,
            I => \N__39984\
        );

    \I__8505\ : Span4Mux_h
    port map (
            O => \N__39984\,
            I => \N__39981\
        );

    \I__8504\ : Odrv4
    port map (
            O => \N__39981\,
            I => n17_adj_1535
        );

    \I__8503\ : CascadeMux
    port map (
            O => \N__39978\,
            I => \N__39975\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39975\,
            I => \N__39972\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39972\,
            I => \N__39969\
        );

    \I__8500\ : Span4Mux_v
    port map (
            O => \N__39969\,
            I => \N__39966\
        );

    \I__8499\ : Sp12to4
    port map (
            O => \N__39966\,
            I => \N__39963\
        );

    \I__8498\ : Odrv12
    port map (
            O => \N__39963\,
            I => n16_adj_1534
        );

    \I__8497\ : CascadeMux
    port map (
            O => \N__39960\,
            I => \N__39957\
        );

    \I__8496\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39954\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39954\,
            I => \N__39951\
        );

    \I__8494\ : Span12Mux_v
    port map (
            O => \N__39951\,
            I => \N__39948\
        );

    \I__8493\ : Span12Mux_h
    port map (
            O => \N__39948\,
            I => \N__39945\
        );

    \I__8492\ : Odrv12
    port map (
            O => \N__39945\,
            I => buf_data_vac_7
        );

    \I__8491\ : InMux
    port map (
            O => \N__39942\,
            I => \N__39939\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__39939\,
            I => \N__39936\
        );

    \I__8489\ : Span4Mux_v
    port map (
            O => \N__39936\,
            I => \N__39933\
        );

    \I__8488\ : Odrv4
    port map (
            O => \N__39933\,
            I => comm_buf_5_7
        );

    \I__8487\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39927\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__39927\,
            I => \N__39924\
        );

    \I__8485\ : Span12Mux_v
    port map (
            O => \N__39924\,
            I => \N__39921\
        );

    \I__8484\ : Span12Mux_h
    port map (
            O => \N__39921\,
            I => \N__39918\
        );

    \I__8483\ : Odrv12
    port map (
            O => \N__39918\,
            I => buf_data_vac_6
        );

    \I__8482\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__39912\,
            I => \N__39909\
        );

    \I__8480\ : Span12Mux_v
    port map (
            O => \N__39909\,
            I => \N__39906\
        );

    \I__8479\ : Span12Mux_h
    port map (
            O => \N__39906\,
            I => \N__39903\
        );

    \I__8478\ : Odrv12
    port map (
            O => \N__39903\,
            I => buf_data_vac_5
        );

    \I__8477\ : InMux
    port map (
            O => \N__39900\,
            I => \N__39897\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39897\,
            I => \N__39894\
        );

    \I__8475\ : Span12Mux_v
    port map (
            O => \N__39894\,
            I => \N__39891\
        );

    \I__8474\ : Span12Mux_h
    port map (
            O => \N__39891\,
            I => \N__39888\
        );

    \I__8473\ : Odrv12
    port map (
            O => \N__39888\,
            I => buf_data_vac_4
        );

    \I__8472\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39882\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__39882\,
            I => \N__39879\
        );

    \I__8470\ : Odrv4
    port map (
            O => \N__39879\,
            I => comm_buf_5_4
        );

    \I__8469\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39873\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39873\,
            I => \N__39870\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__39870\,
            I => \N__39867\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__39867\,
            I => \N__39864\
        );

    \I__8465\ : Odrv4
    port map (
            O => \N__39864\,
            I => buf_data_vac_3
        );

    \I__8464\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39858\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__39858\,
            I => \N__39855\
        );

    \I__8462\ : Span4Mux_h
    port map (
            O => \N__39855\,
            I => \N__39852\
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__39852\,
            I => comm_buf_5_3
        );

    \I__8460\ : InMux
    port map (
            O => \N__39849\,
            I => \N__39846\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__39846\,
            I => \N__39843\
        );

    \I__8458\ : Span4Mux_v
    port map (
            O => \N__39843\,
            I => \N__39840\
        );

    \I__8457\ : Span4Mux_h
    port map (
            O => \N__39840\,
            I => \N__39837\
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__39837\,
            I => buf_data_vac_2
        );

    \I__8455\ : InMux
    port map (
            O => \N__39834\,
            I => \N__39831\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__39831\,
            I => comm_buf_5_2
        );

    \I__8453\ : InMux
    port map (
            O => \N__39828\,
            I => \N__39825\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__39825\,
            I => \N__39822\
        );

    \I__8451\ : Span4Mux_h
    port map (
            O => \N__39822\,
            I => \N__39819\
        );

    \I__8450\ : Span4Mux_h
    port map (
            O => \N__39819\,
            I => \N__39816\
        );

    \I__8449\ : Odrv4
    port map (
            O => \N__39816\,
            I => buf_data_vac_1
        );

    \I__8448\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39810\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__39810\,
            I => comm_buf_5_1
        );

    \I__8446\ : IoInMux
    port map (
            O => \N__39807\,
            I => \N__39804\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39804\,
            I => \N__39801\
        );

    \I__8444\ : Span4Mux_s3_v
    port map (
            O => \N__39801\,
            I => \N__39797\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39794\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__39797\,
            I => \N__39791\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39794\,
            I => \N__39788\
        );

    \I__8440\ : Span4Mux_v
    port map (
            O => \N__39791\,
            I => \N__39784\
        );

    \I__8439\ : Span4Mux_h
    port map (
            O => \N__39788\,
            I => \N__39781\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39787\,
            I => \N__39778\
        );

    \I__8437\ : Span4Mux_v
    port map (
            O => \N__39784\,
            I => \N__39773\
        );

    \I__8436\ : Span4Mux_h
    port map (
            O => \N__39781\,
            I => \N__39773\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__39778\,
            I => \IAC_OSR1\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__39773\,
            I => \IAC_OSR1\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39768\,
            I => \N__39765\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__39765\,
            I => \N__39762\
        );

    \I__8431\ : Span4Mux_h
    port map (
            O => \N__39762\,
            I => \N__39758\
        );

    \I__8430\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39755\
        );

    \I__8429\ : Span4Mux_h
    port map (
            O => \N__39758\,
            I => \N__39749\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39755\,
            I => \N__39749\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39746\
        );

    \I__8426\ : Span4Mux_h
    port map (
            O => \N__39749\,
            I => \N__39743\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__39746\,
            I => buf_adcdata_iac_17
        );

    \I__8424\ : Odrv4
    port map (
            O => \N__39743\,
            I => buf_adcdata_iac_17
        );

    \I__8423\ : InMux
    port map (
            O => \N__39738\,
            I => \N__39735\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39735\,
            I => \N__39732\
        );

    \I__8421\ : Span4Mux_v
    port map (
            O => \N__39732\,
            I => \N__39729\
        );

    \I__8420\ : Span4Mux_h
    port map (
            O => \N__39729\,
            I => \N__39724\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39728\,
            I => \N__39721\
        );

    \I__8418\ : InMux
    port map (
            O => \N__39727\,
            I => \N__39718\
        );

    \I__8417\ : Span4Mux_v
    port map (
            O => \N__39724\,
            I => \N__39715\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__39721\,
            I => buf_dds0_9
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__39718\,
            I => buf_dds0_9
        );

    \I__8414\ : Odrv4
    port map (
            O => \N__39715\,
            I => buf_dds0_9
        );

    \I__8413\ : InMux
    port map (
            O => \N__39708\,
            I => \N__39705\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__39705\,
            I => \N__39702\
        );

    \I__8411\ : Span4Mux_h
    port map (
            O => \N__39702\,
            I => \N__39699\
        );

    \I__8410\ : Odrv4
    port map (
            O => \N__39699\,
            I => comm_buf_2_2
        );

    \I__8409\ : CascadeMux
    port map (
            O => \N__39696\,
            I => \n22393_cascade_\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39693\,
            I => \N__39690\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__39690\,
            I => \N__39687\
        );

    \I__8406\ : Span4Mux_v
    port map (
            O => \N__39687\,
            I => \N__39683\
        );

    \I__8405\ : InMux
    port map (
            O => \N__39686\,
            I => \N__39680\
        );

    \I__8404\ : Span4Mux_h
    port map (
            O => \N__39683\,
            I => \N__39677\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__39680\,
            I => comm_buf_6_2
        );

    \I__8402\ : Odrv4
    port map (
            O => \N__39677\,
            I => comm_buf_6_2
        );

    \I__8401\ : CascadeMux
    port map (
            O => \N__39672\,
            I => \n4_adj_1595_cascade_\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39669\,
            I => \N__39666\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39666\,
            I => n22396
        );

    \I__8398\ : CascadeMux
    port map (
            O => \N__39663\,
            I => \n21196_cascade_\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39660\,
            I => \N__39651\
        );

    \I__8396\ : InMux
    port map (
            O => \N__39659\,
            I => \N__39651\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39658\,
            I => \N__39651\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__39651\,
            I => \N__39648\
        );

    \I__8393\ : Span4Mux_v
    port map (
            O => \N__39648\,
            I => \N__39645\
        );

    \I__8392\ : Odrv4
    port map (
            O => \N__39645\,
            I => comm_tx_buf_2
        );

    \I__8391\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39639\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__39639\,
            I => \N__39635\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39638\,
            I => \N__39632\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__39635\,
            I => \N__39629\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39632\,
            I => comm_buf_6_1
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__39629\,
            I => comm_buf_6_1
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__39624\,
            I => \n4_adj_1596_cascade_\
        );

    \I__8384\ : InMux
    port map (
            O => \N__39621\,
            I => \N__39618\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__39618\,
            I => \N__39615\
        );

    \I__8382\ : Span4Mux_h
    port map (
            O => \N__39615\,
            I => \N__39612\
        );

    \I__8381\ : Odrv4
    port map (
            O => \N__39612\,
            I => n22252
        );

    \I__8380\ : CascadeMux
    port map (
            O => \N__39609\,
            I => \n21052_cascade_\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39606\,
            I => \N__39597\
        );

    \I__8378\ : InMux
    port map (
            O => \N__39605\,
            I => \N__39597\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39604\,
            I => \N__39597\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__39597\,
            I => \N__39594\
        );

    \I__8375\ : Span4Mux_v
    port map (
            O => \N__39594\,
            I => \N__39591\
        );

    \I__8374\ : Odrv4
    port map (
            O => \N__39591\,
            I => comm_tx_buf_1
        );

    \I__8373\ : InMux
    port map (
            O => \N__39588\,
            I => \N__39585\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__39585\,
            I => \N__39582\
        );

    \I__8371\ : Span4Mux_h
    port map (
            O => \N__39582\,
            I => \N__39579\
        );

    \I__8370\ : Span4Mux_h
    port map (
            O => \N__39579\,
            I => \N__39576\
        );

    \I__8369\ : Odrv4
    port map (
            O => \N__39576\,
            I => buf_data_vac_0
        );

    \I__8368\ : SRMux
    port map (
            O => \N__39573\,
            I => \N__39570\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__39570\,
            I => \N__39566\
        );

    \I__8366\ : SRMux
    port map (
            O => \N__39569\,
            I => \N__39563\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__39566\,
            I => \N__39560\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__39563\,
            I => \N__39557\
        );

    \I__8363\ : Span4Mux_h
    port map (
            O => \N__39560\,
            I => \N__39554\
        );

    \I__8362\ : Span4Mux_v
    port map (
            O => \N__39557\,
            I => \N__39551\
        );

    \I__8361\ : Odrv4
    port map (
            O => \N__39554\,
            I => n20378
        );

    \I__8360\ : Odrv4
    port map (
            O => \N__39551\,
            I => n20378
        );

    \I__8359\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39543\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__8357\ : Odrv12
    port map (
            O => \N__39540\,
            I => comm_buf_2_4
        );

    \I__8356\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39534\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__39534\,
            I => \N__39531\
        );

    \I__8354\ : Span4Mux_h
    port map (
            O => \N__39531\,
            I => \N__39527\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39530\,
            I => \N__39524\
        );

    \I__8352\ : Span4Mux_h
    port map (
            O => \N__39527\,
            I => \N__39521\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39524\,
            I => comm_buf_6_4
        );

    \I__8350\ : Odrv4
    port map (
            O => \N__39521\,
            I => comm_buf_6_4
        );

    \I__8349\ : CascadeMux
    port map (
            O => \N__39516\,
            I => \n21538_cascade_\
        );

    \I__8348\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39510\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__39510\,
            I => n1_adj_1591
        );

    \I__8346\ : CascadeMux
    port map (
            O => \N__39507\,
            I => \n22369_cascade_\
        );

    \I__8345\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39501\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__39501\,
            I => n2_adj_1592
        );

    \I__8343\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39495\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__39495\,
            I => n4_adj_1593
        );

    \I__8341\ : SRMux
    port map (
            O => \N__39492\,
            I => \N__39489\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__39489\,
            I => \N__39486\
        );

    \I__8339\ : Odrv4
    port map (
            O => \N__39486\,
            I => \comm_spi.data_tx_7__N_783\
        );

    \I__8338\ : InMux
    port map (
            O => \N__39483\,
            I => \N__39480\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__39480\,
            I => \N__39477\
        );

    \I__8336\ : Span4Mux_v
    port map (
            O => \N__39477\,
            I => \N__39472\
        );

    \I__8335\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39467\
        );

    \I__8334\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39467\
        );

    \I__8333\ : Odrv4
    port map (
            O => \N__39472\,
            I => comm_tx_buf_4
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__39467\,
            I => comm_tx_buf_4
        );

    \I__8331\ : SRMux
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__39459\,
            I => \N__39456\
        );

    \I__8329\ : Span4Mux_v
    port map (
            O => \N__39456\,
            I => \N__39453\
        );

    \I__8328\ : Sp12to4
    port map (
            O => \N__39453\,
            I => \N__39450\
        );

    \I__8327\ : Odrv12
    port map (
            O => \N__39450\,
            I => \comm_spi.data_tx_7__N_769\
        );

    \I__8326\ : CEMux
    port map (
            O => \N__39447\,
            I => \N__39444\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__39444\,
            I => \N__39441\
        );

    \I__8324\ : Odrv12
    port map (
            O => \N__39441\,
            I => n11741
        );

    \I__8323\ : InMux
    port map (
            O => \N__39438\,
            I => \N__39435\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39435\,
            I => n20992
        );

    \I__8321\ : CascadeMux
    port map (
            O => \N__39432\,
            I => \n9255_cascade_\
        );

    \I__8320\ : SRMux
    port map (
            O => \N__39429\,
            I => \N__39426\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39426\,
            I => \N__39423\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__39423\,
            I => \N__39420\
        );

    \I__8317\ : Odrv4
    port map (
            O => \N__39420\,
            I => n14737
        );

    \I__8316\ : SRMux
    port map (
            O => \N__39417\,
            I => \N__39414\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__39414\,
            I => \N__39410\
        );

    \I__8314\ : SRMux
    port map (
            O => \N__39413\,
            I => \N__39407\
        );

    \I__8313\ : Span4Mux_v
    port map (
            O => \N__39410\,
            I => \N__39404\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__39407\,
            I => \N__39401\
        );

    \I__8311\ : Span4Mux_h
    port map (
            O => \N__39404\,
            I => \N__39398\
        );

    \I__8310\ : Span12Mux_v
    port map (
            O => \N__39401\,
            I => \N__39395\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__39398\,
            I => flagcntwd
        );

    \I__8308\ : Odrv12
    port map (
            O => \N__39395\,
            I => flagcntwd
        );

    \I__8307\ : CEMux
    port map (
            O => \N__39390\,
            I => \N__39387\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__39387\,
            I => \N__39384\
        );

    \I__8305\ : Span4Mux_h
    port map (
            O => \N__39384\,
            I => \N__39381\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__39381\,
            I => n11390
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__39378\,
            I => \n12336_cascade_\
        );

    \I__8302\ : SRMux
    port map (
            O => \N__39375\,
            I => \N__39372\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39369\
        );

    \I__8300\ : Span4Mux_h
    port map (
            O => \N__39369\,
            I => \N__39366\
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__39366\,
            I => \comm_spi.data_tx_7__N_772\
        );

    \I__8298\ : SRMux
    port map (
            O => \N__39363\,
            I => \N__39360\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__39360\,
            I => \N__39357\
        );

    \I__8296\ : Span4Mux_h
    port map (
            O => \N__39357\,
            I => \N__39354\
        );

    \I__8295\ : Odrv4
    port map (
            O => \N__39354\,
            I => \comm_spi.data_tx_7__N_792\
        );

    \I__8294\ : InMux
    port map (
            O => \N__39351\,
            I => \N__39348\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__39348\,
            I => \N__39345\
        );

    \I__8292\ : Sp12to4
    port map (
            O => \N__39345\,
            I => \N__39341\
        );

    \I__8291\ : InMux
    port map (
            O => \N__39344\,
            I => \N__39338\
        );

    \I__8290\ : Span12Mux_v
    port map (
            O => \N__39341\,
            I => \N__39334\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__39338\,
            I => \N__39331\
        );

    \I__8288\ : InMux
    port map (
            O => \N__39337\,
            I => \N__39328\
        );

    \I__8287\ : Odrv12
    port map (
            O => \N__39334\,
            I => \comm_spi.n22881\
        );

    \I__8286\ : Odrv4
    port map (
            O => \N__39331\,
            I => \comm_spi.n22881\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__39328\,
            I => \comm_spi.n22881\
        );

    \I__8284\ : SRMux
    port map (
            O => \N__39321\,
            I => \N__39318\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__39318\,
            I => \N__39315\
        );

    \I__8282\ : Span12Mux_s9_v
    port map (
            O => \N__39315\,
            I => \N__39312\
        );

    \I__8281\ : Odrv12
    port map (
            O => \N__39312\,
            I => \comm_spi.data_tx_7__N_789\
        );

    \I__8280\ : SRMux
    port map (
            O => \N__39309\,
            I => \N__39306\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39306\,
            I => \N__39303\
        );

    \I__8278\ : Span4Mux_v
    port map (
            O => \N__39303\,
            I => \N__39300\
        );

    \I__8277\ : Span4Mux_v
    port map (
            O => \N__39300\,
            I => \N__39297\
        );

    \I__8276\ : Span4Mux_v
    port map (
            O => \N__39297\,
            I => \N__39294\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__39294\,
            I => \comm_spi.data_tx_7__N_771\
        );

    \I__8274\ : InMux
    port map (
            O => \N__39291\,
            I => \N__39288\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__39288\,
            I => \N__39284\
        );

    \I__8272\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39281\
        );

    \I__8271\ : Span4Mux_v
    port map (
            O => \N__39284\,
            I => \N__39276\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__39281\,
            I => \N__39276\
        );

    \I__8269\ : Span4Mux_v
    port map (
            O => \N__39276\,
            I => \N__39272\
        );

    \I__8268\ : InMux
    port map (
            O => \N__39275\,
            I => \N__39269\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__39272\,
            I => \comm_spi.n22878\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__39269\,
            I => \comm_spi.n22878\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__39264\,
            I => \N__39261\
        );

    \I__8264\ : InMux
    port map (
            O => \N__39261\,
            I => \N__39256\
        );

    \I__8263\ : InMux
    port map (
            O => \N__39260\,
            I => \N__39251\
        );

    \I__8262\ : InMux
    port map (
            O => \N__39259\,
            I => \N__39251\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__39256\,
            I => wdtick_cnt_2
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__39251\,
            I => wdtick_cnt_2
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__39246\,
            I => \N__39242\
        );

    \I__8258\ : InMux
    port map (
            O => \N__39245\,
            I => \N__39237\
        );

    \I__8257\ : InMux
    port map (
            O => \N__39242\,
            I => \N__39230\
        );

    \I__8256\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39230\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39230\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__39237\,
            I => wdtick_cnt_0
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__39230\,
            I => wdtick_cnt_0
        );

    \I__8252\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39219\
        );

    \I__8251\ : InMux
    port map (
            O => \N__39224\,
            I => \N__39212\
        );

    \I__8250\ : InMux
    port map (
            O => \N__39223\,
            I => \N__39212\
        );

    \I__8249\ : InMux
    port map (
            O => \N__39222\,
            I => \N__39212\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__39219\,
            I => wdtick_cnt_1
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__39212\,
            I => wdtick_cnt_1
        );

    \I__8246\ : IoInMux
    port map (
            O => \N__39207\,
            I => \N__39202\
        );

    \I__8245\ : ClkMux
    port map (
            O => \N__39206\,
            I => \N__39199\
        );

    \I__8244\ : ClkMux
    port map (
            O => \N__39205\,
            I => \N__39196\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__39202\,
            I => \N__39193\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39199\,
            I => \N__39190\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__39196\,
            I => \N__39187\
        );

    \I__8240\ : Span4Mux_s3_v
    port map (
            O => \N__39193\,
            I => \N__39184\
        );

    \I__8239\ : Span4Mux_v
    port map (
            O => \N__39190\,
            I => \N__39181\
        );

    \I__8238\ : Span4Mux_v
    port map (
            O => \N__39187\,
            I => \N__39178\
        );

    \I__8237\ : Sp12to4
    port map (
            O => \N__39184\,
            I => \N__39175\
        );

    \I__8236\ : Span4Mux_h
    port map (
            O => \N__39181\,
            I => \N__39172\
        );

    \I__8235\ : Span4Mux_h
    port map (
            O => \N__39178\,
            I => \N__39169\
        );

    \I__8234\ : Span12Mux_s10_h
    port map (
            O => \N__39175\,
            I => \N__39165\
        );

    \I__8233\ : Span4Mux_h
    port map (
            O => \N__39172\,
            I => \N__39162\
        );

    \I__8232\ : Span4Mux_v
    port map (
            O => \N__39169\,
            I => \N__39159\
        );

    \I__8231\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39156\
        );

    \I__8230\ : Odrv12
    port map (
            O => \N__39165\,
            I => \TEST_LED\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__39162\,
            I => \TEST_LED\
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__39159\,
            I => \TEST_LED\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__39156\,
            I => \TEST_LED\
        );

    \I__8226\ : InMux
    port map (
            O => \N__39147\,
            I => \N__39143\
        );

    \I__8225\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39140\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__39143\,
            I => \comm_spi.n14627\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__39140\,
            I => \comm_spi.n14627\
        );

    \I__8222\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39132\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__39132\,
            I => \N__39128\
        );

    \I__8220\ : InMux
    port map (
            O => \N__39131\,
            I => \N__39125\
        );

    \I__8219\ : Span4Mux_v
    port map (
            O => \N__39128\,
            I => \N__39122\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__39125\,
            I => \N__39119\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__39122\,
            I => \N__39115\
        );

    \I__8216\ : Span4Mux_v
    port map (
            O => \N__39119\,
            I => \N__39112\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39118\,
            I => \N__39109\
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__39115\,
            I => \comm_spi.n22875\
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__39112\,
            I => \comm_spi.n22875\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__39109\,
            I => \comm_spi.n22875\
        );

    \I__8211\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39099\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__39099\,
            I => \N__39096\
        );

    \I__8209\ : Span4Mux_h
    port map (
            O => \N__39096\,
            I => \N__39092\
        );

    \I__8208\ : InMux
    port map (
            O => \N__39095\,
            I => \N__39089\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__39092\,
            I => \N__39086\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__39089\,
            I => \N__39083\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__39086\,
            I => \comm_spi.n14626\
        );

    \I__8204\ : Odrv12
    port map (
            O => \N__39083\,
            I => \comm_spi.n14626\
        );

    \I__8203\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39073\
        );

    \I__8202\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39070\
        );

    \I__8201\ : InMux
    port map (
            O => \N__39076\,
            I => \N__39067\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__39073\,
            I => data_index_9
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__39070\,
            I => data_index_9
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__39067\,
            I => data_index_9
        );

    \I__8197\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39057\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__39057\,
            I => n8_adj_1559
        );

    \I__8195\ : InMux
    port map (
            O => \N__39054\,
            I => \N__39050\
        );

    \I__8194\ : InMux
    port map (
            O => \N__39053\,
            I => \N__39047\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__39050\,
            I => n7_adj_1558
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__39047\,
            I => n7_adj_1558
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__39042\,
            I => \n8_adj_1559_cascade_\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__39039\,
            I => \N__39036\
        );

    \I__8189\ : CascadeBuf
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__8188\ : CascadeMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__8187\ : CascadeBuf
    port map (
            O => \N__39030\,
            I => \N__39027\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__39027\,
            I => \N__39024\
        );

    \I__8185\ : CascadeBuf
    port map (
            O => \N__39024\,
            I => \N__39021\
        );

    \I__8184\ : CascadeMux
    port map (
            O => \N__39021\,
            I => \N__39018\
        );

    \I__8183\ : CascadeBuf
    port map (
            O => \N__39018\,
            I => \N__39015\
        );

    \I__8182\ : CascadeMux
    port map (
            O => \N__39015\,
            I => \N__39012\
        );

    \I__8181\ : CascadeBuf
    port map (
            O => \N__39012\,
            I => \N__39009\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__8179\ : CascadeBuf
    port map (
            O => \N__39006\,
            I => \N__39003\
        );

    \I__8178\ : CascadeMux
    port map (
            O => \N__39003\,
            I => \N__39000\
        );

    \I__8177\ : CascadeBuf
    port map (
            O => \N__39000\,
            I => \N__38996\
        );

    \I__8176\ : CascadeMux
    port map (
            O => \N__38999\,
            I => \N__38993\
        );

    \I__8175\ : CascadeMux
    port map (
            O => \N__38996\,
            I => \N__38990\
        );

    \I__8174\ : CascadeBuf
    port map (
            O => \N__38993\,
            I => \N__38987\
        );

    \I__8173\ : CascadeBuf
    port map (
            O => \N__38990\,
            I => \N__38984\
        );

    \I__8172\ : CascadeMux
    port map (
            O => \N__38987\,
            I => \N__38981\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__38984\,
            I => \N__38978\
        );

    \I__8170\ : InMux
    port map (
            O => \N__38981\,
            I => \N__38975\
        );

    \I__8169\ : CascadeBuf
    port map (
            O => \N__38978\,
            I => \N__38972\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__38975\,
            I => \N__38969\
        );

    \I__8167\ : CascadeMux
    port map (
            O => \N__38972\,
            I => \N__38966\
        );

    \I__8166\ : Span12Mux_h
    port map (
            O => \N__38969\,
            I => \N__38963\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38960\
        );

    \I__8164\ : Span12Mux_v
    port map (
            O => \N__38963\,
            I => \N__38955\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__38960\,
            I => \N__38955\
        );

    \I__8162\ : Odrv12
    port map (
            O => \N__38955\,
            I => \data_index_9_N_216_9\
        );

    \I__8161\ : InMux
    port map (
            O => \N__38952\,
            I => \N__38948\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38945\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38948\,
            I => n7_adj_1560
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__38945\,
            I => n7_adj_1560
        );

    \I__8157\ : CascadeMux
    port map (
            O => \N__38940\,
            I => \N__38937\
        );

    \I__8156\ : CascadeBuf
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__38934\,
            I => \N__38931\
        );

    \I__8154\ : CascadeBuf
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__38928\,
            I => \N__38925\
        );

    \I__8152\ : CascadeBuf
    port map (
            O => \N__38925\,
            I => \N__38922\
        );

    \I__8151\ : CascadeMux
    port map (
            O => \N__38922\,
            I => \N__38919\
        );

    \I__8150\ : CascadeBuf
    port map (
            O => \N__38919\,
            I => \N__38916\
        );

    \I__8149\ : CascadeMux
    port map (
            O => \N__38916\,
            I => \N__38913\
        );

    \I__8148\ : CascadeBuf
    port map (
            O => \N__38913\,
            I => \N__38910\
        );

    \I__8147\ : CascadeMux
    port map (
            O => \N__38910\,
            I => \N__38907\
        );

    \I__8146\ : CascadeBuf
    port map (
            O => \N__38907\,
            I => \N__38904\
        );

    \I__8145\ : CascadeMux
    port map (
            O => \N__38904\,
            I => \N__38901\
        );

    \I__8144\ : CascadeBuf
    port map (
            O => \N__38901\,
            I => \N__38897\
        );

    \I__8143\ : CascadeMux
    port map (
            O => \N__38900\,
            I => \N__38894\
        );

    \I__8142\ : CascadeMux
    port map (
            O => \N__38897\,
            I => \N__38891\
        );

    \I__8141\ : CascadeBuf
    port map (
            O => \N__38894\,
            I => \N__38888\
        );

    \I__8140\ : CascadeBuf
    port map (
            O => \N__38891\,
            I => \N__38885\
        );

    \I__8139\ : CascadeMux
    port map (
            O => \N__38888\,
            I => \N__38882\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__38885\,
            I => \N__38879\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38882\,
            I => \N__38876\
        );

    \I__8136\ : CascadeBuf
    port map (
            O => \N__38879\,
            I => \N__38873\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__38876\,
            I => \N__38870\
        );

    \I__8134\ : CascadeMux
    port map (
            O => \N__38873\,
            I => \N__38867\
        );

    \I__8133\ : Span12Mux_h
    port map (
            O => \N__38870\,
            I => \N__38864\
        );

    \I__8132\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38861\
        );

    \I__8131\ : Span12Mux_v
    port map (
            O => \N__38864\,
            I => \N__38856\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__38861\,
            I => \N__38856\
        );

    \I__8129\ : Odrv12
    port map (
            O => \N__38856\,
            I => \data_index_9_N_216_8\
        );

    \I__8128\ : CascadeMux
    port map (
            O => \N__38853\,
            I => \N__38850\
        );

    \I__8127\ : CascadeBuf
    port map (
            O => \N__38850\,
            I => \N__38847\
        );

    \I__8126\ : CascadeMux
    port map (
            O => \N__38847\,
            I => \N__38844\
        );

    \I__8125\ : CascadeBuf
    port map (
            O => \N__38844\,
            I => \N__38841\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__8123\ : CascadeBuf
    port map (
            O => \N__38838\,
            I => \N__38835\
        );

    \I__8122\ : CascadeMux
    port map (
            O => \N__38835\,
            I => \N__38832\
        );

    \I__8121\ : CascadeBuf
    port map (
            O => \N__38832\,
            I => \N__38829\
        );

    \I__8120\ : CascadeMux
    port map (
            O => \N__38829\,
            I => \N__38826\
        );

    \I__8119\ : CascadeBuf
    port map (
            O => \N__38826\,
            I => \N__38823\
        );

    \I__8118\ : CascadeMux
    port map (
            O => \N__38823\,
            I => \N__38820\
        );

    \I__8117\ : CascadeBuf
    port map (
            O => \N__38820\,
            I => \N__38817\
        );

    \I__8116\ : CascadeMux
    port map (
            O => \N__38817\,
            I => \N__38814\
        );

    \I__8115\ : CascadeBuf
    port map (
            O => \N__38814\,
            I => \N__38810\
        );

    \I__8114\ : CascadeMux
    port map (
            O => \N__38813\,
            I => \N__38807\
        );

    \I__8113\ : CascadeMux
    port map (
            O => \N__38810\,
            I => \N__38804\
        );

    \I__8112\ : CascadeBuf
    port map (
            O => \N__38807\,
            I => \N__38801\
        );

    \I__8111\ : CascadeBuf
    port map (
            O => \N__38804\,
            I => \N__38798\
        );

    \I__8110\ : CascadeMux
    port map (
            O => \N__38801\,
            I => \N__38795\
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__38798\,
            I => \N__38792\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38795\,
            I => \N__38789\
        );

    \I__8107\ : CascadeBuf
    port map (
            O => \N__38792\,
            I => \N__38786\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__38789\,
            I => \N__38783\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__38786\,
            I => \N__38780\
        );

    \I__8104\ : Span12Mux_h
    port map (
            O => \N__38783\,
            I => \N__38777\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38774\
        );

    \I__8102\ : Span12Mux_v
    port map (
            O => \N__38777\,
            I => \N__38769\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__38774\,
            I => \N__38769\
        );

    \I__8100\ : Odrv12
    port map (
            O => \N__38769\,
            I => \data_index_9_N_216_7\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38766\,
            I => \N__38762\
        );

    \I__8098\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38759\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__38762\,
            I => \N__38756\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__38759\,
            I => \N__38742\
        );

    \I__8095\ : Glb2LocalMux
    port map (
            O => \N__38756\,
            I => \N__38706\
        );

    \I__8094\ : ClkMux
    port map (
            O => \N__38755\,
            I => \N__38706\
        );

    \I__8093\ : ClkMux
    port map (
            O => \N__38754\,
            I => \N__38706\
        );

    \I__8092\ : ClkMux
    port map (
            O => \N__38753\,
            I => \N__38706\
        );

    \I__8091\ : ClkMux
    port map (
            O => \N__38752\,
            I => \N__38706\
        );

    \I__8090\ : ClkMux
    port map (
            O => \N__38751\,
            I => \N__38706\
        );

    \I__8089\ : ClkMux
    port map (
            O => \N__38750\,
            I => \N__38706\
        );

    \I__8088\ : ClkMux
    port map (
            O => \N__38749\,
            I => \N__38706\
        );

    \I__8087\ : ClkMux
    port map (
            O => \N__38748\,
            I => \N__38706\
        );

    \I__8086\ : ClkMux
    port map (
            O => \N__38747\,
            I => \N__38706\
        );

    \I__8085\ : ClkMux
    port map (
            O => \N__38746\,
            I => \N__38706\
        );

    \I__8084\ : ClkMux
    port map (
            O => \N__38745\,
            I => \N__38706\
        );

    \I__8083\ : Glb2LocalMux
    port map (
            O => \N__38742\,
            I => \N__38706\
        );

    \I__8082\ : ClkMux
    port map (
            O => \N__38741\,
            I => \N__38706\
        );

    \I__8081\ : ClkMux
    port map (
            O => \N__38740\,
            I => \N__38706\
        );

    \I__8080\ : ClkMux
    port map (
            O => \N__38739\,
            I => \N__38706\
        );

    \I__8079\ : GlobalMux
    port map (
            O => \N__38706\,
            I => \clk_16MHz\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38703\,
            I => \N__38700\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__38700\,
            I => \N__38697\
        );

    \I__8076\ : Span4Mux_v
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__8075\ : Span4Mux_v
    port map (
            O => \N__38694\,
            I => \N__38691\
        );

    \I__8074\ : Span4Mux_v
    port map (
            O => \N__38691\,
            I => \N__38687\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38684\
        );

    \I__8072\ : Odrv4
    port map (
            O => \N__38687\,
            I => dds0_mclk
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__38684\,
            I => dds0_mclk
        );

    \I__8070\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38676\,
            I => \N__38671\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__38675\,
            I => \N__38668\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38665\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__38671\,
            I => \N__38662\
        );

    \I__8065\ : InMux
    port map (
            O => \N__38668\,
            I => \N__38659\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__38665\,
            I => \N__38656\
        );

    \I__8063\ : Odrv4
    port map (
            O => \N__38662\,
            I => buf_control_6
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__38659\,
            I => buf_control_6
        );

    \I__8061\ : Odrv4
    port map (
            O => \N__38656\,
            I => buf_control_6
        );

    \I__8060\ : IoInMux
    port map (
            O => \N__38649\,
            I => \N__38646\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38646\,
            I => \N__38643\
        );

    \I__8058\ : Span4Mux_s2_v
    port map (
            O => \N__38643\,
            I => \N__38640\
        );

    \I__8057\ : Span4Mux_h
    port map (
            O => \N__38640\,
            I => \N__38637\
        );

    \I__8056\ : Span4Mux_h
    port map (
            O => \N__38637\,
            I => \N__38634\
        );

    \I__8055\ : Span4Mux_v
    port map (
            O => \N__38634\,
            I => \N__38631\
        );

    \I__8054\ : Odrv4
    port map (
            O => \N__38631\,
            I => \DDS_MCLK\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38628\,
            I => \N__38625\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__38625\,
            I => \N__38622\
        );

    \I__8051\ : Span4Mux_v
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__8050\ : Span4Mux_v
    port map (
            O => \N__38619\,
            I => \N__38615\
        );

    \I__8049\ : InMux
    port map (
            O => \N__38618\,
            I => \N__38612\
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__38615\,
            I => \comm_spi.n14619\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__38612\,
            I => \comm_spi.n14619\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38603\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38600\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__38603\,
            I => \comm_spi.n22884\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__38600\,
            I => \comm_spi.n22884\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__38595\,
            I => \comm_spi.n22884_cascade_\
        );

    \I__8041\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38588\
        );

    \I__8040\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38585\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__38588\,
            I => \comm_spi.n14593\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__38585\,
            I => \comm_spi.n14593\
        );

    \I__8037\ : InMux
    port map (
            O => \N__38580\,
            I => \N__38577\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__38577\,
            I => \N__38574\
        );

    \I__8035\ : Span4Mux_v
    port map (
            O => \N__38574\,
            I => \N__38570\
        );

    \I__8034\ : InMux
    port map (
            O => \N__38573\,
            I => \N__38567\
        );

    \I__8033\ : Span4Mux_v
    port map (
            O => \N__38570\,
            I => \N__38562\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__38567\,
            I => \N__38562\
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__38562\,
            I => \comm_spi.n14618\
        );

    \I__8030\ : CEMux
    port map (
            O => \N__38559\,
            I => \N__38553\
        );

    \I__8029\ : CEMux
    port map (
            O => \N__38558\,
            I => \N__38549\
        );

    \I__8028\ : CEMux
    port map (
            O => \N__38557\,
            I => \N__38546\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38543\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__38553\,
            I => \N__38540\
        );

    \I__8025\ : CEMux
    port map (
            O => \N__38552\,
            I => \N__38537\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__38549\,
            I => \N__38534\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__38546\,
            I => \N__38531\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__38543\,
            I => \N__38528\
        );

    \I__8021\ : Span4Mux_v
    port map (
            O => \N__38540\,
            I => \N__38525\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__38537\,
            I => \N__38522\
        );

    \I__8019\ : Span4Mux_h
    port map (
            O => \N__38534\,
            I => \N__38519\
        );

    \I__8018\ : Span4Mux_h
    port map (
            O => \N__38531\,
            I => \N__38516\
        );

    \I__8017\ : Span4Mux_h
    port map (
            O => \N__38528\,
            I => \N__38513\
        );

    \I__8016\ : Span4Mux_h
    port map (
            O => \N__38525\,
            I => \N__38508\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__38522\,
            I => \N__38508\
        );

    \I__8014\ : Span4Mux_v
    port map (
            O => \N__38519\,
            I => \N__38501\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__38516\,
            I => \N__38501\
        );

    \I__8012\ : Span4Mux_v
    port map (
            O => \N__38513\,
            I => \N__38501\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__38508\,
            I => n13457
        );

    \I__8010\ : Odrv4
    port map (
            O => \N__38501\,
            I => n13457
        );

    \I__8009\ : SRMux
    port map (
            O => \N__38496\,
            I => \N__38493\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__38493\,
            I => \N__38490\
        );

    \I__8007\ : Span4Mux_v
    port map (
            O => \N__38490\,
            I => \N__38486\
        );

    \I__8006\ : SRMux
    port map (
            O => \N__38489\,
            I => \N__38483\
        );

    \I__8005\ : Span4Mux_h
    port map (
            O => \N__38486\,
            I => \N__38476\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__38483\,
            I => \N__38476\
        );

    \I__8003\ : SRMux
    port map (
            O => \N__38482\,
            I => \N__38473\
        );

    \I__8002\ : SRMux
    port map (
            O => \N__38481\,
            I => \N__38470\
        );

    \I__8001\ : Span4Mux_v
    port map (
            O => \N__38476\,
            I => \N__38465\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N__38465\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__38470\,
            I => \N__38462\
        );

    \I__7998\ : Span4Mux_h
    port map (
            O => \N__38465\,
            I => \N__38459\
        );

    \I__7997\ : Span4Mux_v
    port map (
            O => \N__38462\,
            I => \N__38456\
        );

    \I__7996\ : Odrv4
    port map (
            O => \N__38459\,
            I => n14647
        );

    \I__7995\ : Odrv4
    port map (
            O => \N__38456\,
            I => n14647
        );

    \I__7994\ : CascadeMux
    port map (
            O => \N__38451\,
            I => \N__38447\
        );

    \I__7993\ : InMux
    port map (
            O => \N__38450\,
            I => \N__38444\
        );

    \I__7992\ : InMux
    port map (
            O => \N__38447\,
            I => \N__38441\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__38444\,
            I => \N__38438\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__38441\,
            I => acadc_skipcnt_0
        );

    \I__7989\ : Odrv12
    port map (
            O => \N__38438\,
            I => acadc_skipcnt_0
        );

    \I__7988\ : CascadeMux
    port map (
            O => \N__38433\,
            I => \N__38430\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38430\,
            I => \N__38427\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__38427\,
            I => \N__38423\
        );

    \I__7985\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38420\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__38423\,
            I => \N__38417\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__38420\,
            I => acadc_skipcnt_6
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__38417\,
            I => acadc_skipcnt_6
        );

    \I__7981\ : InMux
    port map (
            O => \N__38412\,
            I => \N__38409\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__38409\,
            I => \N__38406\
        );

    \I__7979\ : Span4Mux_v
    port map (
            O => \N__38406\,
            I => \N__38403\
        );

    \I__7978\ : Span4Mux_h
    port map (
            O => \N__38403\,
            I => \N__38400\
        );

    \I__7977\ : Odrv4
    port map (
            O => \N__38400\,
            I => n17
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__38397\,
            I => \n8_adj_1565_cascade_\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38394\,
            I => \N__38389\
        );

    \I__7974\ : InMux
    port map (
            O => \N__38393\,
            I => \N__38386\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38392\,
            I => \N__38383\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38389\,
            I => data_index_6
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__38386\,
            I => data_index_6
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__38383\,
            I => data_index_6
        );

    \I__7969\ : CascadeMux
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__7968\ : CascadeBuf
    port map (
            O => \N__38373\,
            I => \N__38370\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__38370\,
            I => \N__38367\
        );

    \I__7966\ : CascadeBuf
    port map (
            O => \N__38367\,
            I => \N__38364\
        );

    \I__7965\ : CascadeMux
    port map (
            O => \N__38364\,
            I => \N__38361\
        );

    \I__7964\ : CascadeBuf
    port map (
            O => \N__38361\,
            I => \N__38358\
        );

    \I__7963\ : CascadeMux
    port map (
            O => \N__38358\,
            I => \N__38355\
        );

    \I__7962\ : CascadeBuf
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__38352\,
            I => \N__38349\
        );

    \I__7960\ : CascadeBuf
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__38346\,
            I => \N__38343\
        );

    \I__7958\ : CascadeBuf
    port map (
            O => \N__38343\,
            I => \N__38340\
        );

    \I__7957\ : CascadeMux
    port map (
            O => \N__38340\,
            I => \N__38337\
        );

    \I__7956\ : CascadeBuf
    port map (
            O => \N__38337\,
            I => \N__38334\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__38334\,
            I => \N__38331\
        );

    \I__7954\ : CascadeBuf
    port map (
            O => \N__38331\,
            I => \N__38327\
        );

    \I__7953\ : CascadeMux
    port map (
            O => \N__38330\,
            I => \N__38324\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__38327\,
            I => \N__38321\
        );

    \I__7951\ : CascadeBuf
    port map (
            O => \N__38324\,
            I => \N__38318\
        );

    \I__7950\ : CascadeBuf
    port map (
            O => \N__38321\,
            I => \N__38315\
        );

    \I__7949\ : CascadeMux
    port map (
            O => \N__38318\,
            I => \N__38312\
        );

    \I__7948\ : CascadeMux
    port map (
            O => \N__38315\,
            I => \N__38309\
        );

    \I__7947\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38306\
        );

    \I__7946\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38303\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__38306\,
            I => \N__38300\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__38303\,
            I => \N__38297\
        );

    \I__7943\ : Sp12to4
    port map (
            O => \N__38300\,
            I => \N__38294\
        );

    \I__7942\ : Span4Mux_h
    port map (
            O => \N__38297\,
            I => \N__38291\
        );

    \I__7941\ : Span12Mux_v
    port map (
            O => \N__38294\,
            I => \N__38288\
        );

    \I__7940\ : Span4Mux_h
    port map (
            O => \N__38291\,
            I => \N__38285\
        );

    \I__7939\ : Odrv12
    port map (
            O => \N__38288\,
            I => \data_index_9_N_216_3\
        );

    \I__7938\ : Odrv4
    port map (
            O => \N__38285\,
            I => \data_index_9_N_216_3\
        );

    \I__7937\ : CascadeMux
    port map (
            O => \N__38280\,
            I => \N__38277\
        );

    \I__7936\ : InMux
    port map (
            O => \N__38277\,
            I => \N__38274\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__38274\,
            I => \N__38271\
        );

    \I__7934\ : Odrv4
    port map (
            O => \N__38271\,
            I => n8_adj_1565
        );

    \I__7933\ : InMux
    port map (
            O => \N__38268\,
            I => \N__38264\
        );

    \I__7932\ : InMux
    port map (
            O => \N__38267\,
            I => \N__38261\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__38264\,
            I => n7_adj_1564
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__38261\,
            I => n7_adj_1564
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__38256\,
            I => \N__38253\
        );

    \I__7928\ : CascadeBuf
    port map (
            O => \N__38253\,
            I => \N__38250\
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__38250\,
            I => \N__38247\
        );

    \I__7926\ : CascadeBuf
    port map (
            O => \N__38247\,
            I => \N__38244\
        );

    \I__7925\ : CascadeMux
    port map (
            O => \N__38244\,
            I => \N__38241\
        );

    \I__7924\ : CascadeBuf
    port map (
            O => \N__38241\,
            I => \N__38238\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__38238\,
            I => \N__38235\
        );

    \I__7922\ : CascadeBuf
    port map (
            O => \N__38235\,
            I => \N__38232\
        );

    \I__7921\ : CascadeMux
    port map (
            O => \N__38232\,
            I => \N__38229\
        );

    \I__7920\ : CascadeBuf
    port map (
            O => \N__38229\,
            I => \N__38226\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__7918\ : CascadeBuf
    port map (
            O => \N__38223\,
            I => \N__38220\
        );

    \I__7917\ : CascadeMux
    port map (
            O => \N__38220\,
            I => \N__38217\
        );

    \I__7916\ : CascadeBuf
    port map (
            O => \N__38217\,
            I => \N__38214\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__38214\,
            I => \N__38210\
        );

    \I__7914\ : CascadeMux
    port map (
            O => \N__38213\,
            I => \N__38207\
        );

    \I__7913\ : CascadeBuf
    port map (
            O => \N__38210\,
            I => \N__38204\
        );

    \I__7912\ : CascadeBuf
    port map (
            O => \N__38207\,
            I => \N__38201\
        );

    \I__7911\ : CascadeMux
    port map (
            O => \N__38204\,
            I => \N__38198\
        );

    \I__7910\ : CascadeMux
    port map (
            O => \N__38201\,
            I => \N__38195\
        );

    \I__7909\ : CascadeBuf
    port map (
            O => \N__38198\,
            I => \N__38192\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38195\,
            I => \N__38189\
        );

    \I__7907\ : CascadeMux
    port map (
            O => \N__38192\,
            I => \N__38186\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__38189\,
            I => \N__38183\
        );

    \I__7905\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38180\
        );

    \I__7904\ : Span12Mux_h
    port map (
            O => \N__38183\,
            I => \N__38177\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__38180\,
            I => \N__38174\
        );

    \I__7902\ : Span12Mux_v
    port map (
            O => \N__38177\,
            I => \N__38171\
        );

    \I__7901\ : Span4Mux_h
    port map (
            O => \N__38174\,
            I => \N__38168\
        );

    \I__7900\ : Odrv12
    port map (
            O => \N__38171\,
            I => \data_index_9_N_216_6\
        );

    \I__7899\ : Odrv4
    port map (
            O => \N__38168\,
            I => \data_index_9_N_216_6\
        );

    \I__7898\ : InMux
    port map (
            O => \N__38163\,
            I => n19601
        );

    \I__7897\ : InMux
    port map (
            O => \N__38160\,
            I => \bfn_15_17_0_\
        );

    \I__7896\ : InMux
    port map (
            O => \N__38157\,
            I => n19603
        );

    \I__7895\ : InMux
    port map (
            O => \N__38154\,
            I => n19604
        );

    \I__7894\ : InMux
    port map (
            O => \N__38151\,
            I => n19605
        );

    \I__7893\ : InMux
    port map (
            O => \N__38148\,
            I => \N__38145\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__38145\,
            I => \N__38141\
        );

    \I__7891\ : InMux
    port map (
            O => \N__38144\,
            I => \N__38138\
        );

    \I__7890\ : Span4Mux_h
    port map (
            O => \N__38141\,
            I => \N__38135\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__38138\,
            I => data_cntvec_12
        );

    \I__7888\ : Odrv4
    port map (
            O => \N__38135\,
            I => data_cntvec_12
        );

    \I__7887\ : InMux
    port map (
            O => \N__38130\,
            I => n19606
        );

    \I__7886\ : InMux
    port map (
            O => \N__38127\,
            I => \N__38124\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__38124\,
            I => \N__38120\
        );

    \I__7884\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38117\
        );

    \I__7883\ : Span4Mux_v
    port map (
            O => \N__38120\,
            I => \N__38114\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__38117\,
            I => data_cntvec_13
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__38114\,
            I => data_cntvec_13
        );

    \I__7880\ : InMux
    port map (
            O => \N__38109\,
            I => n19607
        );

    \I__7879\ : InMux
    port map (
            O => \N__38106\,
            I => \N__38102\
        );

    \I__7878\ : InMux
    port map (
            O => \N__38105\,
            I => \N__38099\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__38102\,
            I => data_cntvec_14
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__38099\,
            I => data_cntvec_14
        );

    \I__7875\ : InMux
    port map (
            O => \N__38094\,
            I => n19608
        );

    \I__7874\ : InMux
    port map (
            O => \N__38091\,
            I => n19609
        );

    \I__7873\ : InMux
    port map (
            O => \N__38088\,
            I => \N__38085\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__38085\,
            I => \N__38081\
        );

    \I__7871\ : InMux
    port map (
            O => \N__38084\,
            I => \N__38078\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__38081\,
            I => \N__38075\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__38078\,
            I => data_cntvec_15
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__38075\,
            I => data_cntvec_15
        );

    \I__7867\ : InMux
    port map (
            O => \N__38070\,
            I => \N__38066\
        );

    \I__7866\ : InMux
    port map (
            O => \N__38069\,
            I => \N__38063\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__38066\,
            I => \N__38058\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__38063\,
            I => \N__38058\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__38058\,
            I => \N__38055\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__38055\,
            I => \N__38052\
        );

    \I__7861\ : Odrv4
    port map (
            O => \N__38052\,
            I => n14_adj_1576
        );

    \I__7860\ : CascadeMux
    port map (
            O => \N__38049\,
            I => \N__38045\
        );

    \I__7859\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38042\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38045\,
            I => \N__38039\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__38042\,
            I => \N__38036\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__38039\,
            I => data_idxvec_14
        );

    \I__7855\ : Odrv12
    port map (
            O => \N__38036\,
            I => data_idxvec_14
        );

    \I__7854\ : InMux
    port map (
            O => \N__38031\,
            I => n19647
        );

    \I__7853\ : InMux
    port map (
            O => \N__38028\,
            I => \N__38025\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__38025\,
            I => \N__38022\
        );

    \I__7851\ : Span4Mux_v
    port map (
            O => \N__38022\,
            I => \N__38019\
        );

    \I__7850\ : Span4Mux_h
    port map (
            O => \N__38019\,
            I => \N__38015\
        );

    \I__7849\ : InMux
    port map (
            O => \N__38018\,
            I => \N__38012\
        );

    \I__7848\ : Odrv4
    port map (
            O => \N__38015\,
            I => n14_adj_1549
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__38012\,
            I => n14_adj_1549
        );

    \I__7846\ : InMux
    port map (
            O => \N__38007\,
            I => n19648
        );

    \I__7845\ : InMux
    port map (
            O => \N__38004\,
            I => \N__38001\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__38001\,
            I => \N__37997\
        );

    \I__7843\ : InMux
    port map (
            O => \N__38000\,
            I => \N__37994\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__37997\,
            I => \N__37991\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__37994\,
            I => data_idxvec_15
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__37991\,
            I => data_idxvec_15
        );

    \I__7839\ : CEMux
    port map (
            O => \N__37986\,
            I => \N__37983\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37979\
        );

    \I__7837\ : CEMux
    port map (
            O => \N__37982\,
            I => \N__37976\
        );

    \I__7836\ : Span4Mux_v
    port map (
            O => \N__37979\,
            I => \N__37971\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__37976\,
            I => \N__37971\
        );

    \I__7834\ : Span4Mux_v
    port map (
            O => \N__37971\,
            I => \N__37968\
        );

    \I__7833\ : Span4Mux_v
    port map (
            O => \N__37968\,
            I => \N__37965\
        );

    \I__7832\ : Odrv4
    port map (
            O => \N__37965\,
            I => n12280
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__37962\,
            I => \N__37959\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37959\,
            I => \N__37955\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37958\,
            I => \N__37950\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__37955\,
            I => \N__37947\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37954\,
            I => \N__37944\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37953\,
            I => \N__37941\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37950\,
            I => \N__37934\
        );

    \I__7824\ : Span4Mux_h
    port map (
            O => \N__37947\,
            I => \N__37934\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__37944\,
            I => \N__37934\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__37941\,
            I => \N__37931\
        );

    \I__7821\ : Span4Mux_v
    port map (
            O => \N__37934\,
            I => \N__37928\
        );

    \I__7820\ : Odrv4
    port map (
            O => \N__37931\,
            I => \iac_raw_buf_N_736\
        );

    \I__7819\ : Odrv4
    port map (
            O => \N__37928\,
            I => \iac_raw_buf_N_736\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37920\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37920\,
            I => \N__37915\
        );

    \I__7816\ : InMux
    port map (
            O => \N__37919\,
            I => \N__37912\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37909\
        );

    \I__7814\ : Span4Mux_v
    port map (
            O => \N__37915\,
            I => \N__37906\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37912\,
            I => data_cntvec_1
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__37909\,
            I => data_cntvec_1
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__37906\,
            I => data_cntvec_1
        );

    \I__7810\ : InMux
    port map (
            O => \N__37899\,
            I => n19595
        );

    \I__7809\ : InMux
    port map (
            O => \N__37896\,
            I => n19596
        );

    \I__7808\ : InMux
    port map (
            O => \N__37893\,
            I => n19597
        );

    \I__7807\ : InMux
    port map (
            O => \N__37890\,
            I => n19598
        );

    \I__7806\ : InMux
    port map (
            O => \N__37887\,
            I => n19599
        );

    \I__7805\ : InMux
    port map (
            O => \N__37884\,
            I => n19600
        );

    \I__7804\ : InMux
    port map (
            O => \N__37881\,
            I => n19639
        );

    \I__7803\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37874\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37871\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37874\,
            I => \N__37866\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__37871\,
            I => \N__37866\
        );

    \I__7799\ : Span4Mux_v
    port map (
            O => \N__37866\,
            I => \N__37863\
        );

    \I__7798\ : Span4Mux_h
    port map (
            O => \N__37863\,
            I => \N__37860\
        );

    \I__7797\ : Span4Mux_h
    port map (
            O => \N__37860\,
            I => \N__37857\
        );

    \I__7796\ : Odrv4
    port map (
            O => \N__37857\,
            I => n14_adj_1551
        );

    \I__7795\ : InMux
    port map (
            O => \N__37854\,
            I => n19640
        );

    \I__7794\ : InMux
    port map (
            O => \N__37851\,
            I => \N__37848\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__37848\,
            I => \N__37844\
        );

    \I__7792\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37841\
        );

    \I__7791\ : Span4Mux_h
    port map (
            O => \N__37844\,
            I => \N__37836\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__37841\,
            I => \N__37836\
        );

    \I__7789\ : Span4Mux_v
    port map (
            O => \N__37836\,
            I => \N__37833\
        );

    \I__7788\ : Odrv4
    port map (
            O => \N__37833\,
            I => n14_adj_1550
        );

    \I__7787\ : InMux
    port map (
            O => \N__37830\,
            I => \bfn_15_15_0_\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37827\,
            I => \N__37824\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__37824\,
            I => \N__37820\
        );

    \I__7784\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37817\
        );

    \I__7783\ : Span4Mux_v
    port map (
            O => \N__37820\,
            I => \N__37814\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__37817\,
            I => \N__37811\
        );

    \I__7781\ : Span4Mux_v
    port map (
            O => \N__37814\,
            I => \N__37808\
        );

    \I__7780\ : Sp12to4
    port map (
            O => \N__37811\,
            I => \N__37805\
        );

    \I__7779\ : Sp12to4
    port map (
            O => \N__37808\,
            I => \N__37800\
        );

    \I__7778\ : Span12Mux_v
    port map (
            O => \N__37805\,
            I => \N__37800\
        );

    \I__7777\ : Odrv12
    port map (
            O => \N__37800\,
            I => n14_adj_1580
        );

    \I__7776\ : InMux
    port map (
            O => \N__37797\,
            I => n19642
        );

    \I__7775\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37791\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37791\,
            I => \N__37787\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37784\
        );

    \I__7772\ : Span4Mux_v
    port map (
            O => \N__37787\,
            I => \N__37781\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37784\,
            I => n14_adj_1579
        );

    \I__7770\ : Odrv4
    port map (
            O => \N__37781\,
            I => n14_adj_1579
        );

    \I__7769\ : InMux
    port map (
            O => \N__37776\,
            I => n19643
        );

    \I__7768\ : InMux
    port map (
            O => \N__37773\,
            I => n19644
        );

    \I__7767\ : InMux
    port map (
            O => \N__37770\,
            I => \N__37766\
        );

    \I__7766\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37763\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__37766\,
            I => \N__37760\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37757\
        );

    \I__7763\ : Span4Mux_h
    port map (
            O => \N__37760\,
            I => \N__37754\
        );

    \I__7762\ : Odrv4
    port map (
            O => \N__37757\,
            I => n14_adj_1577
        );

    \I__7761\ : Odrv4
    port map (
            O => \N__37754\,
            I => n14_adj_1577
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__37749\,
            I => \N__37745\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37742\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37739\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37742\,
            I => \N__37736\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__37739\,
            I => data_idxvec_12
        );

    \I__7755\ : Odrv4
    port map (
            O => \N__37736\,
            I => data_idxvec_12
        );

    \I__7754\ : InMux
    port map (
            O => \N__37731\,
            I => n19645
        );

    \I__7753\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37724\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37727\,
            I => \N__37721\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__37724\,
            I => \N__37718\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__37721\,
            I => \N__37714\
        );

    \I__7749\ : Span4Mux_v
    port map (
            O => \N__37718\,
            I => \N__37711\
        );

    \I__7748\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37708\
        );

    \I__7747\ : Span4Mux_h
    port map (
            O => \N__37714\,
            I => \N__37705\
        );

    \I__7746\ : Odrv4
    port map (
            O => \N__37711\,
            I => n14_adj_1583
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__37708\,
            I => n14_adj_1583
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__37705\,
            I => n14_adj_1583
        );

    \I__7743\ : CascadeMux
    port map (
            O => \N__37698\,
            I => \N__37695\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37695\,
            I => \N__37691\
        );

    \I__7741\ : CascadeMux
    port map (
            O => \N__37694\,
            I => \N__37688\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__37691\,
            I => \N__37685\
        );

    \I__7739\ : InMux
    port map (
            O => \N__37688\,
            I => \N__37682\
        );

    \I__7738\ : Span4Mux_h
    port map (
            O => \N__37685\,
            I => \N__37679\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__37682\,
            I => data_idxvec_13
        );

    \I__7736\ : Odrv4
    port map (
            O => \N__37679\,
            I => data_idxvec_13
        );

    \I__7735\ : InMux
    port map (
            O => \N__37674\,
            I => n19646
        );

    \I__7734\ : CascadeMux
    port map (
            O => \N__37671\,
            I => \N__37668\
        );

    \I__7733\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37665\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__37665\,
            I => \N__37662\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__37662\,
            I => \N__37659\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__37659\,
            I => n26_adj_1644
        );

    \I__7729\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37653\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__37653\,
            I => \N__37649\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37646\
        );

    \I__7726\ : Span4Mux_h
    port map (
            O => \N__37649\,
            I => \N__37639\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__37646\,
            I => \N__37639\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37645\,
            I => \N__37636\
        );

    \I__7723\ : InMux
    port map (
            O => \N__37644\,
            I => \N__37633\
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__37639\,
            I => n20893
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__37636\,
            I => n20893
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__37633\,
            I => n20893
        );

    \I__7719\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37623\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__7717\ : Span4Mux_v
    port map (
            O => \N__37620\,
            I => \N__37617\
        );

    \I__7716\ : Odrv4
    port map (
            O => \N__37617\,
            I => n21521
        );

    \I__7715\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37610\
        );

    \I__7714\ : InMux
    port map (
            O => \N__37613\,
            I => \N__37607\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__37610\,
            I => n14_adj_1533
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__37607\,
            I => n14_adj_1533
        );

    \I__7711\ : InMux
    port map (
            O => \N__37602\,
            I => \bfn_15_14_0_\
        );

    \I__7710\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37596\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__37596\,
            I => \N__37593\
        );

    \I__7708\ : Span4Mux_v
    port map (
            O => \N__37593\,
            I => \N__37590\
        );

    \I__7707\ : Span4Mux_h
    port map (
            O => \N__37590\,
            I => \N__37586\
        );

    \I__7706\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37583\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__37586\,
            I => \N__37580\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__37583\,
            I => n14_adj_1556
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__37580\,
            I => n14_adj_1556
        );

    \I__7702\ : CascadeMux
    port map (
            O => \N__37575\,
            I => \N__37571\
        );

    \I__7701\ : CascadeMux
    port map (
            O => \N__37574\,
            I => \N__37568\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37571\,
            I => \N__37565\
        );

    \I__7699\ : InMux
    port map (
            O => \N__37568\,
            I => \N__37562\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__37565\,
            I => \N__37559\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__37562\,
            I => data_idxvec_1
        );

    \I__7696\ : Odrv4
    port map (
            O => \N__37559\,
            I => data_idxvec_1
        );

    \I__7695\ : InMux
    port map (
            O => \N__37554\,
            I => n19634
        );

    \I__7694\ : InMux
    port map (
            O => \N__37551\,
            I => \N__37548\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__37548\,
            I => \N__37544\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37541\
        );

    \I__7691\ : Span4Mux_h
    port map (
            O => \N__37544\,
            I => \N__37538\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__37541\,
            I => n14_adj_1555
        );

    \I__7689\ : Odrv4
    port map (
            O => \N__37538\,
            I => n14_adj_1555
        );

    \I__7688\ : InMux
    port map (
            O => \N__37533\,
            I => n19635
        );

    \I__7687\ : InMux
    port map (
            O => \N__37530\,
            I => n19636
        );

    \I__7686\ : InMux
    port map (
            O => \N__37527\,
            I => \N__37523\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37526\,
            I => \N__37520\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__37523\,
            I => \N__37517\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__37520\,
            I => \N__37514\
        );

    \I__7682\ : Span4Mux_h
    port map (
            O => \N__37517\,
            I => \N__37511\
        );

    \I__7681\ : Span12Mux_h
    port map (
            O => \N__37514\,
            I => \N__37508\
        );

    \I__7680\ : Span4Mux_h
    port map (
            O => \N__37511\,
            I => \N__37505\
        );

    \I__7679\ : Odrv12
    port map (
            O => \N__37508\,
            I => n14_adj_1553
        );

    \I__7678\ : Odrv4
    port map (
            O => \N__37505\,
            I => n14_adj_1553
        );

    \I__7677\ : InMux
    port map (
            O => \N__37500\,
            I => n19637
        );

    \I__7676\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37493\
        );

    \I__7675\ : CascadeMux
    port map (
            O => \N__37496\,
            I => \N__37490\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37493\,
            I => \N__37487\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37490\,
            I => \N__37483\
        );

    \I__7672\ : Span4Mux_v
    port map (
            O => \N__37487\,
            I => \N__37480\
        );

    \I__7671\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37477\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__37483\,
            I => n14_adj_1584
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__37480\,
            I => n14_adj_1584
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__37477\,
            I => n14_adj_1584
        );

    \I__7667\ : InMux
    port map (
            O => \N__37470\,
            I => n19638
        );

    \I__7666\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37464\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__37464\,
            I => n22264
        );

    \I__7664\ : CascadeMux
    port map (
            O => \N__37461\,
            I => \n22414_cascade_\
        );

    \I__7663\ : CascadeMux
    port map (
            O => \N__37458\,
            I => \n30_adj_1524_cascade_\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__37455\,
            I => \N__37452\
        );

    \I__7661\ : InMux
    port map (
            O => \N__37452\,
            I => \N__37449\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__37449\,
            I => \N__37444\
        );

    \I__7659\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37441\
        );

    \I__7658\ : InMux
    port map (
            O => \N__37447\,
            I => \N__37437\
        );

    \I__7657\ : Span4Mux_v
    port map (
            O => \N__37444\,
            I => \N__37432\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__37441\,
            I => \N__37432\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37428\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__37437\,
            I => \N__37425\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__37432\,
            I => \N__37421\
        );

    \I__7652\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37418\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__37428\,
            I => \N__37413\
        );

    \I__7650\ : Span4Mux_v
    port map (
            O => \N__37425\,
            I => \N__37413\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37410\
        );

    \I__7648\ : Sp12to4
    port map (
            O => \N__37421\,
            I => \N__37405\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__37418\,
            I => \N__37405\
        );

    \I__7646\ : Sp12to4
    port map (
            O => \N__37413\,
            I => \N__37400\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__37410\,
            I => \N__37400\
        );

    \I__7644\ : Span12Mux_h
    port map (
            O => \N__37405\,
            I => \N__37397\
        );

    \I__7643\ : Span12Mux_v
    port map (
            O => \N__37400\,
            I => \N__37394\
        );

    \I__7642\ : Odrv12
    port map (
            O => \N__37397\,
            I => comm_buf_1_1
        );

    \I__7641\ : Odrv12
    port map (
            O => \N__37394\,
            I => comm_buf_1_1
        );

    \I__7640\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37386\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__37386\,
            I => \N__37382\
        );

    \I__7638\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37379\
        );

    \I__7637\ : Span12Mux_v
    port map (
            O => \N__37382\,
            I => \N__37374\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__37379\,
            I => \N__37374\
        );

    \I__7635\ : Odrv12
    port map (
            O => \N__37374\,
            I => \comm_spi.n14623\
        );

    \I__7634\ : SRMux
    port map (
            O => \N__37371\,
            I => \N__37368\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__37368\,
            I => \N__37365\
        );

    \I__7632\ : Span4Mux_h
    port map (
            O => \N__37365\,
            I => \N__37362\
        );

    \I__7631\ : Odrv4
    port map (
            O => \N__37362\,
            I => \comm_spi.data_tx_7__N_770\
        );

    \I__7630\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37356\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__37356\,
            I => \N__37352\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37349\
        );

    \I__7627\ : Odrv12
    port map (
            O => \N__37352\,
            I => \comm_spi.n14622\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__37349\,
            I => \comm_spi.n14622\
        );

    \I__7625\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37340\
        );

    \I__7624\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37337\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__37340\,
            I => \N__37332\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37332\
        );

    \I__7621\ : Span4Mux_h
    port map (
            O => \N__37332\,
            I => \N__37329\
        );

    \I__7620\ : Span4Mux_v
    port map (
            O => \N__37329\,
            I => \N__37325\
        );

    \I__7619\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37322\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__37325\,
            I => \comm_spi.n22857\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__37322\,
            I => \comm_spi.n22857\
        );

    \I__7616\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37313\
        );

    \I__7615\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37310\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__37313\,
            I => \N__37304\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__37310\,
            I => \N__37301\
        );

    \I__7612\ : CascadeMux
    port map (
            O => \N__37309\,
            I => \N__37294\
        );

    \I__7611\ : InMux
    port map (
            O => \N__37308\,
            I => \N__37288\
        );

    \I__7610\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37285\
        );

    \I__7609\ : Span4Mux_h
    port map (
            O => \N__37304\,
            I => \N__37282\
        );

    \I__7608\ : Span4Mux_h
    port map (
            O => \N__37301\,
            I => \N__37279\
        );

    \I__7607\ : CascadeMux
    port map (
            O => \N__37300\,
            I => \N__37276\
        );

    \I__7606\ : CascadeMux
    port map (
            O => \N__37299\,
            I => \N__37273\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__37298\,
            I => \N__37269\
        );

    \I__7604\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37266\
        );

    \I__7603\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37263\
        );

    \I__7602\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37258\
        );

    \I__7601\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37258\
        );

    \I__7600\ : InMux
    port map (
            O => \N__37291\,
            I => \N__37255\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__37288\,
            I => \N__37250\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__37285\,
            I => \N__37250\
        );

    \I__7597\ : Span4Mux_v
    port map (
            O => \N__37282\,
            I => \N__37247\
        );

    \I__7596\ : Span4Mux_v
    port map (
            O => \N__37279\,
            I => \N__37244\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37235\
        );

    \I__7594\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37235\
        );

    \I__7593\ : InMux
    port map (
            O => \N__37272\,
            I => \N__37235\
        );

    \I__7592\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37235\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__37266\,
            I => eis_state_1
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__37263\,
            I => eis_state_1
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__37258\,
            I => eis_state_1
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__37255\,
            I => eis_state_1
        );

    \I__7587\ : Odrv4
    port map (
            O => \N__37250\,
            I => eis_state_1
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__37247\,
            I => eis_state_1
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__37244\,
            I => eis_state_1
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__37235\,
            I => eis_state_1
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__37218\,
            I => \n20937_cascade_\
        );

    \I__7582\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37212\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__37212\,
            I => n20939
        );

    \I__7580\ : InMux
    port map (
            O => \N__37209\,
            I => \N__37206\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__37206\,
            I => n19_adj_1522
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__37203\,
            I => \N__37200\
        );

    \I__7577\ : InMux
    port map (
            O => \N__37200\,
            I => \N__37197\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__37197\,
            I => \N__37194\
        );

    \I__7575\ : Span4Mux_h
    port map (
            O => \N__37194\,
            I => \N__37190\
        );

    \I__7574\ : CascadeMux
    port map (
            O => \N__37193\,
            I => \N__37187\
        );

    \I__7573\ : Span4Mux_h
    port map (
            O => \N__37190\,
            I => \N__37184\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37181\
        );

    \I__7571\ : Odrv4
    port map (
            O => \N__37184\,
            I => \buf_readRTD_1\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37181\,
            I => \buf_readRTD_1\
        );

    \I__7569\ : InMux
    port map (
            O => \N__37176\,
            I => \N__37173\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__37173\,
            I => \N__37169\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37172\,
            I => \N__37166\
        );

    \I__7566\ : Span4Mux_v
    port map (
            O => \N__37169\,
            I => \N__37163\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__37166\,
            I => \N__37160\
        );

    \I__7564\ : Span4Mux_h
    port map (
            O => \N__37163\,
            I => \N__37156\
        );

    \I__7563\ : Sp12to4
    port map (
            O => \N__37160\,
            I => \N__37153\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37159\,
            I => \N__37150\
        );

    \I__7561\ : Sp12to4
    port map (
            O => \N__37156\,
            I => \N__37145\
        );

    \I__7560\ : Span12Mux_v
    port map (
            O => \N__37153\,
            I => \N__37145\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__37150\,
            I => buf_adcdata_iac_9
        );

    \I__7558\ : Odrv12
    port map (
            O => \N__37145\,
            I => buf_adcdata_iac_9
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__37140\,
            I => \n22261_cascade_\
        );

    \I__7556\ : InMux
    port map (
            O => \N__37137\,
            I => \N__37134\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__37134\,
            I => \N__37131\
        );

    \I__7554\ : Span4Mux_v
    port map (
            O => \N__37131\,
            I => \N__37128\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__37128\,
            I => n16_adj_1521
        );

    \I__7552\ : CascadeMux
    port map (
            O => \N__37125\,
            I => \n26_adj_1523_cascade_\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37122\,
            I => \N__37119\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__37119\,
            I => \N__37116\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__37116\,
            I => \N__37112\
        );

    \I__7548\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37108\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__37112\,
            I => \N__37105\
        );

    \I__7546\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37102\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__37108\,
            I => \acadc_skipCount_1\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__37105\,
            I => \acadc_skipCount_1\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__37102\,
            I => \acadc_skipCount_1\
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__37095\,
            I => \n22411_cascade_\
        );

    \I__7541\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37089\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37089\,
            I => \N__37086\
        );

    \I__7539\ : Span4Mux_v
    port map (
            O => \N__37086\,
            I => \N__37082\
        );

    \I__7538\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37078\
        );

    \I__7537\ : Span4Mux_v
    port map (
            O => \N__37082\,
            I => \N__37075\
        );

    \I__7536\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37072\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__37078\,
            I => req_data_cnt_1
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__37075\,
            I => req_data_cnt_1
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__37072\,
            I => req_data_cnt_1
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__37065\,
            I => \n21370_cascade_\
        );

    \I__7531\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37059\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__37059\,
            I => n21369
        );

    \I__7529\ : InMux
    port map (
            O => \N__37056\,
            I => \N__37053\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__37053\,
            I => n22426
        );

    \I__7527\ : CEMux
    port map (
            O => \N__37050\,
            I => \N__37047\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__37047\,
            I => \N__37044\
        );

    \I__7525\ : Sp12to4
    port map (
            O => \N__37044\,
            I => \N__37041\
        );

    \I__7524\ : Odrv12
    port map (
            O => \N__37041\,
            I => n14
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__37038\,
            I => \n1264_cascade_\
        );

    \I__7522\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37032\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__37032\,
            I => n4_adj_1643
        );

    \I__7520\ : InMux
    port map (
            O => \N__37029\,
            I => \N__37025\
        );

    \I__7519\ : InMux
    port map (
            O => \N__37028\,
            I => \N__37022\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__37025\,
            I => n1264
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__37022\,
            I => n1264
        );

    \I__7516\ : InMux
    port map (
            O => \N__37017\,
            I => \N__37014\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__37014\,
            I => n8_adj_1582
        );

    \I__7514\ : CascadeMux
    port map (
            O => \N__37011\,
            I => \N__37008\
        );

    \I__7513\ : InMux
    port map (
            O => \N__37008\,
            I => \N__37005\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__37005\,
            I => \comm_state_3_N_420_3\
        );

    \I__7511\ : CascadeMux
    port map (
            O => \N__37002\,
            I => \comm_state_3_N_420_3_cascade_\
        );

    \I__7510\ : CascadeMux
    port map (
            O => \N__36999\,
            I => \n21435_cascade_\
        );

    \I__7509\ : CEMux
    port map (
            O => \N__36996\,
            I => \N__36993\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__36993\,
            I => \N__36990\
        );

    \I__7507\ : Span4Mux_h
    port map (
            O => \N__36990\,
            I => \N__36987\
        );

    \I__7506\ : Odrv4
    port map (
            O => \N__36987\,
            I => n20829
        );

    \I__7505\ : CascadeMux
    port map (
            O => \N__36984\,
            I => \n20944_cascade_\
        );

    \I__7504\ : CEMux
    port map (
            O => \N__36981\,
            I => \N__36978\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__36978\,
            I => n20964
        );

    \I__7502\ : InMux
    port map (
            O => \N__36975\,
            I => \N__36972\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__36972\,
            I => n20962
        );

    \I__7500\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36963\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36963\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36963\,
            I => \N__36960\
        );

    \I__7497\ : Span12Mux_v
    port map (
            O => \N__36960\,
            I => \N__36957\
        );

    \I__7496\ : Odrv12
    port map (
            O => \N__36957\,
            I => n3
        );

    \I__7495\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36951\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__36951\,
            I => n20801
        );

    \I__7493\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36945\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36945\,
            I => n4_adj_1586
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__36942\,
            I => \n20801_cascade_\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36936\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__36936\,
            I => n19902
        );

    \I__7488\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36930\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__36930\,
            I => \N__36927\
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__36927\,
            I => n22423
        );

    \I__7485\ : CascadeMux
    port map (
            O => \N__36924\,
            I => \n2_adj_1581_cascade_\
        );

    \I__7484\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36914\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36920\,
            I => \N__36914\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36909\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__36914\,
            I => \N__36906\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36903\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36900\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__36909\,
            I => \N__36897\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__36906\,
            I => \N__36894\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36903\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__36900\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__36897\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__7473\ : Odrv4
    port map (
            O => \N__36894\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36885\,
            I => \ADC_VDC.n19775\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__36882\,
            I => \N__36876\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36873\
        );

    \I__7469\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36868\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36868\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36865\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__36873\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__36868\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__36865\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36858\,
            I => \ADC_VDC.n19776\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36849\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36844\
        );

    \I__7460\ : InMux
    port map (
            O => \N__36853\,
            I => \N__36844\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36852\,
            I => \N__36841\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36849\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__36844\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__36841\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__7455\ : InMux
    port map (
            O => \N__36834\,
            I => \ADC_VDC.n19777\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36831\,
            I => \ADC_VDC.n19778\
        );

    \I__7453\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36822\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36827\,
            I => \N__36819\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36816\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36825\,
            I => \N__36813\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__36822\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__36819\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__36816\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__36813\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__7445\ : SRMux
    port map (
            O => \N__36804\,
            I => \N__36801\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36801\,
            I => \N__36798\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__36798\,
            I => \ADC_VDC.n18550\
        );

    \I__7442\ : SRMux
    port map (
            O => \N__36795\,
            I => \N__36792\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__36792\,
            I => \N__36789\
        );

    \I__7440\ : Span4Mux_h
    port map (
            O => \N__36789\,
            I => \N__36786\
        );

    \I__7439\ : Span4Mux_v
    port map (
            O => \N__36786\,
            I => \N__36783\
        );

    \I__7438\ : Odrv4
    port map (
            O => \N__36783\,
            I => \comm_spi.data_tx_7__N_786\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36780\,
            I => \N__36777\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36777\,
            I => \N__36774\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__36774\,
            I => \N__36770\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36773\,
            I => \N__36767\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__36770\,
            I => tmp_buf_15
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__36767\,
            I => tmp_buf_15
        );

    \I__7431\ : IoInMux
    port map (
            O => \N__36762\,
            I => \N__36759\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36759\,
            I => \N__36756\
        );

    \I__7429\ : Span12Mux_s1_v
    port map (
            O => \N__36756\,
            I => \N__36753\
        );

    \I__7428\ : Span12Mux_h
    port map (
            O => \N__36753\,
            I => \N__36749\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36746\
        );

    \I__7426\ : Odrv12
    port map (
            O => \N__36749\,
            I => \DDS_MOSI\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36746\,
            I => \DDS_MOSI\
        );

    \I__7424\ : IoInMux
    port map (
            O => \N__36741\,
            I => \N__36738\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__36738\,
            I => \N__36735\
        );

    \I__7422\ : Span4Mux_s2_v
    port map (
            O => \N__36735\,
            I => \N__36732\
        );

    \I__7421\ : Span4Mux_h
    port map (
            O => \N__36732\,
            I => \N__36729\
        );

    \I__7420\ : Span4Mux_v
    port map (
            O => \N__36729\,
            I => \N__36726\
        );

    \I__7419\ : Sp12to4
    port map (
            O => \N__36726\,
            I => \N__36723\
        );

    \I__7418\ : Odrv12
    port map (
            O => \N__36723\,
            I => \DDS_CS\
        );

    \I__7417\ : CEMux
    port map (
            O => \N__36720\,
            I => \N__36717\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__36717\,
            I => \SIG_DDS.n9_adj_1393\
        );

    \I__7415\ : SRMux
    port map (
            O => \N__36714\,
            I => \N__36711\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__36711\,
            I => \comm_spi.data_tx_7__N_795\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36701\
        );

    \I__7412\ : CascadeMux
    port map (
            O => \N__36707\,
            I => \N__36698\
        );

    \I__7411\ : CascadeMux
    port map (
            O => \N__36706\,
            I => \N__36695\
        );

    \I__7410\ : InMux
    port map (
            O => \N__36705\,
            I => \N__36692\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36689\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36686\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36681\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36695\,
            I => \N__36681\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__36692\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__36689\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__36686\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__36681\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36672\,
            I => \bfn_15_4_0_\
        );

    \I__7400\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36663\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36668\,
            I => \N__36658\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36658\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36655\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__36663\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__36658\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__36655\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36648\,
            I => \ADC_VDC.n19772\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36641\
        );

    \I__7391\ : InMux
    port map (
            O => \N__36644\,
            I => \N__36635\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__36641\,
            I => \N__36632\
        );

    \I__7389\ : InMux
    port map (
            O => \N__36640\,
            I => \N__36629\
        );

    \I__7388\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36624\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36624\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__36635\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__36632\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__36629\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__36624\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__7382\ : InMux
    port map (
            O => \N__36615\,
            I => \ADC_VDC.n19773\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36605\
        );

    \I__7380\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36605\
        );

    \I__7379\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36600\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36597\
        );

    \I__7377\ : InMux
    port map (
            O => \N__36604\,
            I => \N__36594\
        );

    \I__7376\ : InMux
    port map (
            O => \N__36603\,
            I => \N__36591\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__36600\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__7374\ : Odrv4
    port map (
            O => \N__36597\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__36594\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__36591\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__7371\ : InMux
    port map (
            O => \N__36582\,
            I => \ADC_VDC.n19774\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36579\,
            I => n19629
        );

    \I__7369\ : InMux
    port map (
            O => \N__36576\,
            I => n19630
        );

    \I__7368\ : InMux
    port map (
            O => \N__36573\,
            I => n19631
        );

    \I__7367\ : InMux
    port map (
            O => \N__36570\,
            I => \bfn_14_19_0_\
        );

    \I__7366\ : CascadeMux
    port map (
            O => \N__36567\,
            I => \N__36563\
        );

    \I__7365\ : CascadeMux
    port map (
            O => \N__36566\,
            I => \N__36555\
        );

    \I__7364\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36552\
        );

    \I__7363\ : CascadeMux
    port map (
            O => \N__36562\,
            I => \N__36549\
        );

    \I__7362\ : CascadeMux
    port map (
            O => \N__36561\,
            I => \N__36546\
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__36560\,
            I => \N__36543\
        );

    \I__7360\ : CascadeMux
    port map (
            O => \N__36559\,
            I => \N__36540\
        );

    \I__7359\ : CascadeMux
    port map (
            O => \N__36558\,
            I => \N__36533\
        );

    \I__7358\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36530\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__36552\,
            I => \N__36527\
        );

    \I__7356\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36518\
        );

    \I__7355\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36518\
        );

    \I__7354\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36518\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36518\
        );

    \I__7352\ : CascadeMux
    port map (
            O => \N__36539\,
            I => \N__36515\
        );

    \I__7351\ : CascadeMux
    port map (
            O => \N__36538\,
            I => \N__36512\
        );

    \I__7350\ : CascadeMux
    port map (
            O => \N__36537\,
            I => \N__36509\
        );

    \I__7349\ : CascadeMux
    port map (
            O => \N__36536\,
            I => \N__36506\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36533\,
            I => \N__36503\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__36530\,
            I => \N__36496\
        );

    \I__7346\ : Span4Mux_h
    port map (
            O => \N__36527\,
            I => \N__36496\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36496\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36515\,
            I => \N__36487\
        );

    \I__7343\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36487\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36509\,
            I => \N__36487\
        );

    \I__7341\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36487\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__36503\,
            I => n10598
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__36496\,
            I => n10598
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__36487\,
            I => n10598
        );

    \I__7337\ : InMux
    port map (
            O => \N__36480\,
            I => n19633
        );

    \I__7336\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36473\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36470\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__36473\,
            I => n7_adj_1572
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36470\,
            I => n7_adj_1572
        );

    \I__7332\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36462\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__36462\,
            I => n8_adj_1573
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__36459\,
            I => \N__36456\
        );

    \I__7329\ : CascadeBuf
    port map (
            O => \N__36456\,
            I => \N__36453\
        );

    \I__7328\ : CascadeMux
    port map (
            O => \N__36453\,
            I => \N__36450\
        );

    \I__7327\ : CascadeBuf
    port map (
            O => \N__36450\,
            I => \N__36447\
        );

    \I__7326\ : CascadeMux
    port map (
            O => \N__36447\,
            I => \N__36444\
        );

    \I__7325\ : CascadeBuf
    port map (
            O => \N__36444\,
            I => \N__36441\
        );

    \I__7324\ : CascadeMux
    port map (
            O => \N__36441\,
            I => \N__36438\
        );

    \I__7323\ : CascadeBuf
    port map (
            O => \N__36438\,
            I => \N__36435\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__7321\ : CascadeBuf
    port map (
            O => \N__36432\,
            I => \N__36429\
        );

    \I__7320\ : CascadeMux
    port map (
            O => \N__36429\,
            I => \N__36426\
        );

    \I__7319\ : CascadeBuf
    port map (
            O => \N__36426\,
            I => \N__36423\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__36423\,
            I => \N__36420\
        );

    \I__7317\ : CascadeBuf
    port map (
            O => \N__36420\,
            I => \N__36417\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__36417\,
            I => \N__36413\
        );

    \I__7315\ : CascadeMux
    port map (
            O => \N__36416\,
            I => \N__36410\
        );

    \I__7314\ : CascadeBuf
    port map (
            O => \N__36413\,
            I => \N__36407\
        );

    \I__7313\ : CascadeBuf
    port map (
            O => \N__36410\,
            I => \N__36404\
        );

    \I__7312\ : CascadeMux
    port map (
            O => \N__36407\,
            I => \N__36401\
        );

    \I__7311\ : CascadeMux
    port map (
            O => \N__36404\,
            I => \N__36398\
        );

    \I__7310\ : CascadeBuf
    port map (
            O => \N__36401\,
            I => \N__36395\
        );

    \I__7309\ : InMux
    port map (
            O => \N__36398\,
            I => \N__36392\
        );

    \I__7308\ : CascadeMux
    port map (
            O => \N__36395\,
            I => \N__36389\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__36392\,
            I => \N__36386\
        );

    \I__7306\ : InMux
    port map (
            O => \N__36389\,
            I => \N__36383\
        );

    \I__7305\ : Span12Mux_h
    port map (
            O => \N__36386\,
            I => \N__36380\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__36383\,
            I => \N__36377\
        );

    \I__7303\ : Span12Mux_v
    port map (
            O => \N__36380\,
            I => \N__36374\
        );

    \I__7302\ : Span4Mux_h
    port map (
            O => \N__36377\,
            I => \N__36371\
        );

    \I__7301\ : Odrv12
    port map (
            O => \N__36374\,
            I => \data_index_9_N_216_1\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__36371\,
            I => \data_index_9_N_216_1\
        );

    \I__7299\ : CascadeMux
    port map (
            O => \N__36366\,
            I => \N__36362\
        );

    \I__7298\ : IoInMux
    port map (
            O => \N__36365\,
            I => \N__36359\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36356\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36359\,
            I => \N__36353\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__36356\,
            I => \N__36349\
        );

    \I__7294\ : Span12Mux_s7_v
    port map (
            O => \N__36353\,
            I => \N__36346\
        );

    \I__7293\ : InMux
    port map (
            O => \N__36352\,
            I => \N__36343\
        );

    \I__7292\ : Span4Mux_h
    port map (
            O => \N__36349\,
            I => \N__36340\
        );

    \I__7291\ : Odrv12
    port map (
            O => \N__36346\,
            I => \DDS_RNG_0\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__36343\,
            I => \DDS_RNG_0\
        );

    \I__7289\ : Odrv4
    port map (
            O => \N__36340\,
            I => \DDS_RNG_0\
        );

    \I__7288\ : InMux
    port map (
            O => \N__36333\,
            I => \N__36330\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__36330\,
            I => n11338
        );

    \I__7286\ : CascadeMux
    port map (
            O => \N__36327\,
            I => \n11338_cascade_\
        );

    \I__7285\ : CascadeMux
    port map (
            O => \N__36324\,
            I => \n8813_cascade_\
        );

    \I__7284\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36316\
        );

    \I__7283\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36313\
        );

    \I__7282\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36310\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__36316\,
            I => data_index_0
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__36313\,
            I => data_index_0
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__36310\,
            I => data_index_0
        );

    \I__7278\ : InMux
    port map (
            O => \N__36303\,
            I => \N__36297\
        );

    \I__7277\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36297\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__36297\,
            I => \N__36294\
        );

    \I__7275\ : Odrv12
    port map (
            O => \N__36294\,
            I => n7
        );

    \I__7274\ : InMux
    port map (
            O => \N__36291\,
            I => \bfn_14_18_0_\
        );

    \I__7273\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36283\
        );

    \I__7272\ : InMux
    port map (
            O => \N__36287\,
            I => \N__36280\
        );

    \I__7271\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36277\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__36283\,
            I => data_index_1
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36280\,
            I => data_index_1
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__36277\,
            I => data_index_1
        );

    \I__7267\ : InMux
    port map (
            O => \N__36270\,
            I => n19625
        );

    \I__7266\ : InMux
    port map (
            O => \N__36267\,
            I => n19626
        );

    \I__7265\ : InMux
    port map (
            O => \N__36264\,
            I => n19627
        );

    \I__7264\ : InMux
    port map (
            O => \N__36261\,
            I => n19628
        );

    \I__7263\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36255\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__36255\,
            I => \N__36251\
        );

    \I__7261\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36248\
        );

    \I__7260\ : Span4Mux_v
    port map (
            O => \N__36251\,
            I => \N__36244\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__36248\,
            I => \N__36241\
        );

    \I__7258\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36238\
        );

    \I__7257\ : Odrv4
    port map (
            O => \N__36244\,
            I => n10520
        );

    \I__7256\ : Odrv12
    port map (
            O => \N__36241\,
            I => n10520
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__36238\,
            I => n10520
        );

    \I__7254\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36227\
        );

    \I__7253\ : CascadeMux
    port map (
            O => \N__36230\,
            I => \N__36224\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__36227\,
            I => \N__36220\
        );

    \I__7251\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36217\
        );

    \I__7250\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36214\
        );

    \I__7249\ : Span4Mux_h
    port map (
            O => \N__36220\,
            I => \N__36209\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__36217\,
            I => \N__36209\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36214\,
            I => req_data_cnt_15
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__36209\,
            I => req_data_cnt_15
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__36204\,
            I => \n8_adj_1532_cascade_\
        );

    \I__7244\ : CascadeMux
    port map (
            O => \N__36201\,
            I => \N__36198\
        );

    \I__7243\ : CascadeBuf
    port map (
            O => \N__36198\,
            I => \N__36195\
        );

    \I__7242\ : CascadeMux
    port map (
            O => \N__36195\,
            I => \N__36192\
        );

    \I__7241\ : CascadeBuf
    port map (
            O => \N__36192\,
            I => \N__36189\
        );

    \I__7240\ : CascadeMux
    port map (
            O => \N__36189\,
            I => \N__36186\
        );

    \I__7239\ : CascadeBuf
    port map (
            O => \N__36186\,
            I => \N__36183\
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__36183\,
            I => \N__36180\
        );

    \I__7237\ : CascadeBuf
    port map (
            O => \N__36180\,
            I => \N__36177\
        );

    \I__7236\ : CascadeMux
    port map (
            O => \N__36177\,
            I => \N__36174\
        );

    \I__7235\ : CascadeBuf
    port map (
            O => \N__36174\,
            I => \N__36171\
        );

    \I__7234\ : CascadeMux
    port map (
            O => \N__36171\,
            I => \N__36168\
        );

    \I__7233\ : CascadeBuf
    port map (
            O => \N__36168\,
            I => \N__36165\
        );

    \I__7232\ : CascadeMux
    port map (
            O => \N__36165\,
            I => \N__36162\
        );

    \I__7231\ : CascadeBuf
    port map (
            O => \N__36162\,
            I => \N__36159\
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__36159\,
            I => \N__36155\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__36158\,
            I => \N__36152\
        );

    \I__7228\ : CascadeBuf
    port map (
            O => \N__36155\,
            I => \N__36149\
        );

    \I__7227\ : CascadeBuf
    port map (
            O => \N__36152\,
            I => \N__36146\
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__36149\,
            I => \N__36143\
        );

    \I__7225\ : CascadeMux
    port map (
            O => \N__36146\,
            I => \N__36140\
        );

    \I__7224\ : CascadeBuf
    port map (
            O => \N__36143\,
            I => \N__36137\
        );

    \I__7223\ : InMux
    port map (
            O => \N__36140\,
            I => \N__36134\
        );

    \I__7222\ : CascadeMux
    port map (
            O => \N__36137\,
            I => \N__36131\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__36134\,
            I => \N__36128\
        );

    \I__7220\ : InMux
    port map (
            O => \N__36131\,
            I => \N__36125\
        );

    \I__7219\ : Span4Mux_h
    port map (
            O => \N__36128\,
            I => \N__36122\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__36125\,
            I => \N__36119\
        );

    \I__7217\ : Sp12to4
    port map (
            O => \N__36122\,
            I => \N__36116\
        );

    \I__7216\ : Span4Mux_v
    port map (
            O => \N__36119\,
            I => \N__36113\
        );

    \I__7215\ : Span12Mux_v
    port map (
            O => \N__36116\,
            I => \N__36110\
        );

    \I__7214\ : Span4Mux_h
    port map (
            O => \N__36113\,
            I => \N__36107\
        );

    \I__7213\ : Odrv12
    port map (
            O => \N__36110\,
            I => \data_index_9_N_216_0\
        );

    \I__7212\ : Odrv4
    port map (
            O => \N__36107\,
            I => \data_index_9_N_216_0\
        );

    \I__7211\ : InMux
    port map (
            O => \N__36102\,
            I => \N__36099\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__36099\,
            I => n8_adj_1532
        );

    \I__7209\ : CEMux
    port map (
            O => \N__36096\,
            I => \N__36093\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__36093\,
            I => \N__36089\
        );

    \I__7207\ : CEMux
    port map (
            O => \N__36092\,
            I => \N__36086\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__36089\,
            I => \N__36083\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__36086\,
            I => \N__36080\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__36083\,
            I => \N__36075\
        );

    \I__7203\ : Span4Mux_h
    port map (
            O => \N__36080\,
            I => \N__36075\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__36075\,
            I => \SIG_DDS.n9\
        );

    \I__7201\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36069\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__36069\,
            I => n22_adj_1499
        );

    \I__7199\ : InMux
    port map (
            O => \N__36066\,
            I => \N__36063\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__36063\,
            I => n18
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__36060\,
            I => \N__36057\
        );

    \I__7196\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36052\
        );

    \I__7195\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36047\
        );

    \I__7194\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36047\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__36052\,
            I => \N__36044\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__36047\,
            I => req_data_cnt_14
        );

    \I__7191\ : Odrv4
    port map (
            O => \N__36044\,
            I => req_data_cnt_14
        );

    \I__7190\ : InMux
    port map (
            O => \N__36039\,
            I => \N__36036\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__36036\,
            I => n23_adj_1614
        );

    \I__7188\ : CascadeMux
    port map (
            O => \N__36033\,
            I => \n10_adj_1554_cascade_\
        );

    \I__7187\ : CEMux
    port map (
            O => \N__36030\,
            I => \N__36027\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__36027\,
            I => \N__36024\
        );

    \I__7185\ : Span4Mux_v
    port map (
            O => \N__36024\,
            I => \N__36021\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__36021\,
            I => n11850
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__36018\,
            I => \n20914_cascade_\
        );

    \I__7182\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36012\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__36012\,
            I => n21014
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__36009\,
            I => \N__36006\
        );

    \I__7179\ : InMux
    port map (
            O => \N__36006\,
            I => \N__36003\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__36003\,
            I => n17_adj_1489
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__36000\,
            I => \n16891_cascade_\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35994\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__35994\,
            I => \N__35991\
        );

    \I__7174\ : Span4Mux_v
    port map (
            O => \N__35991\,
            I => \N__35988\
        );

    \I__7173\ : Span4Mux_h
    port map (
            O => \N__35988\,
            I => \N__35985\
        );

    \I__7172\ : Odrv4
    port map (
            O => \N__35985\,
            I => \SIG_DDS.n21571\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35979\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35979\,
            I => \N__35976\
        );

    \I__7169\ : Span4Mux_v
    port map (
            O => \N__35976\,
            I => \N__35973\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__35973\,
            I => \N__35969\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35966\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__35969\,
            I => buf_adcdata_vdc_10
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35966\,
            I => buf_adcdata_vdc_10
        );

    \I__7164\ : InMux
    port map (
            O => \N__35961\,
            I => \N__35958\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__35958\,
            I => \N__35955\
        );

    \I__7162\ : Span4Mux_v
    port map (
            O => \N__35955\,
            I => \N__35951\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__35954\,
            I => \N__35948\
        );

    \I__7160\ : Span4Mux_h
    port map (
            O => \N__35951\,
            I => \N__35944\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35948\,
            I => \N__35941\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35947\,
            I => \N__35938\
        );

    \I__7157\ : Span4Mux_h
    port map (
            O => \N__35944\,
            I => \N__35935\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__35941\,
            I => buf_adcdata_vac_10
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__35938\,
            I => buf_adcdata_vac_10
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__35935\,
            I => buf_adcdata_vac_10
        );

    \I__7153\ : IoInMux
    port map (
            O => \N__35928\,
            I => \N__35925\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35925\,
            I => \N__35922\
        );

    \I__7151\ : Span4Mux_s2_h
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__7150\ : Sp12to4
    port map (
            O => \N__35919\,
            I => \N__35916\
        );

    \I__7149\ : Span12Mux_v
    port map (
            O => \N__35916\,
            I => \N__35913\
        );

    \I__7148\ : Span12Mux_h
    port map (
            O => \N__35913\,
            I => \N__35910\
        );

    \I__7147\ : Odrv12
    port map (
            O => \N__35910\,
            I => \ICE_GPMI_0\
        );

    \I__7146\ : CEMux
    port map (
            O => \N__35907\,
            I => \N__35904\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35904\,
            I => \N__35901\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__35901\,
            I => n11385
        );

    \I__7143\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35895\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__35895\,
            I => \N__35885\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35894\,
            I => \N__35869\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35893\,
            I => \N__35869\
        );

    \I__7139\ : InMux
    port map (
            O => \N__35892\,
            I => \N__35869\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35869\
        );

    \I__7137\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35869\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35869\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35869\
        );

    \I__7134\ : Span4Mux_v
    port map (
            O => \N__35885\,
            I => \N__35866\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35863\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__35869\,
            I => \N__35860\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__35866\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35863\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__35860\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35850\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__35850\,
            I => \N__35847\
        );

    \I__7126\ : Span4Mux_v
    port map (
            O => \N__35847\,
            I => \N__35837\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35822\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35822\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35822\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35822\
        );

    \I__7121\ : InMux
    port map (
            O => \N__35842\,
            I => \N__35822\
        );

    \I__7120\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35822\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35822\
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__35837\,
            I => \comm_spi.n17036\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35822\,
            I => \comm_spi.n17036\
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__35817\,
            I => \N__35812\
        );

    \I__7115\ : CascadeMux
    port map (
            O => \N__35816\,
            I => \N__35809\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35815\,
            I => \N__35799\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35792\
        );

    \I__7112\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35792\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35808\,
            I => \N__35789\
        );

    \I__7110\ : InMux
    port map (
            O => \N__35807\,
            I => \N__35786\
        );

    \I__7109\ : InMux
    port map (
            O => \N__35806\,
            I => \N__35783\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35805\,
            I => \N__35780\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35804\,
            I => \N__35771\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35803\,
            I => \N__35771\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35802\,
            I => \N__35768\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__35799\,
            I => \N__35765\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35760\
        );

    \I__7102\ : InMux
    port map (
            O => \N__35797\,
            I => \N__35760\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__35792\,
            I => \N__35751\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__35789\,
            I => \N__35751\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__35786\,
            I => \N__35748\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__35783\,
            I => \N__35743\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__35780\,
            I => \N__35743\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35735\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35735\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35735\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35732\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35729\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35768\,
            I => \N__35726\
        );

    \I__7090\ : Span4Mux_v
    port map (
            O => \N__35765\,
            I => \N__35723\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__35760\,
            I => \N__35720\
        );

    \I__7088\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35712\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35758\,
            I => \N__35712\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35712\
        );

    \I__7085\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35709\
        );

    \I__7084\ : Span4Mux_v
    port map (
            O => \N__35751\,
            I => \N__35706\
        );

    \I__7083\ : Span4Mux_v
    port map (
            O => \N__35748\,
            I => \N__35703\
        );

    \I__7082\ : Span4Mux_h
    port map (
            O => \N__35743\,
            I => \N__35698\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35742\,
            I => \N__35695\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__35735\,
            I => \N__35688\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__35732\,
            I => \N__35688\
        );

    \I__7078\ : Span4Mux_h
    port map (
            O => \N__35729\,
            I => \N__35688\
        );

    \I__7077\ : Span4Mux_v
    port map (
            O => \N__35726\,
            I => \N__35681\
        );

    \I__7076\ : Span4Mux_h
    port map (
            O => \N__35723\,
            I => \N__35681\
        );

    \I__7075\ : Span4Mux_v
    port map (
            O => \N__35720\,
            I => \N__35681\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35678\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__35712\,
            I => \N__35675\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__35709\,
            I => \N__35668\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__35706\,
            I => \N__35668\
        );

    \I__7070\ : Span4Mux_h
    port map (
            O => \N__35703\,
            I => \N__35668\
        );

    \I__7069\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35663\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35663\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__35698\,
            I => \N__35660\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35695\,
            I => \N__35653\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__35688\,
            I => \N__35653\
        );

    \I__7064\ : Span4Mux_v
    port map (
            O => \N__35681\,
            I => \N__35653\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__35678\,
            I => \N__35646\
        );

    \I__7062\ : Span4Mux_h
    port map (
            O => \N__35675\,
            I => \N__35646\
        );

    \I__7061\ : Span4Mux_h
    port map (
            O => \N__35668\,
            I => \N__35646\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__35663\,
            I => n20858
        );

    \I__7059\ : Odrv4
    port map (
            O => \N__35660\,
            I => n20858
        );

    \I__7058\ : Odrv4
    port map (
            O => \N__35653\,
            I => n20858
        );

    \I__7057\ : Odrv4
    port map (
            O => \N__35646\,
            I => n20858
        );

    \I__7056\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35613\
        );

    \I__7055\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35608\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35635\,
            I => \N__35608\
        );

    \I__7053\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35599\
        );

    \I__7052\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35599\
        );

    \I__7051\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35599\
        );

    \I__7050\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35599\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35595\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35586\
        );

    \I__7047\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35586\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35586\
        );

    \I__7045\ : InMux
    port map (
            O => \N__35626\,
            I => \N__35586\
        );

    \I__7044\ : InMux
    port map (
            O => \N__35625\,
            I => \N__35580\
        );

    \I__7043\ : InMux
    port map (
            O => \N__35624\,
            I => \N__35580\
        );

    \I__7042\ : InMux
    port map (
            O => \N__35623\,
            I => \N__35574\
        );

    \I__7041\ : InMux
    port map (
            O => \N__35622\,
            I => \N__35574\
        );

    \I__7040\ : CascadeMux
    port map (
            O => \N__35621\,
            I => \N__35571\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35620\,
            I => \N__35560\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35560\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35560\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35560\
        );

    \I__7035\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35548\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__35613\,
            I => \N__35545\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__35608\,
            I => \N__35542\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__35599\,
            I => \N__35539\
        );

    \I__7031\ : CascadeMux
    port map (
            O => \N__35598\,
            I => \N__35532\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35595\,
            I => \N__35521\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35586\,
            I => \N__35521\
        );

    \I__7028\ : CascadeMux
    port map (
            O => \N__35585\,
            I => \N__35517\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__35580\,
            I => \N__35514\
        );

    \I__7026\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35511\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35574\,
            I => \N__35508\
        );

    \I__7024\ : InMux
    port map (
            O => \N__35571\,
            I => \N__35503\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35503\
        );

    \I__7022\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35500\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__35560\,
            I => \N__35497\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35487\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35487\
        );

    \I__7018\ : InMux
    port map (
            O => \N__35557\,
            I => \N__35478\
        );

    \I__7017\ : InMux
    port map (
            O => \N__35556\,
            I => \N__35478\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35478\
        );

    \I__7015\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35478\
        );

    \I__7014\ : InMux
    port map (
            O => \N__35553\,
            I => \N__35473\
        );

    \I__7013\ : InMux
    port map (
            O => \N__35552\,
            I => \N__35473\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35470\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35465\
        );

    \I__7010\ : Span4Mux_h
    port map (
            O => \N__35545\,
            I => \N__35465\
        );

    \I__7009\ : Span4Mux_h
    port map (
            O => \N__35542\,
            I => \N__35460\
        );

    \I__7008\ : Span4Mux_h
    port map (
            O => \N__35539\,
            I => \N__35460\
        );

    \I__7007\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35449\
        );

    \I__7006\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35449\
        );

    \I__7005\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35449\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35535\,
            I => \N__35449\
        );

    \I__7003\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35446\
        );

    \I__7002\ : InMux
    port map (
            O => \N__35531\,
            I => \N__35443\
        );

    \I__7001\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35432\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35529\,
            I => \N__35432\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35528\,
            I => \N__35432\
        );

    \I__6998\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35432\
        );

    \I__6997\ : InMux
    port map (
            O => \N__35526\,
            I => \N__35432\
        );

    \I__6996\ : Span4Mux_v
    port map (
            O => \N__35521\,
            I => \N__35429\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35426\
        );

    \I__6994\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35423\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__35514\,
            I => \N__35420\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35511\,
            I => \N__35417\
        );

    \I__6991\ : Span4Mux_v
    port map (
            O => \N__35508\,
            I => \N__35412\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35503\,
            I => \N__35412\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35398\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__35497\,
            I => \N__35395\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35496\,
            I => \N__35383\
        );

    \I__6986\ : InMux
    port map (
            O => \N__35495\,
            I => \N__35383\
        );

    \I__6985\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35383\
        );

    \I__6984\ : InMux
    port map (
            O => \N__35493\,
            I => \N__35383\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35383\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__35487\,
            I => \N__35380\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__35478\,
            I => \N__35369\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__35473\,
            I => \N__35369\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__35470\,
            I => \N__35369\
        );

    \I__6978\ : Span4Mux_h
    port map (
            O => \N__35465\,
            I => \N__35369\
        );

    \I__6977\ : Span4Mux_v
    port map (
            O => \N__35460\,
            I => \N__35369\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35366\
        );

    \I__6975\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35363\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__35449\,
            I => \N__35360\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__35446\,
            I => \N__35353\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__35443\,
            I => \N__35353\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__35432\,
            I => \N__35353\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__35429\,
            I => \N__35350\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__35426\,
            I => \N__35339\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__35423\,
            I => \N__35339\
        );

    \I__6967\ : Span4Mux_v
    port map (
            O => \N__35420\,
            I => \N__35339\
        );

    \I__6966\ : Span4Mux_h
    port map (
            O => \N__35417\,
            I => \N__35339\
        );

    \I__6965\ : Span4Mux_h
    port map (
            O => \N__35412\,
            I => \N__35339\
        );

    \I__6964\ : InMux
    port map (
            O => \N__35411\,
            I => \N__35326\
        );

    \I__6963\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35326\
        );

    \I__6962\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35326\
        );

    \I__6961\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35326\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35326\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35326\
        );

    \I__6958\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35321\
        );

    \I__6957\ : InMux
    port map (
            O => \N__35404\,
            I => \N__35318\
        );

    \I__6956\ : InMux
    port map (
            O => \N__35403\,
            I => \N__35315\
        );

    \I__6955\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35312\
        );

    \I__6954\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35309\
        );

    \I__6953\ : Span4Mux_h
    port map (
            O => \N__35398\,
            I => \N__35304\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__35395\,
            I => \N__35304\
        );

    \I__6951\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35301\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__35383\,
            I => \N__35294\
        );

    \I__6949\ : Span4Mux_h
    port map (
            O => \N__35380\,
            I => \N__35294\
        );

    \I__6948\ : Span4Mux_v
    port map (
            O => \N__35369\,
            I => \N__35294\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35281\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__35363\,
            I => \N__35281\
        );

    \I__6945\ : Span4Mux_h
    port map (
            O => \N__35360\,
            I => \N__35281\
        );

    \I__6944\ : Span4Mux_h
    port map (
            O => \N__35353\,
            I => \N__35281\
        );

    \I__6943\ : Span4Mux_h
    port map (
            O => \N__35350\,
            I => \N__35281\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__35339\,
            I => \N__35281\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__35326\,
            I => \N__35278\
        );

    \I__6940\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35273\
        );

    \I__6939\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35273\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__35321\,
            I => adc_state_0
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__35318\,
            I => adc_state_0
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__35315\,
            I => adc_state_0
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__35312\,
            I => adc_state_0
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__35309\,
            I => adc_state_0
        );

    \I__6933\ : Odrv4
    port map (
            O => \N__35304\,
            I => adc_state_0
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__35301\,
            I => adc_state_0
        );

    \I__6931\ : Odrv4
    port map (
            O => \N__35294\,
            I => adc_state_0
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__35281\,
            I => adc_state_0
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__35278\,
            I => adc_state_0
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__35273\,
            I => adc_state_0
        );

    \I__6927\ : CascadeMux
    port map (
            O => \N__35250\,
            I => \N__35247\
        );

    \I__6926\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35244\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__35244\,
            I => \N__35241\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__35241\,
            I => \N__35237\
        );

    \I__6923\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35234\
        );

    \I__6922\ : Span4Mux_h
    port map (
            O => \N__35237\,
            I => \N__35228\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35228\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__35233\,
            I => \N__35225\
        );

    \I__6919\ : Span4Mux_h
    port map (
            O => \N__35228\,
            I => \N__35222\
        );

    \I__6918\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35219\
        );

    \I__6917\ : Odrv4
    port map (
            O => \N__35222\,
            I => cmd_rdadctmp_21
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__35219\,
            I => cmd_rdadctmp_21
        );

    \I__6915\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35208\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__35208\,
            I => \N__35205\
        );

    \I__6912\ : Span4Mux_h
    port map (
            O => \N__35205\,
            I => \N__35202\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__35202\,
            I => \N__35199\
        );

    \I__6910\ : Odrv4
    port map (
            O => \N__35199\,
            I => buf_data_iac_21
        );

    \I__6909\ : CascadeMux
    port map (
            O => \N__35196\,
            I => \N__35193\
        );

    \I__6908\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35190\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__35190\,
            I => \N__35187\
        );

    \I__6906\ : Span4Mux_v
    port map (
            O => \N__35187\,
            I => \N__35184\
        );

    \I__6905\ : Span4Mux_h
    port map (
            O => \N__35184\,
            I => \N__35181\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__35181\,
            I => n21124
        );

    \I__6903\ : InMux
    port map (
            O => \N__35178\,
            I => \N__35173\
        );

    \I__6902\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35169\
        );

    \I__6901\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35166\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__35173\,
            I => \N__35162\
        );

    \I__6899\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35159\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__35169\,
            I => \N__35156\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__35166\,
            I => \N__35153\
        );

    \I__6896\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35150\
        );

    \I__6895\ : Span4Mux_h
    port map (
            O => \N__35162\,
            I => \N__35147\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__35159\,
            I => \N__35143\
        );

    \I__6893\ : Span4Mux_h
    port map (
            O => \N__35156\,
            I => \N__35140\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__35153\,
            I => \N__35137\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__35150\,
            I => \N__35134\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__35147\,
            I => \N__35131\
        );

    \I__6889\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35128\
        );

    \I__6888\ : Span4Mux_h
    port map (
            O => \N__35143\,
            I => \N__35125\
        );

    \I__6887\ : Span4Mux_h
    port map (
            O => \N__35140\,
            I => \N__35120\
        );

    \I__6886\ : Span4Mux_v
    port map (
            O => \N__35137\,
            I => \N__35120\
        );

    \I__6885\ : Odrv12
    port map (
            O => \N__35134\,
            I => \comm_spi.n14603\
        );

    \I__6884\ : Odrv4
    port map (
            O => \N__35131\,
            I => \comm_spi.n14603\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__35128\,
            I => \comm_spi.n14603\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__35125\,
            I => \comm_spi.n14603\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__35120\,
            I => \comm_spi.n14603\
        );

    \I__6880\ : SRMux
    port map (
            O => \N__35109\,
            I => \N__35104\
        );

    \I__6879\ : SRMux
    port map (
            O => \N__35108\,
            I => \N__35101\
        );

    \I__6878\ : SRMux
    port map (
            O => \N__35107\,
            I => \N__35098\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__35104\,
            I => \N__35095\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__35101\,
            I => \N__35092\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__35098\,
            I => \N__35089\
        );

    \I__6874\ : Span4Mux_h
    port map (
            O => \N__35095\,
            I => \N__35086\
        );

    \I__6873\ : Span4Mux_v
    port map (
            O => \N__35092\,
            I => \N__35083\
        );

    \I__6872\ : Span4Mux_h
    port map (
            O => \N__35089\,
            I => \N__35080\
        );

    \I__6871\ : Span4Mux_v
    port map (
            O => \N__35086\,
            I => \N__35077\
        );

    \I__6870\ : Span4Mux_h
    port map (
            O => \N__35083\,
            I => \N__35072\
        );

    \I__6869\ : Span4Mux_v
    port map (
            O => \N__35080\,
            I => \N__35072\
        );

    \I__6868\ : Odrv4
    port map (
            O => \N__35077\,
            I => \comm_spi.data_tx_7__N_774\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__35072\,
            I => \comm_spi.data_tx_7__N_774\
        );

    \I__6866\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35062\
        );

    \I__6865\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35057\
        );

    \I__6864\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35057\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__35062\,
            I => \N__35052\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__35057\,
            I => \N__35052\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__35052\,
            I => comm_tx_buf_7
        );

    \I__6860\ : SRMux
    port map (
            O => \N__35049\,
            I => \N__35046\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__35046\,
            I => \N__35041\
        );

    \I__6858\ : SRMux
    port map (
            O => \N__35045\,
            I => \N__35038\
        );

    \I__6857\ : SRMux
    port map (
            O => \N__35044\,
            I => \N__35035\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__35041\,
            I => \N__35032\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__35038\,
            I => \N__35029\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N__35026\
        );

    \I__6853\ : Span4Mux_v
    port map (
            O => \N__35032\,
            I => \N__35023\
        );

    \I__6852\ : Span4Mux_h
    port map (
            O => \N__35029\,
            I => \N__35020\
        );

    \I__6851\ : Span4Mux_v
    port map (
            O => \N__35026\,
            I => \N__35017\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__35023\,
            I => \N__35014\
        );

    \I__6849\ : Span4Mux_h
    port map (
            O => \N__35020\,
            I => \N__35011\
        );

    \I__6848\ : Odrv4
    port map (
            O => \N__35017\,
            I => \comm_spi.data_tx_7__N_766\
        );

    \I__6847\ : Odrv4
    port map (
            O => \N__35014\,
            I => \comm_spi.data_tx_7__N_766\
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__35011\,
            I => \comm_spi.data_tx_7__N_766\
        );

    \I__6845\ : InMux
    port map (
            O => \N__35004\,
            I => \N__34998\
        );

    \I__6844\ : InMux
    port map (
            O => \N__35003\,
            I => \N__34998\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34998\,
            I => \N__34990\
        );

    \I__6842\ : InMux
    port map (
            O => \N__34997\,
            I => \N__34987\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34996\,
            I => \N__34980\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34980\
        );

    \I__6839\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34980\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34977\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__34990\,
            I => n12228
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34987\,
            I => n12228
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34980\,
            I => n12228
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34977\,
            I => n12228
        );

    \I__6833\ : InMux
    port map (
            O => \N__34968\,
            I => \N__34965\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__34965\,
            I => \N__34962\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__34962\,
            I => \N__34959\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__34959\,
            I => \N__34955\
        );

    \I__6829\ : CascadeMux
    port map (
            O => \N__34958\,
            I => \N__34952\
        );

    \I__6828\ : Span4Mux_h
    port map (
            O => \N__34955\,
            I => \N__34949\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34946\
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__34949\,
            I => buf_adcdata_vdc_9
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__34946\,
            I => buf_adcdata_vdc_9
        );

    \I__6824\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34938\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__34938\,
            I => \N__34934\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34930\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__34934\,
            I => \N__34927\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__34933\,
            I => \N__34924\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__34930\,
            I => \N__34921\
        );

    \I__6818\ : Sp12to4
    port map (
            O => \N__34927\,
            I => \N__34918\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34924\,
            I => \N__34915\
        );

    \I__6816\ : Span4Mux_v
    port map (
            O => \N__34921\,
            I => \N__34912\
        );

    \I__6815\ : Span12Mux_v
    port map (
            O => \N__34918\,
            I => \N__34909\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__34915\,
            I => buf_adcdata_vac_9
        );

    \I__6813\ : Odrv4
    port map (
            O => \N__34912\,
            I => buf_adcdata_vac_9
        );

    \I__6812\ : Odrv12
    port map (
            O => \N__34909\,
            I => buf_adcdata_vac_9
        );

    \I__6811\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34898\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34894\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__34898\,
            I => \N__34891\
        );

    \I__6808\ : InMux
    port map (
            O => \N__34897\,
            I => \N__34888\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34894\,
            I => \N__34881\
        );

    \I__6806\ : Span4Mux_h
    port map (
            O => \N__34891\,
            I => \N__34881\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__34888\,
            I => \N__34881\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__34881\,
            I => comm_tx_buf_3
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__34878\,
            I => \n21122_cascade_\
        );

    \I__6802\ : CascadeMux
    port map (
            O => \N__34875\,
            I => \N__34872\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34869\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__34869\,
            I => n21120
        );

    \I__6799\ : CEMux
    port map (
            O => \N__34866\,
            I => \N__34863\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34863\,
            I => \N__34860\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__34860\,
            I => n11361
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__34857\,
            I => \n7_adj_1616_cascade_\
        );

    \I__6795\ : CascadeMux
    port map (
            O => \N__34854\,
            I => \N__34851\
        );

    \I__6794\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34848\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__34848\,
            I => \ADC_VDC.n17509\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34842\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34842\,
            I => \ADC_VDC.n11265\
        );

    \I__6790\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34836\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__34836\,
            I => \ADC_VDC.n6\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__34833\,
            I => \ADC_VDC.n11265_cascade_\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34827\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__34827\,
            I => \N__34823\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34820\
        );

    \I__6784\ : Span4Mux_h
    port map (
            O => \N__34823\,
            I => \N__34817\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34814\
        );

    \I__6782\ : Odrv4
    port map (
            O => \N__34817\,
            I => \ADC_VDC.n15\
        );

    \I__6781\ : Odrv4
    port map (
            O => \N__34814\,
            I => \ADC_VDC.n15\
        );

    \I__6780\ : CascadeMux
    port map (
            O => \N__34809\,
            I => \ADC_VDC.n15_cascade_\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34803\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34800\
        );

    \I__6777\ : Odrv4
    port map (
            O => \N__34800\,
            I => \ADC_VDC.n20996\
        );

    \I__6776\ : CascadeMux
    port map (
            O => \N__34797\,
            I => \N__34777\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34773\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34768\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34753\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34793\,
            I => \N__34753\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34753\
        );

    \I__6770\ : InMux
    port map (
            O => \N__34791\,
            I => \N__34753\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34790\,
            I => \N__34753\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34753\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34753\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34787\,
            I => \N__34732\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34732\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34785\,
            I => \N__34732\
        );

    \I__6763\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34732\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34732\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34732\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34732\
        );

    \I__6759\ : InMux
    port map (
            O => \N__34780\,
            I => \N__34732\
        );

    \I__6758\ : InMux
    port map (
            O => \N__34777\,
            I => \N__34727\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34727\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__34773\,
            I => \N__34724\
        );

    \I__6755\ : SRMux
    port map (
            O => \N__34772\,
            I => \N__34721\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34718\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34715\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34753\,
            I => \N__34712\
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__34752\,
            I => \N__34707\
        );

    \I__6750\ : CEMux
    port map (
            O => \N__34751\,
            I => \N__34703\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34700\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34749\,
            I => \N__34697\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__34732\,
            I => \N__34692\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__34727\,
            I => \N__34692\
        );

    \I__6745\ : Span4Mux_v
    port map (
            O => \N__34724\,
            I => \N__34687\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34687\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__34718\,
            I => \N__34684\
        );

    \I__6742\ : Span4Mux_v
    port map (
            O => \N__34715\,
            I => \N__34679\
        );

    \I__6741\ : Span4Mux_v
    port map (
            O => \N__34712\,
            I => \N__34679\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34676\
        );

    \I__6739\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34673\
        );

    \I__6738\ : InMux
    port map (
            O => \N__34707\,
            I => \N__34670\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34667\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__34703\,
            I => \N__34664\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__34700\,
            I => \N__34661\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__34697\,
            I => \N__34656\
        );

    \I__6733\ : Span4Mux_v
    port map (
            O => \N__34692\,
            I => \N__34656\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__34687\,
            I => \N__34651\
        );

    \I__6731\ : Span4Mux_v
    port map (
            O => \N__34684\,
            I => \N__34651\
        );

    \I__6730\ : Span4Mux_h
    port map (
            O => \N__34679\,
            I => \N__34646\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__34676\,
            I => \N__34646\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34643\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__34670\,
            I => \N__34638\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__34667\,
            I => \N__34638\
        );

    \I__6725\ : Span4Mux_v
    port map (
            O => \N__34664\,
            I => \N__34629\
        );

    \I__6724\ : Span4Mux_h
    port map (
            O => \N__34661\,
            I => \N__34629\
        );

    \I__6723\ : Span4Mux_v
    port map (
            O => \N__34656\,
            I => \N__34629\
        );

    \I__6722\ : Span4Mux_h
    port map (
            O => \N__34651\,
            I => \N__34629\
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__34646\,
            I => dds_state_1_adj_1453
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__34643\,
            I => dds_state_1_adj_1453
        );

    \I__6719\ : Odrv12
    port map (
            O => \N__34638\,
            I => dds_state_1_adj_1453
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__34629\,
            I => dds_state_1_adj_1453
        );

    \I__6717\ : InMux
    port map (
            O => \N__34620\,
            I => \N__34606\
        );

    \I__6716\ : CascadeMux
    port map (
            O => \N__34619\,
            I => \N__34603\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34618\,
            I => \N__34577\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34617\,
            I => \N__34577\
        );

    \I__6713\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34577\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34615\,
            I => \N__34577\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34577\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34577\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34577\
        );

    \I__6708\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34577\
        );

    \I__6707\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34574\
        );

    \I__6706\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34571\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__34606\,
            I => \N__34568\
        );

    \I__6704\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34564\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34549\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34549\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34549\
        );

    \I__6700\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34549\
        );

    \I__6699\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34549\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34549\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34596\,
            I => \N__34549\
        );

    \I__6696\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34542\
        );

    \I__6695\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34542\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__34577\,
            I => \N__34537\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__34574\,
            I => \N__34537\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__34571\,
            I => \N__34533\
        );

    \I__6691\ : Span4Mux_h
    port map (
            O => \N__34568\,
            I => \N__34530\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34526\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34521\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__34549\,
            I => \N__34521\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34518\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34515\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34542\,
            I => \N__34512\
        );

    \I__6684\ : Span4Mux_v
    port map (
            O => \N__34537\,
            I => \N__34509\
        );

    \I__6683\ : InMux
    port map (
            O => \N__34536\,
            I => \N__34506\
        );

    \I__6682\ : Span4Mux_v
    port map (
            O => \N__34533\,
            I => \N__34501\
        );

    \I__6681\ : Span4Mux_h
    port map (
            O => \N__34530\,
            I => \N__34501\
        );

    \I__6680\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34498\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34526\,
            I => \N__34495\
        );

    \I__6678\ : Span12Mux_v
    port map (
            O => \N__34521\,
            I => \N__34492\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__34518\,
            I => \N__34489\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34484\
        );

    \I__6675\ : Span4Mux_v
    port map (
            O => \N__34512\,
            I => \N__34484\
        );

    \I__6674\ : Span4Mux_h
    port map (
            O => \N__34509\,
            I => \N__34477\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__34506\,
            I => \N__34477\
        );

    \I__6672\ : Span4Mux_h
    port map (
            O => \N__34501\,
            I => \N__34477\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__34498\,
            I => dds_state_2_adj_1452
        );

    \I__6670\ : Odrv4
    port map (
            O => \N__34495\,
            I => dds_state_2_adj_1452
        );

    \I__6669\ : Odrv12
    port map (
            O => \N__34492\,
            I => dds_state_2_adj_1452
        );

    \I__6668\ : Odrv4
    port map (
            O => \N__34489\,
            I => dds_state_2_adj_1452
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__34484\,
            I => dds_state_2_adj_1452
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__34477\,
            I => dds_state_2_adj_1452
        );

    \I__6665\ : InMux
    port map (
            O => \N__34464\,
            I => \N__34460\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34463\,
            I => \N__34454\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__34460\,
            I => \N__34450\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34459\,
            I => \N__34447\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34444\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34441\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__34454\,
            I => \N__34438\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34434\
        );

    \I__6657\ : Span4Mux_h
    port map (
            O => \N__34450\,
            I => \N__34431\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__34447\,
            I => \N__34426\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34444\,
            I => \N__34426\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__34441\,
            I => \N__34420\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__34438\,
            I => \N__34417\
        );

    \I__6652\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34414\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34407\
        );

    \I__6650\ : Span4Mux_h
    port map (
            O => \N__34431\,
            I => \N__34407\
        );

    \I__6649\ : Span4Mux_v
    port map (
            O => \N__34426\,
            I => \N__34407\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34404\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34399\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34399\
        );

    \I__6645\ : Odrv4
    port map (
            O => \N__34420\,
            I => dds_state_0_adj_1454
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__34417\,
            I => dds_state_0_adj_1454
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__34414\,
            I => dds_state_0_adj_1454
        );

    \I__6642\ : Odrv4
    port map (
            O => \N__34407\,
            I => dds_state_0_adj_1454
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__34404\,
            I => dds_state_0_adj_1454
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__34399\,
            I => dds_state_0_adj_1454
        );

    \I__6639\ : CEMux
    port map (
            O => \N__34386\,
            I => \N__34383\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__34383\,
            I => \N__34379\
        );

    \I__6637\ : CEMux
    port map (
            O => \N__34382\,
            I => \N__34376\
        );

    \I__6636\ : Span4Mux_v
    port map (
            O => \N__34379\,
            I => \N__34373\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__34376\,
            I => \N__34370\
        );

    \I__6634\ : Span4Mux_h
    port map (
            O => \N__34373\,
            I => \N__34367\
        );

    \I__6633\ : Span12Mux_v
    port map (
            O => \N__34370\,
            I => \N__34364\
        );

    \I__6632\ : Odrv4
    port map (
            O => \N__34367\,
            I => \CLK_DDS.n12784\
        );

    \I__6631\ : Odrv12
    port map (
            O => \N__34364\,
            I => \CLK_DDS.n12784\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34356\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__6628\ : Span4Mux_v
    port map (
            O => \N__34353\,
            I => \N__34349\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34346\
        );

    \I__6626\ : Span4Mux_v
    port map (
            O => \N__34349\,
            I => \N__34341\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__34346\,
            I => \N__34341\
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__34341\,
            I => \comm_spi.n14607\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34335\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__34335\,
            I => \ADC_VDC.n19_adj_1401\
        );

    \I__6621\ : CascadeMux
    port map (
            O => \N__34332\,
            I => \ADC_VDC.n21323_cascade_\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34326\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__34326\,
            I => \ADC_VDC.n21320\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34323\,
            I => \N__34320\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34320\,
            I => \N__34317\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__34317\,
            I => \ADC_VDC.n20965\
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__34314\,
            I => \ADC_VDC.n10_cascade_\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34308\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__34308\,
            I => \ADC_VDC.n20812\
        );

    \I__6612\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34302\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__34302\,
            I => \ADC_VDC.n20784\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__34299\,
            I => \n8_adj_1573_cascade_\
        );

    \I__6609\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34292\
        );

    \I__6608\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34289\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__34292\,
            I => \N__34286\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__34289\,
            I => \N__34281\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__34286\,
            I => \N__34278\
        );

    \I__6604\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34273\
        );

    \I__6603\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34273\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__34281\,
            I => eis_stop
        );

    \I__6601\ : Odrv4
    port map (
            O => \N__34278\,
            I => eis_stop
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__34273\,
            I => eis_stop
        );

    \I__6599\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34262\
        );

    \I__6598\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34258\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__34262\,
            I => \N__34255\
        );

    \I__6596\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34252\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__34258\,
            I => req_data_cnt_9
        );

    \I__6594\ : Odrv4
    port map (
            O => \N__34255\,
            I => req_data_cnt_9
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__34252\,
            I => req_data_cnt_9
        );

    \I__6592\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34242\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__34242\,
            I => n22375
        );

    \I__6590\ : CascadeMux
    port map (
            O => \N__34239\,
            I => \N__34236\
        );

    \I__6589\ : InMux
    port map (
            O => \N__34236\,
            I => \N__34233\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__34233\,
            I => \N__34230\
        );

    \I__6587\ : Span4Mux_v
    port map (
            O => \N__34230\,
            I => \N__34227\
        );

    \I__6586\ : Span4Mux_v
    port map (
            O => \N__34227\,
            I => \N__34224\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__34224\,
            I => n22381
        );

    \I__6584\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34218\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__34218\,
            I => \N__34215\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__34215\,
            I => \N__34212\
        );

    \I__6581\ : Span4Mux_v
    port map (
            O => \N__34212\,
            I => \N__34209\
        );

    \I__6580\ : Odrv4
    port map (
            O => \N__34209\,
            I => n22384
        );

    \I__6579\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34203\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__34203\,
            I => \N__34200\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__34200\,
            I => n11396
        );

    \I__6576\ : IoInMux
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34194\,
            I => \N__34191\
        );

    \I__6574\ : IoSpan4Mux
    port map (
            O => \N__34191\,
            I => \N__34188\
        );

    \I__6573\ : IoSpan4Mux
    port map (
            O => \N__34188\,
            I => \N__34185\
        );

    \I__6572\ : Span4Mux_s3_v
    port map (
            O => \N__34185\,
            I => \N__34182\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__34182\,
            I => \N__34179\
        );

    \I__6570\ : Span4Mux_v
    port map (
            O => \N__34179\,
            I => \N__34175\
        );

    \I__6569\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34172\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__34175\,
            I => \DDS_SCK\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__34172\,
            I => \DDS_SCK\
        );

    \I__6566\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34164\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__34164\,
            I => \N__34161\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__34161\,
            I => \N__34158\
        );

    \I__6563\ : Odrv4
    port map (
            O => \N__34158\,
            I => \comm_spi.n14605\
        );

    \I__6562\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34152\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__34152\,
            I => \N__34149\
        );

    \I__6560\ : Span4Mux_h
    port map (
            O => \N__34149\,
            I => \N__34146\
        );

    \I__6559\ : Odrv4
    port map (
            O => \N__34146\,
            I => \comm_spi.n14604\
        );

    \I__6558\ : IoInMux
    port map (
            O => \N__34143\,
            I => \N__34140\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__34140\,
            I => \N__34137\
        );

    \I__6556\ : IoSpan4Mux
    port map (
            O => \N__34137\,
            I => \N__34134\
        );

    \I__6555\ : Span4Mux_s3_h
    port map (
            O => \N__34134\,
            I => \N__34131\
        );

    \I__6554\ : Sp12to4
    port map (
            O => \N__34131\,
            I => \N__34128\
        );

    \I__6553\ : Span12Mux_h
    port map (
            O => \N__34128\,
            I => \N__34125\
        );

    \I__6552\ : Odrv12
    port map (
            O => \N__34125\,
            I => \ICE_SPI_MISO\
        );

    \I__6551\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34119\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__34119\,
            I => n20_adj_1617
        );

    \I__6549\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34113\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__34113\,
            I => \N__34108\
        );

    \I__6547\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34105\
        );

    \I__6546\ : InMux
    port map (
            O => \N__34111\,
            I => \N__34102\
        );

    \I__6545\ : Span4Mux_h
    port map (
            O => \N__34108\,
            I => \N__34099\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__34105\,
            I => \N__34094\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__34102\,
            I => \N__34094\
        );

    \I__6542\ : Odrv4
    port map (
            O => \N__34099\,
            I => n10717
        );

    \I__6541\ : Odrv12
    port map (
            O => \N__34094\,
            I => n10717
        );

    \I__6540\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34084\
        );

    \I__6539\ : InMux
    port map (
            O => \N__34088\,
            I => \N__34079\
        );

    \I__6538\ : InMux
    port map (
            O => \N__34087\,
            I => \N__34079\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__34084\,
            I => req_data_cnt_12
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__34079\,
            I => req_data_cnt_12
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__34074\,
            I => \N__34069\
        );

    \I__6534\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34066\
        );

    \I__6533\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34063\
        );

    \I__6532\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34060\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__34066\,
            I => \acadc_skipCount_9\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__34063\,
            I => \acadc_skipCount_9\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__34060\,
            I => \acadc_skipCount_9\
        );

    \I__6528\ : InMux
    port map (
            O => \N__34053\,
            I => \N__34050\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__34050\,
            I => \N__34047\
        );

    \I__6526\ : Odrv12
    port map (
            O => \N__34047\,
            I => n19_adj_1607
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__34044\,
            I => \n29_cascade_\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__34041\,
            I => \N__34038\
        );

    \I__6523\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34034\
        );

    \I__6522\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34031\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__34034\,
            I => \N__34025\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34025\
        );

    \I__6519\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34022\
        );

    \I__6518\ : Span4Mux_v
    port map (
            O => \N__34025\,
            I => \N__34019\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__34022\,
            I => n16_adj_1603
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__34019\,
            I => n16_adj_1603
        );

    \I__6515\ : InMux
    port map (
            O => \N__34014\,
            I => \N__34011\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__34011\,
            I => n24
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__34008\,
            I => \n21_adj_1492_cascade_\
        );

    \I__6512\ : InMux
    port map (
            O => \N__34005\,
            I => \N__34002\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__34002\,
            I => n30_adj_1618
        );

    \I__6510\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33996\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__33996\,
            I => \N__33993\
        );

    \I__6508\ : Span4Mux_v
    port map (
            O => \N__33993\,
            I => \N__33989\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33992\,
            I => \N__33985\
        );

    \I__6506\ : Span4Mux_h
    port map (
            O => \N__33989\,
            I => \N__33982\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33979\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33985\,
            I => buf_dds1_4
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__33982\,
            I => buf_dds1_4
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__33979\,
            I => buf_dds1_4
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__33972\,
            I => \N__33969\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33964\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33961\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33967\,
            I => \N__33958\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33964\,
            I => \N__33953\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33953\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33958\,
            I => buf_dds0_0
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__33953\,
            I => buf_dds0_0
        );

    \I__6493\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33945\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__33945\,
            I => \N__33941\
        );

    \I__6491\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33937\
        );

    \I__6490\ : Span4Mux_h
    port map (
            O => \N__33941\,
            I => \N__33934\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33931\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__33937\,
            I => req_data_cnt_13
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__33934\,
            I => req_data_cnt_13
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33931\,
            I => req_data_cnt_13
        );

    \I__6485\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33920\
        );

    \I__6484\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33916\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__33920\,
            I => \N__33913\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33919\,
            I => \N__33910\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__33916\,
            I => buf_dds1_0
        );

    \I__6480\ : Odrv12
    port map (
            O => \N__33913\,
            I => buf_dds1_0
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33910\,
            I => buf_dds1_0
        );

    \I__6478\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33900\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33900\,
            I => n22_adj_1615
        );

    \I__6476\ : CascadeMux
    port map (
            O => \N__33897\,
            I => \n10717_cascade_\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33894\,
            I => \N__33891\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33891\,
            I => \N__33888\
        );

    \I__6473\ : Odrv4
    port map (
            O => \N__33888\,
            I => n21344
        );

    \I__6472\ : InMux
    port map (
            O => \N__33885\,
            I => \N__33880\
        );

    \I__6471\ : InMux
    port map (
            O => \N__33884\,
            I => \N__33877\
        );

    \I__6470\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33874\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__33880\,
            I => \N__33871\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33877\,
            I => \N__33868\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__33874\,
            I => \N__33863\
        );

    \I__6466\ : Span4Mux_v
    port map (
            O => \N__33871\,
            I => \N__33863\
        );

    \I__6465\ : Span4Mux_h
    port map (
            O => \N__33868\,
            I => \N__33860\
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__33863\,
            I => buf_dds1_5
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__33860\,
            I => buf_dds1_5
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__33855\,
            I => \N__33852\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33852\,
            I => \N__33849\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__33849\,
            I => \N__33844\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33841\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33847\,
            I => \N__33838\
        );

    \I__6457\ : Span4Mux_v
    port map (
            O => \N__33844\,
            I => \N__33833\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__33841\,
            I => \N__33833\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__33838\,
            I => buf_dds1_7
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__33833\,
            I => buf_dds1_7
        );

    \I__6453\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33825\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__33825\,
            I => \N__33822\
        );

    \I__6451\ : Span4Mux_v
    port map (
            O => \N__33822\,
            I => \N__33817\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33812\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33812\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__33817\,
            I => \acadc_skipCount_14\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__33812\,
            I => \acadc_skipCount_14\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33807\,
            I => \N__33803\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33799\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__33803\,
            I => \N__33796\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33793\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__33799\,
            I => \N__33790\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__33796\,
            I => \N__33787\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__33793\,
            I => buf_dds0_4
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__33790\,
            I => buf_dds0_4
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__33787\,
            I => buf_dds0_4
        );

    \I__6437\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33777\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33777\,
            I => \N__33773\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33770\
        );

    \I__6434\ : Span4Mux_v
    port map (
            O => \N__33773\,
            I => \N__33767\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__33770\,
            I => comm_buf_6_3
        );

    \I__6432\ : Odrv4
    port map (
            O => \N__33767\,
            I => comm_buf_6_3
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__33762\,
            I => \N__33759\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33759\,
            I => \N__33755\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33751\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__33755\,
            I => \N__33748\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33754\,
            I => \N__33745\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__33751\,
            I => buf_dds1_1
        );

    \I__6425\ : Odrv4
    port map (
            O => \N__33748\,
            I => buf_dds1_1
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33745\,
            I => buf_dds1_1
        );

    \I__6423\ : InMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33730\
        );

    \I__6421\ : InMux
    port map (
            O => \N__33734\,
            I => \N__33727\
        );

    \I__6420\ : InMux
    port map (
            O => \N__33733\,
            I => \N__33724\
        );

    \I__6419\ : Odrv12
    port map (
            O => \N__33730\,
            I => cmd_rdadctmp_9_adj_1441
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__33727\,
            I => cmd_rdadctmp_9_adj_1441
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__33724\,
            I => cmd_rdadctmp_9_adj_1441
        );

    \I__6416\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33714\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__33714\,
            I => \N__33710\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33706\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__33710\,
            I => \N__33703\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__33709\,
            I => \N__33700\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__33706\,
            I => \N__33697\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__33703\,
            I => \N__33694\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33691\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__33697\,
            I => \N__33686\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__33694\,
            I => \N__33686\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33691\,
            I => buf_adcdata_vac_1
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__33686\,
            I => buf_adcdata_vac_1
        );

    \I__6404\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33667\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33664\
        );

    \I__6402\ : CascadeMux
    port map (
            O => \N__33679\,
            I => \N__33659\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33652\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33652\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33644\
        );

    \I__6398\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33641\
        );

    \I__6397\ : CascadeMux
    port map (
            O => \N__33674\,
            I => \N__33638\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33631\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33631\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33631\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33628\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33667\,
            I => \N__33625\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__33664\,
            I => \N__33622\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33615\
        );

    \I__6389\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33615\
        );

    \I__6388\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33610\
        );

    \I__6387\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33610\
        );

    \I__6386\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33607\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__33652\,
            I => \N__33604\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33598\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33650\,
            I => \N__33598\
        );

    \I__6382\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33591\
        );

    \I__6381\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33591\
        );

    \I__6380\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33591\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__33644\,
            I => \N__33588\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__33641\,
            I => \N__33585\
        );

    \I__6377\ : InMux
    port map (
            O => \N__33638\,
            I => \N__33582\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33579\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33576\
        );

    \I__6374\ : Span4Mux_h
    port map (
            O => \N__33625\,
            I => \N__33571\
        );

    \I__6373\ : Span4Mux_h
    port map (
            O => \N__33622\,
            I => \N__33571\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33566\
        );

    \I__6371\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33566\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__33615\,
            I => \N__33563\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__33610\,
            I => \N__33556\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33556\
        );

    \I__6367\ : Span4Mux_h
    port map (
            O => \N__33604\,
            I => \N__33556\
        );

    \I__6366\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33553\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__33598\,
            I => \N__33544\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__33591\,
            I => \N__33544\
        );

    \I__6363\ : Span4Mux_h
    port map (
            O => \N__33588\,
            I => \N__33544\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__33585\,
            I => \N__33544\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__33582\,
            I => \N__33535\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__33579\,
            I => \N__33535\
        );

    \I__6359\ : Span4Mux_h
    port map (
            O => \N__33576\,
            I => \N__33535\
        );

    \I__6358\ : Span4Mux_v
    port map (
            O => \N__33571\,
            I => \N__33535\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__33566\,
            I => \N__33530\
        );

    \I__6356\ : Span4Mux_h
    port map (
            O => \N__33563\,
            I => \N__33530\
        );

    \I__6355\ : Span4Mux_h
    port map (
            O => \N__33556\,
            I => \N__33527\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__33553\,
            I => \N__33522\
        );

    \I__6353\ : Span4Mux_v
    port map (
            O => \N__33544\,
            I => \N__33522\
        );

    \I__6352\ : Span4Mux_v
    port map (
            O => \N__33535\,
            I => \N__33519\
        );

    \I__6351\ : Span4Mux_v
    port map (
            O => \N__33530\,
            I => \N__33514\
        );

    \I__6350\ : Span4Mux_h
    port map (
            O => \N__33527\,
            I => \N__33514\
        );

    \I__6349\ : Odrv4
    port map (
            O => \N__33522\,
            I => n20853
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__33519\,
            I => n20853
        );

    \I__6347\ : Odrv4
    port map (
            O => \N__33514\,
            I => n20853
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__33507\,
            I => \N__33498\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__33506\,
            I => \N__33495\
        );

    \I__6344\ : InMux
    port map (
            O => \N__33505\,
            I => \N__33466\
        );

    \I__6343\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33466\
        );

    \I__6342\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33466\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33466\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33463\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33460\
        );

    \I__6338\ : InMux
    port map (
            O => \N__33495\,
            I => \N__33451\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33494\,
            I => \N__33451\
        );

    \I__6336\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33439\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33439\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33439\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33439\
        );

    \I__6332\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33439\
        );

    \I__6331\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33432\
        );

    \I__6330\ : InMux
    port map (
            O => \N__33487\,
            I => \N__33432\
        );

    \I__6329\ : InMux
    port map (
            O => \N__33486\,
            I => \N__33432\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33485\,
            I => \N__33421\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33421\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33421\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33421\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33481\,
            I => \N__33421\
        );

    \I__6323\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33410\
        );

    \I__6322\ : InMux
    port map (
            O => \N__33479\,
            I => \N__33410\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33410\
        );

    \I__6320\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33410\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33410\
        );

    \I__6318\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33407\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33404\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33463\,
            I => \N__33399\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__33460\,
            I => \N__33399\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33394\
        );

    \I__6313\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33394\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__33457\,
            I => \N__33391\
        );

    \I__6311\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33384\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__33451\,
            I => \N__33381\
        );

    \I__6309\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33370\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__33439\,
            I => \N__33367\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__33432\,
            I => \N__33360\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__33421\,
            I => \N__33360\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__33410\,
            I => \N__33360\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__33407\,
            I => \N__33357\
        );

    \I__6303\ : Span4Mux_h
    port map (
            O => \N__33404\,
            I => \N__33354\
        );

    \I__6302\ : Span4Mux_v
    port map (
            O => \N__33399\,
            I => \N__33351\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__33394\,
            I => \N__33348\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33340\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33335\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33389\,
            I => \N__33335\
        );

    \I__6297\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33332\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33329\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__33384\,
            I => \N__33324\
        );

    \I__6294\ : Span4Mux_v
    port map (
            O => \N__33381\,
            I => \N__33324\
        );

    \I__6293\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33313\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33313\
        );

    \I__6291\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33313\
        );

    \I__6290\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33313\
        );

    \I__6289\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33313\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__33375\,
            I => \N__33310\
        );

    \I__6287\ : InMux
    port map (
            O => \N__33374\,
            I => \N__33301\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33373\,
            I => \N__33301\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__33370\,
            I => \N__33292\
        );

    \I__6284\ : Span4Mux_h
    port map (
            O => \N__33367\,
            I => \N__33292\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__33360\,
            I => \N__33292\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__33357\,
            I => \N__33292\
        );

    \I__6281\ : Span4Mux_v
    port map (
            O => \N__33354\,
            I => \N__33285\
        );

    \I__6280\ : Span4Mux_v
    port map (
            O => \N__33351\,
            I => \N__33285\
        );

    \I__6279\ : Span4Mux_h
    port map (
            O => \N__33348\,
            I => \N__33285\
        );

    \I__6278\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33278\
        );

    \I__6277\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33278\
        );

    \I__6276\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33278\
        );

    \I__6275\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33275\
        );

    \I__6274\ : CascadeMux
    port map (
            O => \N__33343\,
            I => \N__33269\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__33340\,
            I => \N__33261\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__33335\,
            I => \N__33254\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33254\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__33329\,
            I => \N__33251\
        );

    \I__6269\ : Span4Mux_h
    port map (
            O => \N__33324\,
            I => \N__33246\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33246\
        );

    \I__6267\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33234\
        );

    \I__6266\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33234\
        );

    \I__6265\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33234\
        );

    \I__6264\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33234\
        );

    \I__6263\ : InMux
    port map (
            O => \N__33306\,
            I => \N__33234\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33301\,
            I => \N__33227\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__33292\,
            I => \N__33227\
        );

    \I__6260\ : Span4Mux_h
    port map (
            O => \N__33285\,
            I => \N__33227\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33222\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__33275\,
            I => \N__33222\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33213\
        );

    \I__6256\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33213\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33210\
        );

    \I__6254\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33207\
        );

    \I__6253\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33202\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33202\
        );

    \I__6251\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33195\
        );

    \I__6250\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33195\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33195\
        );

    \I__6248\ : Span4Mux_h
    port map (
            O => \N__33261\,
            I => \N__33192\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33189\
        );

    \I__6246\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33186\
        );

    \I__6245\ : Span12Mux_v
    port map (
            O => \N__33254\,
            I => \N__33183\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__33251\,
            I => \N__33178\
        );

    \I__6243\ : Span4Mux_v
    port map (
            O => \N__33246\,
            I => \N__33178\
        );

    \I__6242\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33175\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__33234\,
            I => \N__33168\
        );

    \I__6240\ : Sp12to4
    port map (
            O => \N__33227\,
            I => \N__33168\
        );

    \I__6239\ : Span12Mux_h
    port map (
            O => \N__33222\,
            I => \N__33168\
        );

    \I__6238\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33161\
        );

    \I__6237\ : InMux
    port map (
            O => \N__33220\,
            I => \N__33161\
        );

    \I__6236\ : InMux
    port map (
            O => \N__33219\,
            I => \N__33161\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33218\,
            I => \N__33158\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__33213\,
            I => adc_state_0_adj_1418
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__33210\,
            I => adc_state_0_adj_1418
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__33207\,
            I => adc_state_0_adj_1418
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__33202\,
            I => adc_state_0_adj_1418
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__33195\,
            I => adc_state_0_adj_1418
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__33192\,
            I => adc_state_0_adj_1418
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__33189\,
            I => adc_state_0_adj_1418
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__33186\,
            I => adc_state_0_adj_1418
        );

    \I__6226\ : Odrv12
    port map (
            O => \N__33183\,
            I => adc_state_0_adj_1418
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__33178\,
            I => adc_state_0_adj_1418
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__33175\,
            I => adc_state_0_adj_1418
        );

    \I__6223\ : Odrv12
    port map (
            O => \N__33168\,
            I => adc_state_0_adj_1418
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__33161\,
            I => adc_state_0_adj_1418
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__33158\,
            I => adc_state_0_adj_1418
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__33129\,
            I => \N__33124\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33121\
        );

    \I__6218\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33116\
        );

    \I__6217\ : InMux
    port map (
            O => \N__33124\,
            I => \N__33116\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__33121\,
            I => cmd_rdadctmp_18_adj_1432
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__33116\,
            I => cmd_rdadctmp_18_adj_1432
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__33111\,
            I => \N__33108\
        );

    \I__6213\ : InMux
    port map (
            O => \N__33108\,
            I => \N__33105\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__33105\,
            I => \N__33102\
        );

    \I__6211\ : Span12Mux_h
    port map (
            O => \N__33102\,
            I => \N__33099\
        );

    \I__6210\ : Odrv12
    port map (
            O => \N__33099\,
            I => n9_adj_1416
        );

    \I__6209\ : CascadeMux
    port map (
            O => \N__33096\,
            I => \n31_adj_1613_cascade_\
        );

    \I__6208\ : CEMux
    port map (
            O => \N__33093\,
            I => \N__33089\
        );

    \I__6207\ : CEMux
    port map (
            O => \N__33092\,
            I => \N__33086\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__33089\,
            I => \N__33083\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__33086\,
            I => \N__33080\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__33083\,
            I => n12085
        );

    \I__6203\ : Odrv12
    port map (
            O => \N__33080\,
            I => n12085
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__33075\,
            I => \n12085_cascade_\
        );

    \I__6201\ : SRMux
    port map (
            O => \N__33072\,
            I => \N__33068\
        );

    \I__6200\ : SRMux
    port map (
            O => \N__33071\,
            I => \N__33065\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__33068\,
            I => \N__33062\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__33065\,
            I => \N__33059\
        );

    \I__6197\ : Span4Mux_h
    port map (
            O => \N__33062\,
            I => \N__33056\
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__33059\,
            I => n14764
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__33056\,
            I => n14764
        );

    \I__6194\ : CascadeMux
    port map (
            O => \N__33051\,
            I => \n12228_cascade_\
        );

    \I__6193\ : InMux
    port map (
            O => \N__33048\,
            I => \N__33044\
        );

    \I__6192\ : InMux
    port map (
            O => \N__33047\,
            I => \N__33041\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__33044\,
            I => comm_buf_6_7
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__33041\,
            I => comm_buf_6_7
        );

    \I__6189\ : InMux
    port map (
            O => \N__33036\,
            I => \N__33033\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__33033\,
            I => n20850
        );

    \I__6187\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33027\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__33027\,
            I => n20852
        );

    \I__6185\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__33021\,
            I => comm_buf_2_3
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__33018\,
            I => \n22387_cascade_\
        );

    \I__6182\ : InMux
    port map (
            O => \N__33015\,
            I => \N__33012\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__33012\,
            I => n21193
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__33009\,
            I => \n22390_cascade_\
        );

    \I__6179\ : CascadeMux
    port map (
            O => \N__33006\,
            I => \n4_adj_1587_cascade_\
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__33003\,
            I => \n21175_cascade_\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__33000\,
            I => \n2358_cascade_\
        );

    \I__6176\ : CascadeMux
    port map (
            O => \N__32997\,
            I => \n20850_cascade_\
        );

    \I__6175\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32991\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32988\
        );

    \I__6173\ : Span4Mux_v
    port map (
            O => \N__32988\,
            I => \N__32985\
        );

    \I__6172\ : Odrv4
    port map (
            O => \N__32985\,
            I => n30_adj_1482
        );

    \I__6171\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32979\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__32979\,
            I => \N__32976\
        );

    \I__6169\ : Span4Mux_h
    port map (
            O => \N__32976\,
            I => \N__32973\
        );

    \I__6168\ : Span4Mux_h
    port map (
            O => \N__32973\,
            I => \N__32970\
        );

    \I__6167\ : Odrv4
    port map (
            O => \N__32970\,
            I => n30_adj_1625
        );

    \I__6166\ : InMux
    port map (
            O => \N__32967\,
            I => \N__32964\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__32964\,
            I => comm_buf_2_7
        );

    \I__6164\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32958\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32958\,
            I => \N__32955\
        );

    \I__6162\ : Span4Mux_h
    port map (
            O => \N__32955\,
            I => \N__32952\
        );

    \I__6161\ : Span4Mux_h
    port map (
            O => \N__32952\,
            I => \N__32949\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__32949\,
            I => n30_adj_1628
        );

    \I__6159\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32943\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32943\,
            I => \N__32940\
        );

    \I__6157\ : Span4Mux_h
    port map (
            O => \N__32940\,
            I => \N__32937\
        );

    \I__6156\ : Odrv4
    port map (
            O => \N__32937\,
            I => n30_adj_1631
        );

    \I__6155\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32931\,
            I => \N__32928\
        );

    \I__6153\ : Odrv12
    port map (
            O => \N__32928\,
            I => n30_adj_1634
        );

    \I__6152\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__6150\ : Odrv4
    port map (
            O => \N__32919\,
            I => n30_adj_1638
        );

    \I__6149\ : InMux
    port map (
            O => \N__32916\,
            I => \N__32913\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__32913\,
            I => \N__32910\
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__32910\,
            I => n30_adj_1641
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__32907\,
            I => \n4_adj_1594_cascade_\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32901\,
            I => \ADC_VDC.n21229\
        );

    \I__6143\ : CEMux
    port map (
            O => \N__32898\,
            I => \N__32895\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32892\
        );

    \I__6141\ : Odrv12
    port map (
            O => \N__32892\,
            I => \ADC_VDC.n47\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32886\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32883\
        );

    \I__6138\ : Span4Mux_v
    port map (
            O => \N__32883\,
            I => \N__32879\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32876\
        );

    \I__6136\ : Odrv4
    port map (
            O => \N__32879\,
            I => \comm_spi.n14608\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__32876\,
            I => \comm_spi.n14608\
        );

    \I__6134\ : CascadeMux
    port map (
            O => \N__32871\,
            I => \N__32868\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32865\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32861\
        );

    \I__6131\ : CascadeMux
    port map (
            O => \N__32864\,
            I => \N__32858\
        );

    \I__6130\ : Span4Mux_v
    port map (
            O => \N__32861\,
            I => \N__32855\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32852\
        );

    \I__6128\ : Odrv4
    port map (
            O => \N__32855\,
            I => buf_adcdata_vdc_1
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__32852\,
            I => buf_adcdata_vdc_1
        );

    \I__6126\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32843\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32839\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32836\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32833\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32839\,
            I => \N__32828\
        );

    \I__6121\ : Span12Mux_s9_h
    port map (
            O => \N__32836\,
            I => \N__32828\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__32833\,
            I => buf_adcdata_iac_1
        );

    \I__6119\ : Odrv12
    port map (
            O => \N__32828\,
            I => buf_adcdata_iac_1
        );

    \I__6118\ : CascadeMux
    port map (
            O => \N__32823\,
            I => \n19_adj_1491_cascade_\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32817\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__32817\,
            I => \N__32814\
        );

    \I__6115\ : Span4Mux_h
    port map (
            O => \N__32814\,
            I => \N__32811\
        );

    \I__6114\ : Span4Mux_h
    port map (
            O => \N__32811\,
            I => \N__32808\
        );

    \I__6113\ : Odrv4
    port map (
            O => \N__32808\,
            I => buf_data_iac_1
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__32805\,
            I => \n22_adj_1488_cascade_\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32799\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32799\,
            I => n30_adj_1506
        );

    \I__6109\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32793\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32793\,
            I => comm_buf_2_1
        );

    \I__6107\ : CascadeMux
    port map (
            O => \N__32790\,
            I => \n22249_cascade_\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__32787\,
            I => \ADC_VDC.n77_cascade_\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__32781\,
            I => \ADC_VDC.n12\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32778\,
            I => \N__32775\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__32775\,
            I => \ADC_VDC.n20899\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__32772\,
            I => \ADC_VDC.n72_cascade_\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__32769\,
            I => \ADC_VDC.n31_cascade_\
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__32766\,
            I => \ADC_VDC.n22195_cascade_\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__32763\,
            I => \ADC_VDC.n22198_cascade_\
        );

    \I__6097\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32757\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__32757\,
            I => \N__32754\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__32754\,
            I => \N__32751\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__32751\,
            I => \N__32748\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__32748\,
            I => \ADC_VDC.n18566\
        );

    \I__6092\ : CEMux
    port map (
            O => \N__32745\,
            I => \N__32742\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__32742\,
            I => \N__32739\
        );

    \I__6090\ : Odrv4
    port map (
            O => \N__32739\,
            I => \ADC_VDC.n20811\
        );

    \I__6089\ : CascadeMux
    port map (
            O => \N__32736\,
            I => \ADC_VDC.n6_adj_1399_cascade_\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32730\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__32730\,
            I => \N__32727\
        );

    \I__6086\ : Span4Mux_h
    port map (
            O => \N__32727\,
            I => \N__32723\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32726\,
            I => \N__32720\
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__32723\,
            I => \ADC_VDC.n10536\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__32720\,
            I => \ADC_VDC.n10536\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32712\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__32712\,
            I => \N__32708\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32705\
        );

    \I__6079\ : Span4Mux_v
    port map (
            O => \N__32708\,
            I => \N__32702\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__32705\,
            I => acadc_skipcnt_13
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__32702\,
            I => acadc_skipcnt_13
        );

    \I__6076\ : InMux
    port map (
            O => \N__32697\,
            I => n19622
        );

    \I__6075\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32690\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32687\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__32690\,
            I => \N__32684\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32687\,
            I => acadc_skipcnt_14
        );

    \I__6071\ : Odrv4
    port map (
            O => \N__32684\,
            I => acadc_skipcnt_14
        );

    \I__6070\ : InMux
    port map (
            O => \N__32679\,
            I => n19623
        );

    \I__6069\ : InMux
    port map (
            O => \N__32676\,
            I => n19624
        );

    \I__6068\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32669\
        );

    \I__6067\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32666\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__32669\,
            I => \N__32663\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__32666\,
            I => acadc_skipcnt_15
        );

    \I__6064\ : Odrv12
    port map (
            O => \N__32663\,
            I => acadc_skipcnt_15
        );

    \I__6063\ : CEMux
    port map (
            O => \N__32658\,
            I => \N__32653\
        );

    \I__6062\ : CEMux
    port map (
            O => \N__32657\,
            I => \N__32650\
        );

    \I__6061\ : CEMux
    port map (
            O => \N__32656\,
            I => \N__32647\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32643\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32650\,
            I => \N__32638\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32638\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32635\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__32643\,
            I => \N__32630\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__32638\,
            I => \N__32630\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32627\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__32630\,
            I => n11654
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__32627\,
            I => n11654
        );

    \I__6051\ : SRMux
    port map (
            O => \N__32622\,
            I => \N__32619\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__32619\,
            I => \N__32615\
        );

    \I__6049\ : SRMux
    port map (
            O => \N__32618\,
            I => \N__32612\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__32615\,
            I => \N__32609\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__32612\,
            I => \N__32606\
        );

    \I__6046\ : Span4Mux_h
    port map (
            O => \N__32609\,
            I => \N__32601\
        );

    \I__6045\ : Span4Mux_v
    port map (
            O => \N__32606\,
            I => \N__32601\
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__32601\,
            I => n14671
        );

    \I__6043\ : CEMux
    port map (
            O => \N__32598\,
            I => \N__32595\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__32595\,
            I => \N__32592\
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__32592\,
            I => \ADC_VDC.n17\
        );

    \I__6040\ : SRMux
    port map (
            O => \N__32589\,
            I => \N__32586\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__32586\,
            I => \N__32583\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__32583\,
            I => \N__32580\
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__32580\,
            I => \ADC_VDC.n4\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32577\,
            I => \N__32574\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__32574\,
            I => \ADC_VDC.n7_adj_1398\
        );

    \I__6034\ : CascadeMux
    port map (
            O => \N__32571\,
            I => \ADC_VDC.n7_adj_1398_cascade_\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32564\
        );

    \I__6032\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32561\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__32564\,
            I => \ADC_VDC.n77\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__32561\,
            I => \ADC_VDC.n77\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__32556\,
            I => \N__32552\
        );

    \I__6028\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32549\
        );

    \I__6027\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32546\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__32549\,
            I => acadc_skipcnt_4
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__32546\,
            I => acadc_skipcnt_4
        );

    \I__6024\ : InMux
    port map (
            O => \N__32541\,
            I => n19613
        );

    \I__6023\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32534\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32531\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32528\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__32531\,
            I => acadc_skipcnt_5
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__32528\,
            I => acadc_skipcnt_5
        );

    \I__6018\ : InMux
    port map (
            O => \N__32523\,
            I => n19614
        );

    \I__6017\ : InMux
    port map (
            O => \N__32520\,
            I => n19615
        );

    \I__6016\ : InMux
    port map (
            O => \N__32517\,
            I => n19616
        );

    \I__6015\ : InMux
    port map (
            O => \N__32514\,
            I => \N__32510\
        );

    \I__6014\ : InMux
    port map (
            O => \N__32513\,
            I => \N__32507\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__32510\,
            I => \N__32504\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__32507\,
            I => acadc_skipcnt_8
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__32504\,
            I => acadc_skipcnt_8
        );

    \I__6010\ : InMux
    port map (
            O => \N__32499\,
            I => n19617
        );

    \I__6009\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32492\
        );

    \I__6008\ : InMux
    port map (
            O => \N__32495\,
            I => \N__32489\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__32492\,
            I => \N__32486\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__32489\,
            I => acadc_skipcnt_9
        );

    \I__6005\ : Odrv4
    port map (
            O => \N__32486\,
            I => acadc_skipcnt_9
        );

    \I__6004\ : InMux
    port map (
            O => \N__32481\,
            I => \bfn_12_20_0_\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32478\,
            I => \N__32475\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__32475\,
            I => \N__32471\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32468\
        );

    \I__6000\ : Span4Mux_h
    port map (
            O => \N__32471\,
            I => \N__32465\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__32468\,
            I => acadc_skipcnt_10
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__32465\,
            I => acadc_skipcnt_10
        );

    \I__5997\ : InMux
    port map (
            O => \N__32460\,
            I => n19619
        );

    \I__5996\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32453\
        );

    \I__5995\ : InMux
    port map (
            O => \N__32456\,
            I => \N__32450\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32453\,
            I => \N__32447\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__32450\,
            I => acadc_skipcnt_11
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__32447\,
            I => acadc_skipcnt_11
        );

    \I__5991\ : InMux
    port map (
            O => \N__32442\,
            I => n19620
        );

    \I__5990\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32436\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__32436\,
            I => \N__32432\
        );

    \I__5988\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32429\
        );

    \I__5987\ : Span4Mux_h
    port map (
            O => \N__32432\,
            I => \N__32426\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__32429\,
            I => acadc_skipcnt_12
        );

    \I__5985\ : Odrv4
    port map (
            O => \N__32426\,
            I => acadc_skipcnt_12
        );

    \I__5984\ : InMux
    port map (
            O => \N__32421\,
            I => n19621
        );

    \I__5983\ : InMux
    port map (
            O => \N__32418\,
            I => \N__32414\
        );

    \I__5982\ : InMux
    port map (
            O => \N__32417\,
            I => \N__32411\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__32414\,
            I => acadc_skipcnt_1
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__32411\,
            I => acadc_skipcnt_1
        );

    \I__5979\ : InMux
    port map (
            O => \N__32406\,
            I => \bfn_12_19_0_\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32403\,
            I => n19611
        );

    \I__5977\ : InMux
    port map (
            O => \N__32400\,
            I => \N__32396\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32393\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__32396\,
            I => \N__32390\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__32393\,
            I => acadc_skipcnt_3
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__32390\,
            I => acadc_skipcnt_3
        );

    \I__5972\ : InMux
    port map (
            O => \N__32385\,
            I => n19612
        );

    \I__5971\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32379\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__32379\,
            I => n23_adj_1501
        );

    \I__5969\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__32373\,
            I => n24_adj_1642
        );

    \I__5967\ : InMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__5965\ : Span4Mux_h
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__5964\ : Span4Mux_v
    port map (
            O => \N__32361\,
            I => \N__32356\
        );

    \I__5963\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32351\
        );

    \I__5962\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32351\
        );

    \I__5961\ : Odrv4
    port map (
            O => \N__32356\,
            I => \acadc_skipCount_15\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__32351\,
            I => \acadc_skipCount_15\
        );

    \I__5959\ : SRMux
    port map (
            O => \N__32346\,
            I => \N__32343\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32340\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__32340\,
            I => \N__32337\
        );

    \I__5956\ : Span4Mux_v
    port map (
            O => \N__32337\,
            I => \N__32334\
        );

    \I__5955\ : Odrv4
    port map (
            O => \N__32334\,
            I => n21037
        );

    \I__5954\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32328\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__32328\,
            I => \SIG_DDS.tmp_buf_6\
        );

    \I__5952\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32322\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__32322\,
            I => \N__32318\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32321\,
            I => \N__32314\
        );

    \I__5949\ : Span4Mux_v
    port map (
            O => \N__32318\,
            I => \N__32311\
        );

    \I__5948\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32308\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__32314\,
            I => buf_dds0_7
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__32311\,
            I => buf_dds0_7
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__32308\,
            I => buf_dds0_7
        );

    \I__5944\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32298\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32298\,
            I => \SIG_DDS.tmp_buf_7\
        );

    \I__5942\ : InMux
    port map (
            O => \N__32295\,
            I => \N__32291\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32287\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__32291\,
            I => \N__32284\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32281\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32287\,
            I => \acadc_skipCount_12\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__32284\,
            I => \acadc_skipCount_12\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__32281\,
            I => \acadc_skipCount_12\
        );

    \I__5935\ : CascadeMux
    port map (
            O => \N__32274\,
            I => \N__32269\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__32273\,
            I => \N__32266\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32272\,
            I => \N__32263\
        );

    \I__5932\ : InMux
    port map (
            O => \N__32269\,
            I => \N__32260\
        );

    \I__5931\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32257\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__32263\,
            I => \N__32252\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__32260\,
            I => \N__32252\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__32257\,
            I => \acadc_skipCount_10\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__32252\,
            I => \acadc_skipCount_10\
        );

    \I__5926\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32244\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N__32240\
        );

    \I__5924\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32236\
        );

    \I__5923\ : Span4Mux_h
    port map (
            O => \N__32240\,
            I => \N__32233\
        );

    \I__5922\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32230\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32236\,
            I => \acadc_skipCount_13\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__32233\,
            I => \acadc_skipCount_13\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__32230\,
            I => \acadc_skipCount_13\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32220\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__32220\,
            I => n20
        );

    \I__5916\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32214\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__32214\,
            I => \N__32208\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32201\
        );

    \I__5913\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32201\
        );

    \I__5912\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32198\
        );

    \I__5911\ : Span4Mux_h
    port map (
            O => \N__32208\,
            I => \N__32195\
        );

    \I__5910\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32190\
        );

    \I__5909\ : InMux
    port map (
            O => \N__32206\,
            I => \N__32190\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32187\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__32198\,
            I => acadc_dtrig_v
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__32195\,
            I => acadc_dtrig_v
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__32190\,
            I => acadc_dtrig_v
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__32187\,
            I => acadc_dtrig_v
        );

    \I__5903\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32170\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32165\
        );

    \I__5901\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32165\
        );

    \I__5900\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32158\
        );

    \I__5899\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32158\
        );

    \I__5898\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32158\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__32170\,
            I => acadc_dtrig_i
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__32165\,
            I => acadc_dtrig_i
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__32158\,
            I => acadc_dtrig_i
        );

    \I__5894\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__32148\,
            I => n4_adj_1546
        );

    \I__5892\ : InMux
    port map (
            O => \N__32145\,
            I => \N__32141\
        );

    \I__5891\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32138\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__32141\,
            I => \N__32135\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__32138\,
            I => \N__32131\
        );

    \I__5888\ : Span4Mux_h
    port map (
            O => \N__32135\,
            I => \N__32128\
        );

    \I__5887\ : InMux
    port map (
            O => \N__32134\,
            I => \N__32125\
        );

    \I__5886\ : Span4Mux_h
    port map (
            O => \N__32131\,
            I => \N__32122\
        );

    \I__5885\ : Span4Mux_v
    port map (
            O => \N__32128\,
            I => \N__32119\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__32125\,
            I => buf_dds0_1
        );

    \I__5883\ : Odrv4
    port map (
            O => \N__32122\,
            I => buf_dds0_1
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__32119\,
            I => buf_dds0_1
        );

    \I__5881\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32109\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__32109\,
            I => \SIG_DDS.tmp_buf_0\
        );

    \I__5879\ : InMux
    port map (
            O => \N__32106\,
            I => \N__32103\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__32103\,
            I => \SIG_DDS.tmp_buf_1\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32100\,
            I => \N__32097\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__32097\,
            I => \SIG_DDS.tmp_buf_2\
        );

    \I__5875\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32091\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__32091\,
            I => \SIG_DDS.tmp_buf_14\
        );

    \I__5873\ : CascadeMux
    port map (
            O => \N__32088\,
            I => \N__32085\
        );

    \I__5872\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32082\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__32082\,
            I => \N__32079\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__32079\,
            I => \N__32075\
        );

    \I__5869\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32071\
        );

    \I__5868\ : Span4Mux_v
    port map (
            O => \N__32075\,
            I => \N__32068\
        );

    \I__5867\ : InMux
    port map (
            O => \N__32074\,
            I => \N__32065\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__32071\,
            I => buf_dds0_15
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__32068\,
            I => buf_dds0_15
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__32065\,
            I => buf_dds0_15
        );

    \I__5863\ : InMux
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__32055\,
            I => \SIG_DDS.tmp_buf_3\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__32052\,
            I => \N__32049\
        );

    \I__5860\ : InMux
    port map (
            O => \N__32049\,
            I => \N__32046\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__32046\,
            I => \SIG_DDS.tmp_buf_4\
        );

    \I__5858\ : CascadeMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__5857\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__32032\
        );

    \I__5855\ : InMux
    port map (
            O => \N__32036\,
            I => \N__32029\
        );

    \I__5854\ : InMux
    port map (
            O => \N__32035\,
            I => \N__32026\
        );

    \I__5853\ : Span12Mux_h
    port map (
            O => \N__32032\,
            I => \N__32023\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__32029\,
            I => \N__32020\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__32026\,
            I => buf_dds0_8
        );

    \I__5850\ : Odrv12
    port map (
            O => \N__32023\,
            I => buf_dds0_8
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__32020\,
            I => buf_dds0_8
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__32013\,
            I => \N__32010\
        );

    \I__5847\ : InMux
    port map (
            O => \N__32010\,
            I => \N__32007\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__32004\,
            I => \SIG_DDS.tmp_buf_8\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__32001\,
            I => \N__31998\
        );

    \I__5843\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31995\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__31995\,
            I => \N__31990\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31987\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__31993\,
            I => \N__31984\
        );

    \I__5839\ : Span12Mux_v
    port map (
            O => \N__31990\,
            I => \N__31981\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31987\,
            I => \N__31978\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31975\
        );

    \I__5836\ : Odrv12
    port map (
            O => \N__31981\,
            I => cmd_rdadctmp_19
        );

    \I__5835\ : Odrv4
    port map (
            O => \N__31978\,
            I => cmd_rdadctmp_19
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__31975\,
            I => cmd_rdadctmp_19
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__31968\,
            I => \N__31965\
        );

    \I__5832\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31960\
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__31964\,
            I => \N__31957\
        );

    \I__5830\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31954\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31960\,
            I => \N__31951\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31948\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31943\
        );

    \I__5826\ : Span4Mux_h
    port map (
            O => \N__31951\,
            I => \N__31943\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31948\,
            I => cmd_rdadctmp_25
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__31943\,
            I => cmd_rdadctmp_25
        );

    \I__5823\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31934\
        );

    \I__5822\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31930\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__31934\,
            I => \N__31927\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__31933\,
            I => \N__31924\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__31930\,
            I => \N__31921\
        );

    \I__5818\ : Span12Mux_h
    port map (
            O => \N__31927\,
            I => \N__31918\
        );

    \I__5817\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31915\
        );

    \I__5816\ : Span4Mux_h
    port map (
            O => \N__31921\,
            I => \N__31912\
        );

    \I__5815\ : Span12Mux_v
    port map (
            O => \N__31918\,
            I => \N__31909\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31915\,
            I => buf_adcdata_iac_22
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__31912\,
            I => buf_adcdata_iac_22
        );

    \I__5812\ : Odrv12
    port map (
            O => \N__31909\,
            I => buf_adcdata_iac_22
        );

    \I__5811\ : IoInMux
    port map (
            O => \N__31902\,
            I => \N__31899\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__5809\ : Span4Mux_s2_h
    port map (
            O => \N__31896\,
            I => \N__31892\
        );

    \I__5808\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31889\
        );

    \I__5807\ : Sp12to4
    port map (
            O => \N__31892\,
            I => \N__31886\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__31889\,
            I => \N__31882\
        );

    \I__5805\ : Span12Mux_v
    port map (
            O => \N__31886\,
            I => \N__31879\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31876\
        );

    \I__5803\ : Span4Mux_h
    port map (
            O => \N__31882\,
            I => \N__31873\
        );

    \I__5802\ : Odrv12
    port map (
            O => \N__31879\,
            I => \VAC_FLT0\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31876\,
            I => \VAC_FLT0\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__31873\,
            I => \VAC_FLT0\
        );

    \I__5799\ : IoInMux
    port map (
            O => \N__31866\,
            I => \N__31863\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31860\
        );

    \I__5797\ : Span4Mux_s0_h
    port map (
            O => \N__31860\,
            I => \N__31856\
        );

    \I__5796\ : CascadeMux
    port map (
            O => \N__31859\,
            I => \N__31853\
        );

    \I__5795\ : Sp12to4
    port map (
            O => \N__31856\,
            I => \N__31850\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31853\,
            I => \N__31846\
        );

    \I__5793\ : Span12Mux_v
    port map (
            O => \N__31850\,
            I => \N__31843\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__31849\,
            I => \N__31840\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__31846\,
            I => \N__31837\
        );

    \I__5790\ : Span12Mux_h
    port map (
            O => \N__31843\,
            I => \N__31834\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31831\
        );

    \I__5788\ : Span4Mux_v
    port map (
            O => \N__31837\,
            I => \N__31828\
        );

    \I__5787\ : Odrv12
    port map (
            O => \N__31834\,
            I => \VDC_RNG0\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31831\,
            I => \VDC_RNG0\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__31828\,
            I => \VDC_RNG0\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__31821\,
            I => \N__31818\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31815\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31815\,
            I => \N__31812\
        );

    \I__5781\ : Span4Mux_v
    port map (
            O => \N__31812\,
            I => \N__31809\
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__31809\,
            I => \SIG_DDS.n10\
        );

    \I__5779\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31803\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__31803\,
            I => \N__31799\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31795\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__31799\,
            I => \N__31792\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31798\,
            I => \N__31789\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31795\,
            I => buf_dds1_10
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__31792\,
            I => buf_dds1_10
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__31789\,
            I => buf_dds1_10
        );

    \I__5771\ : IoInMux
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31776\
        );

    \I__5769\ : Span4Mux_s1_v
    port map (
            O => \N__31776\,
            I => \N__31772\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31769\
        );

    \I__5767\ : Sp12to4
    port map (
            O => \N__31772\,
            I => \N__31766\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__31769\,
            I => \N__31762\
        );

    \I__5765\ : Span12Mux_h
    port map (
            O => \N__31766\,
            I => \N__31759\
        );

    \I__5764\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31756\
        );

    \I__5763\ : Span4Mux_v
    port map (
            O => \N__31762\,
            I => \N__31753\
        );

    \I__5762\ : Odrv12
    port map (
            O => \N__31759\,
            I => \SELIRNG0\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__31756\,
            I => \SELIRNG0\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__31753\,
            I => \SELIRNG0\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31743\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__31740\,
            I => \N__31737\
        );

    \I__5756\ : Span4Mux_h
    port map (
            O => \N__31737\,
            I => \N__31734\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__31731\,
            I => buf_data_iac_3
        );

    \I__5753\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__31725\,
            I => n22_adj_1637
        );

    \I__5751\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31718\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31721\,
            I => \N__31715\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__31718\,
            I => \N__31712\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31706\
        );

    \I__5747\ : Span4Mux_v
    port map (
            O => \N__31712\,
            I => \N__31706\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__31711\,
            I => \N__31703\
        );

    \I__5745\ : Span4Mux_h
    port map (
            O => \N__31706\,
            I => \N__31700\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31703\,
            I => \N__31697\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__31700\,
            I => cmd_rdadctmp_17_adj_1433
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__31697\,
            I => cmd_rdadctmp_17_adj_1433
        );

    \I__5741\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31678\
        );

    \I__5740\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31678\
        );

    \I__5739\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31673\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31673\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31661\
        );

    \I__5736\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31661\
        );

    \I__5735\ : InMux
    port map (
            O => \N__31686\,
            I => \N__31661\
        );

    \I__5734\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31648\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31648\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31648\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__31678\,
            I => \N__31645\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31642\
        );

    \I__5729\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31637\
        );

    \I__5728\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31637\
        );

    \I__5727\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31630\
        );

    \I__5726\ : InMux
    port map (
            O => \N__31669\,
            I => \N__31630\
        );

    \I__5725\ : InMux
    port map (
            O => \N__31668\,
            I => \N__31630\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__31661\,
            I => \N__31625\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31620\
        );

    \I__5722\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31620\
        );

    \I__5721\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31610\
        );

    \I__5720\ : InMux
    port map (
            O => \N__31657\,
            I => \N__31610\
        );

    \I__5719\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31610\
        );

    \I__5718\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31610\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__31648\,
            I => \N__31607\
        );

    \I__5716\ : Span4Mux_v
    port map (
            O => \N__31645\,
            I => \N__31598\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__31642\,
            I => \N__31598\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__31637\,
            I => \N__31598\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__31630\,
            I => \N__31598\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31629\,
            I => \N__31593\
        );

    \I__5711\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31593\
        );

    \I__5710\ : Span4Mux_v
    port map (
            O => \N__31625\,
            I => \N__31587\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__31620\,
            I => \N__31587\
        );

    \I__5708\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31584\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__31610\,
            I => \N__31581\
        );

    \I__5706\ : Span4Mux_v
    port map (
            O => \N__31607\,
            I => \N__31574\
        );

    \I__5705\ : Span4Mux_h
    port map (
            O => \N__31598\,
            I => \N__31574\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__31593\,
            I => \N__31574\
        );

    \I__5703\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31571\
        );

    \I__5702\ : Span4Mux_h
    port map (
            O => \N__31587\,
            I => \N__31566\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__31584\,
            I => \N__31566\
        );

    \I__5700\ : Span12Mux_v
    port map (
            O => \N__31581\,
            I => \N__31556\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__31574\,
            I => \N__31553\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31550\
        );

    \I__5697\ : Span4Mux_h
    port map (
            O => \N__31566\,
            I => \N__31547\
        );

    \I__5696\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31542\
        );

    \I__5695\ : InMux
    port map (
            O => \N__31564\,
            I => \N__31542\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31537\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31562\,
            I => \N__31537\
        );

    \I__5692\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31530\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31530\
        );

    \I__5690\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31530\
        );

    \I__5689\ : Odrv12
    port map (
            O => \N__31556\,
            I => n12653
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__31553\,
            I => n12653
        );

    \I__5687\ : Odrv12
    port map (
            O => \N__31550\,
            I => n12653
        );

    \I__5686\ : Odrv4
    port map (
            O => \N__31547\,
            I => n12653
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__31542\,
            I => n12653
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__31537\,
            I => n12653
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__31530\,
            I => n12653
        );

    \I__5682\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31511\
        );

    \I__5681\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31508\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31505\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__31508\,
            I => \N__31502\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__31505\,
            I => \N__31499\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__31502\,
            I => \N__31495\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__31499\,
            I => \N__31492\
        );

    \I__5675\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31489\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__31495\,
            I => cmd_rdadctmp_19_adj_1431
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__31492\,
            I => cmd_rdadctmp_19_adj_1431
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__31489\,
            I => cmd_rdadctmp_19_adj_1431
        );

    \I__5671\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31478\
        );

    \I__5670\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31475\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__31478\,
            I => secclk_cnt_21
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__31475\,
            I => secclk_cnt_21
        );

    \I__5667\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31466\
        );

    \I__5666\ : InMux
    port map (
            O => \N__31469\,
            I => \N__31463\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__31466\,
            I => secclk_cnt_19
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__31463\,
            I => secclk_cnt_19
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__31458\,
            I => \N__31454\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31451\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31448\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__31451\,
            I => secclk_cnt_12
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__31448\,
            I => secclk_cnt_12
        );

    \I__5658\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31439\
        );

    \I__5657\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31436\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__31439\,
            I => secclk_cnt_22
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__31436\,
            I => secclk_cnt_22
        );

    \I__5654\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31428\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__31428\,
            I => \N__31425\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__31425\,
            I => n14_adj_1599
        );

    \I__5651\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31419\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__31419\,
            I => \N__31415\
        );

    \I__5649\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31412\
        );

    \I__5648\ : Sp12to4
    port map (
            O => \N__31415\,
            I => \N__31407\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__31412\,
            I => \N__31407\
        );

    \I__5646\ : Odrv12
    port map (
            O => \N__31407\,
            I => \comm_spi.n14610\
        );

    \I__5645\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31400\
        );

    \I__5644\ : CascadeMux
    port map (
            O => \N__31403\,
            I => \N__31397\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__31400\,
            I => \N__31394\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31391\
        );

    \I__5641\ : Odrv12
    port map (
            O => \N__31394\,
            I => \buf_readRTD_14\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__31391\,
            I => \buf_readRTD_14\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31386\,
            I => \N__31382\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__31385\,
            I => \N__31379\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__31382\,
            I => \N__31375\
        );

    \I__5636\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31372\
        );

    \I__5635\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31368\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__31375\,
            I => \N__31365\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__31372\,
            I => \N__31362\
        );

    \I__5632\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31359\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__31368\,
            I => \N__31356\
        );

    \I__5630\ : Span4Mux_v
    port map (
            O => \N__31365\,
            I => \N__31353\
        );

    \I__5629\ : Span4Mux_v
    port map (
            O => \N__31362\,
            I => \N__31349\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__31359\,
            I => \N__31346\
        );

    \I__5627\ : Span12Mux_s11_h
    port map (
            O => \N__31356\,
            I => \N__31343\
        );

    \I__5626\ : Span4Mux_v
    port map (
            O => \N__31353\,
            I => \N__31340\
        );

    \I__5625\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31337\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__31349\,
            I => \N__31332\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__31346\,
            I => \N__31332\
        );

    \I__5622\ : Odrv12
    port map (
            O => \N__31343\,
            I => \buf_cfgRTD_6\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__31340\,
            I => \buf_cfgRTD_6\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__31337\,
            I => \buf_cfgRTD_6\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__31332\,
            I => \buf_cfgRTD_6\
        );

    \I__5618\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31316\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__31319\,
            I => \N__31313\
        );

    \I__5615\ : Span4Mux_h
    port map (
            O => \N__31316\,
            I => \N__31310\
        );

    \I__5614\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31307\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__31310\,
            I => \buf_readRTD_15\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__31307\,
            I => \buf_readRTD_15\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__31302\,
            I => \N__31297\
        );

    \I__5610\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31294\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__31300\,
            I => \N__31291\
        );

    \I__5608\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31288\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__31294\,
            I => \N__31284\
        );

    \I__5606\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31281\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31277\
        );

    \I__5604\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31274\
        );

    \I__5603\ : Sp12to4
    port map (
            O => \N__31284\,
            I => \N__31269\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31269\
        );

    \I__5601\ : CascadeMux
    port map (
            O => \N__31280\,
            I => \N__31266\
        );

    \I__5600\ : Span4Mux_v
    port map (
            O => \N__31277\,
            I => \N__31263\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31274\,
            I => \N__31260\
        );

    \I__5598\ : Span12Mux_v
    port map (
            O => \N__31269\,
            I => \N__31257\
        );

    \I__5597\ : InMux
    port map (
            O => \N__31266\,
            I => \N__31254\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__31263\,
            I => \N__31249\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__31260\,
            I => \N__31249\
        );

    \I__5594\ : Odrv12
    port map (
            O => \N__31257\,
            I => \buf_cfgRTD_7\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__31254\,
            I => \buf_cfgRTD_7\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__31249\,
            I => \buf_cfgRTD_7\
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__31242\,
            I => \N__31239\
        );

    \I__5590\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31236\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__5588\ : Span4Mux_h
    port map (
            O => \N__31233\,
            I => \N__31230\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__31230\,
            I => n20_adj_1528
        );

    \I__5586\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31223\
        );

    \I__5585\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31220\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31223\,
            I => secclk_cnt_16
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__31220\,
            I => secclk_cnt_16
        );

    \I__5582\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31211\
        );

    \I__5581\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31208\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__31211\,
            I => secclk_cnt_2
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__31208\,
            I => secclk_cnt_2
        );

    \I__5578\ : CascadeMux
    port map (
            O => \N__31203\,
            I => \N__31200\
        );

    \I__5577\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31196\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31193\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__31196\,
            I => secclk_cnt_7
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31193\,
            I => secclk_cnt_7
        );

    \I__5573\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31184\
        );

    \I__5572\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31181\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__31184\,
            I => secclk_cnt_13
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__31181\,
            I => secclk_cnt_13
        );

    \I__5569\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31173\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__31173\,
            I => n27_adj_1597
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__31170\,
            I => \n26_adj_1575_cascade_\
        );

    \I__5566\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__31164\,
            I => n25_adj_1574
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__31161\,
            I => \n19856_cascade_\
        );

    \I__5563\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31154\
        );

    \I__5562\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31151\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__31154\,
            I => secclk_cnt_20
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__31151\,
            I => secclk_cnt_20
        );

    \I__5559\ : SRMux
    port map (
            O => \N__31146\,
            I => \N__31142\
        );

    \I__5558\ : SRMux
    port map (
            O => \N__31145\,
            I => \N__31139\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__31142\,
            I => \N__31134\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__31139\,
            I => \N__31131\
        );

    \I__5555\ : SRMux
    port map (
            O => \N__31138\,
            I => \N__31128\
        );

    \I__5554\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31125\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__31134\,
            I => \N__31122\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__31131\,
            I => \N__31117\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31117\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__31125\,
            I => \N__31114\
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__31122\,
            I => n14715
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__31117\,
            I => n14715
        );

    \I__5547\ : Odrv12
    port map (
            O => \N__31114\,
            I => n14715
        );

    \I__5546\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31103\
        );

    \I__5545\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31100\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__31103\,
            I => secclk_cnt_0
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__31100\,
            I => secclk_cnt_0
        );

    \I__5542\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31091\
        );

    \I__5541\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31088\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__31091\,
            I => secclk_cnt_18
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__31088\,
            I => secclk_cnt_18
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__31083\,
            I => \N__31079\
        );

    \I__5537\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31076\
        );

    \I__5536\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31073\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__31076\,
            I => secclk_cnt_11
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__31073\,
            I => secclk_cnt_11
        );

    \I__5533\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31064\
        );

    \I__5532\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31061\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__31064\,
            I => secclk_cnt_4
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__31061\,
            I => secclk_cnt_4
        );

    \I__5529\ : InMux
    port map (
            O => \N__31056\,
            I => \N__31053\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__31053\,
            I => n28_adj_1505
        );

    \I__5527\ : InMux
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__5525\ : Span4Mux_h
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__5524\ : Span4Mux_h
    port map (
            O => \N__31041\,
            I => \N__31036\
        );

    \I__5523\ : InMux
    port map (
            O => \N__31040\,
            I => \N__31033\
        );

    \I__5522\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31030\
        );

    \I__5521\ : Span4Mux_h
    port map (
            O => \N__31036\,
            I => \N__31027\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__31033\,
            I => \N__31024\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__31030\,
            I => buf_adcdata_iac_3
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__31027\,
            I => buf_adcdata_iac_3
        );

    \I__5517\ : Odrv4
    port map (
            O => \N__31024\,
            I => buf_adcdata_iac_3
        );

    \I__5516\ : InMux
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__31014\,
            I => \N__31011\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__31011\,
            I => n19_adj_1636
        );

    \I__5513\ : InMux
    port map (
            O => \N__31008\,
            I => \N__31004\
        );

    \I__5512\ : InMux
    port map (
            O => \N__31007\,
            I => \N__31001\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__31004\,
            I => secclk_cnt_17
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__31001\,
            I => secclk_cnt_17
        );

    \I__5509\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30992\
        );

    \I__5508\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30989\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__30992\,
            I => secclk_cnt_9
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__30989\,
            I => secclk_cnt_9
        );

    \I__5505\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30981\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__30981\,
            I => n10_adj_1601
        );

    \I__5503\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__30975\,
            I => \N__30971\
        );

    \I__5501\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30968\
        );

    \I__5500\ : Odrv12
    port map (
            O => \N__30971\,
            I => dds0_mclkcnt_6
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__30968\,
            I => dds0_mclkcnt_6
        );

    \I__5498\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30960\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__30960\,
            I => \N__30957\
        );

    \I__5496\ : Odrv12
    port map (
            O => \N__30957\,
            I => n20799
        );

    \I__5495\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30950\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30947\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30950\,
            I => secclk_cnt_6
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__30947\,
            I => secclk_cnt_6
        );

    \I__5491\ : InMux
    port map (
            O => \N__30942\,
            I => \N__30938\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30935\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30938\,
            I => secclk_cnt_14
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__30935\,
            I => secclk_cnt_14
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__30930\,
            I => \N__30926\
        );

    \I__5486\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30923\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30920\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__30923\,
            I => secclk_cnt_10
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30920\,
            I => secclk_cnt_10
        );

    \I__5482\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30911\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30908\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30911\,
            I => secclk_cnt_3
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__30908\,
            I => secclk_cnt_3
        );

    \I__5478\ : InMux
    port map (
            O => \N__30903\,
            I => \N__30899\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30896\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__30899\,
            I => secclk_cnt_15
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30896\,
            I => secclk_cnt_15
        );

    \I__5474\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30887\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30884\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30887\,
            I => secclk_cnt_8
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__30884\,
            I => secclk_cnt_8
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__30879\,
            I => \N__30875\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30872\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30869\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30872\,
            I => secclk_cnt_1
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30869\,
            I => secclk_cnt_1
        );

    \I__5465\ : InMux
    port map (
            O => \N__30864\,
            I => \N__30860\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30857\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30860\,
            I => secclk_cnt_5
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__30857\,
            I => secclk_cnt_5
        );

    \I__5461\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30848\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30851\,
            I => \N__30845\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__30848\,
            I => dds0_mclkcnt_5
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__30845\,
            I => dds0_mclkcnt_5
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__30840\,
            I => \N__30836\
        );

    \I__5456\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30833\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30830\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__30833\,
            I => dds0_mclkcnt_1
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__30830\,
            I => dds0_mclkcnt_1
        );

    \I__5452\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30821\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30824\,
            I => \N__30818\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30821\,
            I => dds0_mclkcnt_4
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__30818\,
            I => dds0_mclkcnt_4
        );

    \I__5448\ : InMux
    port map (
            O => \N__30813\,
            I => \N__30809\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30812\,
            I => \N__30806\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__30809\,
            I => dds0_mclkcnt_2
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__30806\,
            I => dds0_mclkcnt_2
        );

    \I__5444\ : InMux
    port map (
            O => \N__30801\,
            I => \N__30797\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30794\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__30797\,
            I => dds0_mclkcnt_0
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__30794\,
            I => dds0_mclkcnt_0
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__30789\,
            I => \n12_adj_1480_cascade_\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30782\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30779\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__30782\,
            I => dds0_mclkcnt_7
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__30779\,
            I => dds0_mclkcnt_7
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__30774\,
            I => \n20799_cascade_\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30768\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30768\,
            I => n10
        );

    \I__5432\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30762\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30762\,
            I => \N__30758\
        );

    \I__5430\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30755\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__30758\,
            I => \comm_spi.n14611\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30755\,
            I => \comm_spi.n14611\
        );

    \I__5427\ : InMux
    port map (
            O => \N__30750\,
            I => \N__30746\
        );

    \I__5426\ : CEMux
    port map (
            O => \N__30749\,
            I => \N__30743\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30740\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30743\,
            I => \N__30737\
        );

    \I__5423\ : Span12Mux_h
    port map (
            O => \N__30740\,
            I => \N__30734\
        );

    \I__5422\ : Odrv4
    port map (
            O => \N__30737\,
            I => \ADC_VAC.n12594\
        );

    \I__5421\ : Odrv12
    port map (
            O => \N__30734\,
            I => \ADC_VAC.n12594\
        );

    \I__5420\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30725\
        );

    \I__5419\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30722\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__30725\,
            I => \N__30717\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30722\,
            I => \N__30714\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30710\
        );

    \I__5415\ : CascadeMux
    port map (
            O => \N__30720\,
            I => \N__30703\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__30717\,
            I => \N__30697\
        );

    \I__5413\ : Sp12to4
    port map (
            O => \N__30714\,
            I => \N__30694\
        );

    \I__5412\ : InMux
    port map (
            O => \N__30713\,
            I => \N__30691\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__30710\,
            I => \N__30688\
        );

    \I__5410\ : InMux
    port map (
            O => \N__30709\,
            I => \N__30685\
        );

    \I__5409\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30682\
        );

    \I__5408\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30679\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30706\,
            I => \N__30676\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30673\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30666\
        );

    \I__5404\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30666\
        );

    \I__5403\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30666\
        );

    \I__5402\ : Sp12to4
    port map (
            O => \N__30697\,
            I => \N__30661\
        );

    \I__5401\ : Span12Mux_v
    port map (
            O => \N__30694\,
            I => \N__30661\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__30691\,
            I => \N__30654\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__30688\,
            I => \N__30654\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__30685\,
            I => \N__30654\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__30682\,
            I => \DTRIG_N_918_adj_1451\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__30679\,
            I => \DTRIG_N_918_adj_1451\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__30676\,
            I => \DTRIG_N_918_adj_1451\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__30673\,
            I => \DTRIG_N_918_adj_1451\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__30666\,
            I => \DTRIG_N_918_adj_1451\
        );

    \I__5392\ : Odrv12
    port map (
            O => \N__30661\,
            I => \DTRIG_N_918_adj_1451\
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__30654\,
            I => \DTRIG_N_918_adj_1451\
        );

    \I__5390\ : SRMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__5387\ : Span4Mux_h
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__5386\ : Span4Mux_v
    port map (
            O => \N__30627\,
            I => \N__30624\
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__30624\,
            I => \ADC_VAC.n14844\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30621\,
            I => n19741
        );

    \I__5383\ : InMux
    port map (
            O => \N__30618\,
            I => n19742
        );

    \I__5382\ : InMux
    port map (
            O => \N__30615\,
            I => n19743
        );

    \I__5381\ : InMux
    port map (
            O => \N__30612\,
            I => n19744
        );

    \I__5380\ : InMux
    port map (
            O => \N__30609\,
            I => n19745
        );

    \I__5379\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30602\
        );

    \I__5378\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30599\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__30602\,
            I => clk_cnt_0
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__30599\,
            I => clk_cnt_0
        );

    \I__5375\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30590\
        );

    \I__5374\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30587\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__30590\,
            I => clk_cnt_4
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__30587\,
            I => clk_cnt_4
        );

    \I__5371\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30578\
        );

    \I__5370\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30575\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30578\,
            I => clk_cnt_2
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__30575\,
            I => clk_cnt_2
        );

    \I__5367\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30566\
        );

    \I__5366\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30563\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__30566\,
            I => clk_cnt_1
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__30563\,
            I => clk_cnt_1
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__30558\,
            I => \n6_cascade_\
        );

    \I__5362\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30551\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30548\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__30551\,
            I => clk_cnt_3
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__30548\,
            I => clk_cnt_3
        );

    \I__5358\ : SRMux
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30537\
        );

    \I__5356\ : Sp12to4
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__5355\ : Odrv12
    port map (
            O => \N__30534\,
            I => n14714
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__30531\,
            I => \n14714_cascade_\
        );

    \I__5353\ : ClkMux
    port map (
            O => \N__30528\,
            I => \N__30522\
        );

    \I__5352\ : ClkMux
    port map (
            O => \N__30527\,
            I => \N__30519\
        );

    \I__5351\ : ClkMux
    port map (
            O => \N__30526\,
            I => \N__30514\
        );

    \I__5350\ : ClkMux
    port map (
            O => \N__30525\,
            I => \N__30510\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__30522\,
            I => \N__30501\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30501\
        );

    \I__5347\ : ClkMux
    port map (
            O => \N__30518\,
            I => \N__30498\
        );

    \I__5346\ : ClkMux
    port map (
            O => \N__30517\,
            I => \N__30495\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__30514\,
            I => \N__30489\
        );

    \I__5344\ : ClkMux
    port map (
            O => \N__30513\,
            I => \N__30486\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__30510\,
            I => \N__30483\
        );

    \I__5342\ : ClkMux
    port map (
            O => \N__30509\,
            I => \N__30480\
        );

    \I__5341\ : ClkMux
    port map (
            O => \N__30508\,
            I => \N__30477\
        );

    \I__5340\ : ClkMux
    port map (
            O => \N__30507\,
            I => \N__30473\
        );

    \I__5339\ : ClkMux
    port map (
            O => \N__30506\,
            I => \N__30469\
        );

    \I__5338\ : Span4Mux_v
    port map (
            O => \N__30501\,
            I => \N__30460\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__30498\,
            I => \N__30460\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30460\
        );

    \I__5335\ : ClkMux
    port map (
            O => \N__30494\,
            I => \N__30456\
        );

    \I__5334\ : ClkMux
    port map (
            O => \N__30493\,
            I => \N__30453\
        );

    \I__5333\ : ClkMux
    port map (
            O => \N__30492\,
            I => \N__30450\
        );

    \I__5332\ : Span4Mux_v
    port map (
            O => \N__30489\,
            I => \N__30446\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__30486\,
            I => \N__30443\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__30483\,
            I => \N__30438\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__30480\,
            I => \N__30438\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__30477\,
            I => \N__30435\
        );

    \I__5327\ : ClkMux
    port map (
            O => \N__30476\,
            I => \N__30432\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30473\,
            I => \N__30429\
        );

    \I__5325\ : ClkMux
    port map (
            O => \N__30472\,
            I => \N__30426\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__30469\,
            I => \N__30423\
        );

    \I__5323\ : ClkMux
    port map (
            O => \N__30468\,
            I => \N__30420\
        );

    \I__5322\ : ClkMux
    port map (
            O => \N__30467\,
            I => \N__30417\
        );

    \I__5321\ : Span4Mux_v
    port map (
            O => \N__30460\,
            I => \N__30413\
        );

    \I__5320\ : ClkMux
    port map (
            O => \N__30459\,
            I => \N__30410\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__30456\,
            I => \N__30403\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30453\,
            I => \N__30403\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__30450\,
            I => \N__30403\
        );

    \I__5316\ : ClkMux
    port map (
            O => \N__30449\,
            I => \N__30400\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__30446\,
            I => \N__30395\
        );

    \I__5314\ : Span4Mux_v
    port map (
            O => \N__30443\,
            I => \N__30395\
        );

    \I__5313\ : Span4Mux_v
    port map (
            O => \N__30438\,
            I => \N__30392\
        );

    \I__5312\ : Span4Mux_h
    port map (
            O => \N__30435\,
            I => \N__30387\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__30432\,
            I => \N__30387\
        );

    \I__5310\ : Span4Mux_v
    port map (
            O => \N__30429\,
            I => \N__30382\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__30426\,
            I => \N__30382\
        );

    \I__5308\ : Span4Mux_v
    port map (
            O => \N__30423\,
            I => \N__30375\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__30420\,
            I => \N__30375\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__30417\,
            I => \N__30375\
        );

    \I__5305\ : ClkMux
    port map (
            O => \N__30416\,
            I => \N__30372\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__30413\,
            I => \N__30369\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__30410\,
            I => \N__30362\
        );

    \I__5302\ : Sp12to4
    port map (
            O => \N__30403\,
            I => \N__30362\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__30400\,
            I => \N__30362\
        );

    \I__5300\ : Span4Mux_h
    port map (
            O => \N__30395\,
            I => \N__30359\
        );

    \I__5299\ : Span4Mux_h
    port map (
            O => \N__30392\,
            I => \N__30354\
        );

    \I__5298\ : Span4Mux_h
    port map (
            O => \N__30387\,
            I => \N__30354\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__30382\,
            I => \N__30347\
        );

    \I__5296\ : Span4Mux_v
    port map (
            O => \N__30375\,
            I => \N__30347\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__30372\,
            I => \N__30347\
        );

    \I__5294\ : Sp12to4
    port map (
            O => \N__30369\,
            I => \N__30341\
        );

    \I__5293\ : Span12Mux_v
    port map (
            O => \N__30362\,
            I => \N__30341\
        );

    \I__5292\ : Span4Mux_v
    port map (
            O => \N__30359\,
            I => \N__30336\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__30354\,
            I => \N__30336\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__30347\,
            I => \N__30333\
        );

    \I__5289\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30330\
        );

    \I__5288\ : Odrv12
    port map (
            O => \N__30341\,
            I => \clk_RTD\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__30336\,
            I => \clk_RTD\
        );

    \I__5286\ : Odrv4
    port map (
            O => \N__30333\,
            I => \clk_RTD\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__30330\,
            I => \clk_RTD\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30317\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30314\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__30317\,
            I => dds0_mclkcnt_3
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__30314\,
            I => dds0_mclkcnt_3
        );

    \I__5280\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30303\
        );

    \I__5279\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30299\
        );

    \I__5278\ : InMux
    port map (
            O => \N__30307\,
            I => \N__30290\
        );

    \I__5277\ : InMux
    port map (
            O => \N__30306\,
            I => \N__30290\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__30303\,
            I => \N__30287\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__30302\,
            I => \N__30282\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__30299\,
            I => \N__30278\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__30298\,
            I => \N__30275\
        );

    \I__5272\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30267\
        );

    \I__5271\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30267\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30264\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__30290\,
            I => \N__30259\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__30287\,
            I => \N__30259\
        );

    \I__5267\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30250\
        );

    \I__5266\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30250\
        );

    \I__5265\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30250\
        );

    \I__5264\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30250\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__30278\,
            I => \N__30247\
        );

    \I__5262\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30244\
        );

    \I__5261\ : InMux
    port map (
            O => \N__30274\,
            I => \N__30239\
        );

    \I__5260\ : InMux
    port map (
            O => \N__30273\,
            I => \N__30239\
        );

    \I__5259\ : InMux
    port map (
            O => \N__30272\,
            I => \N__30236\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30233\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__30264\,
            I => \N__30226\
        );

    \I__5256\ : Span4Mux_v
    port map (
            O => \N__30259\,
            I => \N__30226\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__30250\,
            I => \N__30226\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__30247\,
            I => \eis_end_N_724\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__30244\,
            I => \eis_end_N_724\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__30239\,
            I => \eis_end_N_724\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__30236\,
            I => \eis_end_N_724\
        );

    \I__5250\ : Odrv12
    port map (
            O => \N__30233\,
            I => \eis_end_N_724\
        );

    \I__5249\ : Odrv4
    port map (
            O => \N__30226\,
            I => \eis_end_N_724\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__30213\,
            I => \ADC_VDC.n10119_cascade_\
        );

    \I__5247\ : CEMux
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__30207\,
            I => \ADC_VDC.n12807\
        );

    \I__5245\ : InMux
    port map (
            O => \N__30204\,
            I => \bfn_12_4_0_\
        );

    \I__5244\ : InMux
    port map (
            O => \N__30201\,
            I => n19739
        );

    \I__5243\ : InMux
    port map (
            O => \N__30198\,
            I => n19740
        );

    \I__5242\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30192\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__30192\,
            I => \N__30188\
        );

    \I__5240\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30185\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__30188\,
            I => n20915
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__30185\,
            I => n20915
        );

    \I__5237\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30177\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__30177\,
            I => \N__30174\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__30174\,
            I => n20985
        );

    \I__5234\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30167\
        );

    \I__5233\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30164\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__30167\,
            I => n16571
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__30164\,
            I => n16571
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__30159\,
            I => \n13_cascade_\
        );

    \I__5229\ : InMux
    port map (
            O => \N__30156\,
            I => \N__30153\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__30153\,
            I => n21337
        );

    \I__5227\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__30147\,
            I => \N__30144\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__30144\,
            I => n17507
        );

    \I__5224\ : CascadeMux
    port map (
            O => \N__30141\,
            I => \N__30136\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30128\
        );

    \I__5222\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30128\
        );

    \I__5221\ : InMux
    port map (
            O => \N__30136\,
            I => \N__30128\
        );

    \I__5220\ : CascadeMux
    port map (
            O => \N__30135\,
            I => \N__30123\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__30128\,
            I => \N__30119\
        );

    \I__5218\ : InMux
    port map (
            O => \N__30127\,
            I => \N__30111\
        );

    \I__5217\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30108\
        );

    \I__5216\ : InMux
    port map (
            O => \N__30123\,
            I => \N__30103\
        );

    \I__5215\ : InMux
    port map (
            O => \N__30122\,
            I => \N__30103\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__30119\,
            I => \N__30100\
        );

    \I__5213\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30089\
        );

    \I__5212\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30089\
        );

    \I__5211\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30089\
        );

    \I__5210\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30089\
        );

    \I__5209\ : InMux
    port map (
            O => \N__30114\,
            I => \N__30089\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__30111\,
            I => eis_state_0
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__30108\,
            I => eis_state_0
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__30103\,
            I => eis_state_0
        );

    \I__5205\ : Odrv4
    port map (
            O => \N__30100\,
            I => eis_state_0
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__30089\,
            I => eis_state_0
        );

    \I__5203\ : CascadeMux
    port map (
            O => \N__30078\,
            I => \n11_adj_1621_cascade_\
        );

    \I__5202\ : CEMux
    port map (
            O => \N__30075\,
            I => \N__30071\
        );

    \I__5201\ : CEMux
    port map (
            O => \N__30074\,
            I => \N__30068\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__30071\,
            I => \N__30065\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__30068\,
            I => \N__30062\
        );

    \I__5198\ : Span4Mux_h
    port map (
            O => \N__30065\,
            I => \N__30059\
        );

    \I__5197\ : Sp12to4
    port map (
            O => \N__30062\,
            I => \N__30056\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__30059\,
            I => n11744
        );

    \I__5195\ : Odrv12
    port map (
            O => \N__30056\,
            I => n11744
        );

    \I__5194\ : InMux
    port map (
            O => \N__30051\,
            I => \N__30045\
        );

    \I__5193\ : InMux
    port map (
            O => \N__30050\,
            I => \N__30045\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__30045\,
            I => eis_end
        );

    \I__5191\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30039\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__30039\,
            I => n26_adj_1530
        );

    \I__5189\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30033\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__30033\,
            I => n21234
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__30030\,
            I => \N__30027\
        );

    \I__5186\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30024\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__30024\,
            I => n21
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__30021\,
            I => \n30_adj_1604_cascade_\
        );

    \I__5183\ : InMux
    port map (
            O => \N__30018\,
            I => \N__30014\
        );

    \I__5182\ : InMux
    port map (
            O => \N__30017\,
            I => \N__30011\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__30014\,
            I => n31
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__30011\,
            I => n31
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__30006\,
            I => \N__30003\
        );

    \I__5178\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29997\
        );

    \I__5177\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29990\
        );

    \I__5176\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29987\
        );

    \I__5175\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29984\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29997\,
            I => \N__29981\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__29996\,
            I => \N__29978\
        );

    \I__5172\ : CascadeMux
    port map (
            O => \N__29995\,
            I => \N__29975\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29968\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29968\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29960\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__29987\,
            I => \N__29960\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__29984\,
            I => \N__29960\
        );

    \I__5166\ : Span4Mux_h
    port map (
            O => \N__29981\,
            I => \N__29956\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29953\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29948\
        );

    \I__5163\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29948\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29945\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29968\,
            I => \N__29942\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29939\
        );

    \I__5159\ : Span4Mux_v
    port map (
            O => \N__29960\,
            I => \N__29936\
        );

    \I__5158\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29933\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__29956\,
            I => \DTRIG_N_918\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__29953\,
            I => \DTRIG_N_918\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__29948\,
            I => \DTRIG_N_918\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29945\,
            I => \DTRIG_N_918\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__29942\,
            I => \DTRIG_N_918\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__29939\,
            I => \DTRIG_N_918\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__29936\,
            I => \DTRIG_N_918\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29933\,
            I => \DTRIG_N_918\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__29916\,
            I => \N__29913\
        );

    \I__5148\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29906\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29903\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29896\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29891\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29891\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__29906\,
            I => \N__29887\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__29903\,
            I => \N__29884\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29902\,
            I => \N__29879\
        );

    \I__5140\ : InMux
    port map (
            O => \N__29901\,
            I => \N__29874\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29874\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29899\,
            I => \N__29871\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__29896\,
            I => \N__29866\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29891\,
            I => \N__29866\
        );

    \I__5135\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29863\
        );

    \I__5134\ : Span4Mux_v
    port map (
            O => \N__29887\,
            I => \N__29858\
        );

    \I__5133\ : Span4Mux_h
    port map (
            O => \N__29884\,
            I => \N__29858\
        );

    \I__5132\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29853\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29853\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__29879\,
            I => \N__29850\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__29874\,
            I => \N__29843\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__29871\,
            I => \N__29843\
        );

    \I__5127\ : Span4Mux_v
    port map (
            O => \N__29866\,
            I => \N__29843\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__29863\,
            I => adc_state_1
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__29858\,
            I => adc_state_1
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__29853\,
            I => adc_state_1
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__29850\,
            I => adc_state_1
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__29843\,
            I => adc_state_1
        );

    \I__5121\ : CascadeMux
    port map (
            O => \N__29832\,
            I => \n14_adj_1509_cascade_\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29826\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__29826\,
            I => n26_adj_1508
        );

    \I__5118\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29820\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29820\,
            I => n18_adj_1609
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__29817\,
            I => \N__29814\
        );

    \I__5115\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29811\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__29811\,
            I => \SIG_DDS.tmp_buf_9\
        );

    \I__5113\ : CascadeMux
    port map (
            O => \N__29808\,
            I => \N__29805\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29802\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__29802\,
            I => \SIG_DDS.tmp_buf_5\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29793\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29798\,
            I => \N__29793\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__29793\,
            I => n16554
        );

    \I__5107\ : CascadeMux
    port map (
            O => \N__29790\,
            I => \iac_raw_buf_N_736_cascade_\
        );

    \I__5106\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29784\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__29784\,
            I => n17_adj_1622
        );

    \I__5104\ : CascadeMux
    port map (
            O => \N__29781\,
            I => \n20826_cascade_\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__5102\ : CascadeBuf
    port map (
            O => \N__29775\,
            I => \N__29772\
        );

    \I__5101\ : CascadeMux
    port map (
            O => \N__29772\,
            I => \N__29769\
        );

    \I__5100\ : CascadeBuf
    port map (
            O => \N__29769\,
            I => \N__29766\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__29766\,
            I => \N__29763\
        );

    \I__5098\ : CascadeBuf
    port map (
            O => \N__29763\,
            I => \N__29760\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__29760\,
            I => \N__29757\
        );

    \I__5096\ : CascadeBuf
    port map (
            O => \N__29757\,
            I => \N__29754\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__29754\,
            I => \N__29751\
        );

    \I__5094\ : CascadeBuf
    port map (
            O => \N__29751\,
            I => \N__29748\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__29748\,
            I => \N__29745\
        );

    \I__5092\ : CascadeBuf
    port map (
            O => \N__29745\,
            I => \N__29742\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__29742\,
            I => \N__29739\
        );

    \I__5090\ : CascadeBuf
    port map (
            O => \N__29739\,
            I => \N__29736\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__29736\,
            I => \N__29732\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__29735\,
            I => \N__29729\
        );

    \I__5087\ : CascadeBuf
    port map (
            O => \N__29732\,
            I => \N__29726\
        );

    \I__5086\ : CascadeBuf
    port map (
            O => \N__29729\,
            I => \N__29723\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__29726\,
            I => \N__29720\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__29723\,
            I => \N__29717\
        );

    \I__5083\ : CascadeBuf
    port map (
            O => \N__29720\,
            I => \N__29714\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29711\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__29714\,
            I => \N__29708\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29705\
        );

    \I__5079\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29702\
        );

    \I__5078\ : Sp12to4
    port map (
            O => \N__29705\,
            I => \N__29698\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__29702\,
            I => \N__29695\
        );

    \I__5076\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29692\
        );

    \I__5075\ : Span12Mux_h
    port map (
            O => \N__29698\,
            I => \N__29687\
        );

    \I__5074\ : Span12Mux_h
    port map (
            O => \N__29695\,
            I => \N__29687\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__29692\,
            I => data_count_7
        );

    \I__5072\ : Odrv12
    port map (
            O => \N__29687\,
            I => data_count_7
        );

    \I__5071\ : InMux
    port map (
            O => \N__29682\,
            I => n19592
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__29679\,
            I => \N__29676\
        );

    \I__5069\ : CascadeBuf
    port map (
            O => \N__29676\,
            I => \N__29673\
        );

    \I__5068\ : CascadeMux
    port map (
            O => \N__29673\,
            I => \N__29670\
        );

    \I__5067\ : CascadeBuf
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__29667\,
            I => \N__29664\
        );

    \I__5065\ : CascadeBuf
    port map (
            O => \N__29664\,
            I => \N__29661\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__29661\,
            I => \N__29658\
        );

    \I__5063\ : CascadeBuf
    port map (
            O => \N__29658\,
            I => \N__29655\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__29655\,
            I => \N__29652\
        );

    \I__5061\ : CascadeBuf
    port map (
            O => \N__29652\,
            I => \N__29649\
        );

    \I__5060\ : CascadeMux
    port map (
            O => \N__29649\,
            I => \N__29646\
        );

    \I__5059\ : CascadeBuf
    port map (
            O => \N__29646\,
            I => \N__29643\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__29643\,
            I => \N__29640\
        );

    \I__5057\ : CascadeBuf
    port map (
            O => \N__29640\,
            I => \N__29637\
        );

    \I__5056\ : CascadeMux
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__5055\ : CascadeBuf
    port map (
            O => \N__29634\,
            I => \N__29630\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__29633\,
            I => \N__29627\
        );

    \I__5053\ : CascadeMux
    port map (
            O => \N__29630\,
            I => \N__29624\
        );

    \I__5052\ : CascadeBuf
    port map (
            O => \N__29627\,
            I => \N__29621\
        );

    \I__5051\ : CascadeBuf
    port map (
            O => \N__29624\,
            I => \N__29618\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__29621\,
            I => \N__29615\
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__29618\,
            I => \N__29612\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29609\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29606\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__29609\,
            I => \N__29603\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__29606\,
            I => \N__29600\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__29603\,
            I => \N__29597\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__29600\,
            I => \N__29594\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__29597\,
            I => \N__29590\
        );

    \I__5041\ : Sp12to4
    port map (
            O => \N__29594\,
            I => \N__29587\
        );

    \I__5040\ : InMux
    port map (
            O => \N__29593\,
            I => \N__29584\
        );

    \I__5039\ : Sp12to4
    port map (
            O => \N__29590\,
            I => \N__29579\
        );

    \I__5038\ : Span12Mux_h
    port map (
            O => \N__29587\,
            I => \N__29579\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__29584\,
            I => data_count_8
        );

    \I__5036\ : Odrv12
    port map (
            O => \N__29579\,
            I => data_count_8
        );

    \I__5035\ : InMux
    port map (
            O => \N__29574\,
            I => \bfn_11_14_0_\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29571\,
            I => n19594
        );

    \I__5033\ : CascadeMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__5032\ : CascadeBuf
    port map (
            O => \N__29565\,
            I => \N__29562\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__29562\,
            I => \N__29559\
        );

    \I__5030\ : CascadeBuf
    port map (
            O => \N__29559\,
            I => \N__29556\
        );

    \I__5029\ : CascadeMux
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__5028\ : CascadeBuf
    port map (
            O => \N__29553\,
            I => \N__29550\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__29550\,
            I => \N__29547\
        );

    \I__5026\ : CascadeBuf
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__5025\ : CascadeMux
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__5024\ : CascadeBuf
    port map (
            O => \N__29541\,
            I => \N__29538\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__5022\ : CascadeBuf
    port map (
            O => \N__29535\,
            I => \N__29532\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__29532\,
            I => \N__29529\
        );

    \I__5020\ : CascadeBuf
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__5018\ : CascadeBuf
    port map (
            O => \N__29523\,
            I => \N__29519\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__29522\,
            I => \N__29516\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__29519\,
            I => \N__29513\
        );

    \I__5015\ : CascadeBuf
    port map (
            O => \N__29516\,
            I => \N__29510\
        );

    \I__5014\ : CascadeBuf
    port map (
            O => \N__29513\,
            I => \N__29507\
        );

    \I__5013\ : CascadeMux
    port map (
            O => \N__29510\,
            I => \N__29504\
        );

    \I__5012\ : CascadeMux
    port map (
            O => \N__29507\,
            I => \N__29501\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29498\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29501\,
            I => \N__29495\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__29498\,
            I => \N__29492\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29489\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__29492\,
            I => \N__29486\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__29489\,
            I => \N__29483\
        );

    \I__5005\ : Sp12to4
    port map (
            O => \N__29486\,
            I => \N__29479\
        );

    \I__5004\ : Sp12to4
    port map (
            O => \N__29483\,
            I => \N__29476\
        );

    \I__5003\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29473\
        );

    \I__5002\ : Span12Mux_h
    port map (
            O => \N__29479\,
            I => \N__29468\
        );

    \I__5001\ : Span12Mux_h
    port map (
            O => \N__29476\,
            I => \N__29468\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__29473\,
            I => data_count_9
        );

    \I__4999\ : Odrv12
    port map (
            O => \N__29468\,
            I => data_count_9
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__29463\,
            I => \N__29460\
        );

    \I__4997\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29457\,
            I => \SIG_DDS.tmp_buf_10\
        );

    \I__4995\ : CascadeMux
    port map (
            O => \N__29454\,
            I => \N__29450\
        );

    \I__4994\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29446\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29441\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29441\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__29446\,
            I => buf_dds0_5
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__29441\,
            I => buf_dds0_5
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__29436\,
            I => \N__29433\
        );

    \I__4988\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29425\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29429\,
            I => \N__29420\
        );

    \I__4985\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29420\
        );

    \I__4984\ : Odrv12
    port map (
            O => \N__29425\,
            I => buf_dds0_14
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__29420\,
            I => buf_dds0_14
        );

    \I__4982\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__29412\,
            I => \SIG_DDS.tmp_buf_13\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__29409\,
            I => \N__29406\
        );

    \I__4979\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29403\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__29403\,
            I => \SIG_DDS.tmp_buf_11\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__29400\,
            I => \N__29397\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29394\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__29394\,
            I => \SIG_DDS.tmp_buf_12\
        );

    \I__4974\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29388\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__29388\,
            I => \CLK_DDS.tmp_buf_8\
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__29385\,
            I => \N__29382\
        );

    \I__4971\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29379\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__29379\,
            I => \CLK_DDS.tmp_buf_9\
        );

    \I__4969\ : CascadeMux
    port map (
            O => \N__29376\,
            I => \N__29373\
        );

    \I__4968\ : CascadeBuf
    port map (
            O => \N__29373\,
            I => \N__29370\
        );

    \I__4967\ : CascadeMux
    port map (
            O => \N__29370\,
            I => \N__29367\
        );

    \I__4966\ : CascadeBuf
    port map (
            O => \N__29367\,
            I => \N__29364\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__29364\,
            I => \N__29361\
        );

    \I__4964\ : CascadeBuf
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__29358\,
            I => \N__29355\
        );

    \I__4962\ : CascadeBuf
    port map (
            O => \N__29355\,
            I => \N__29352\
        );

    \I__4961\ : CascadeMux
    port map (
            O => \N__29352\,
            I => \N__29349\
        );

    \I__4960\ : CascadeBuf
    port map (
            O => \N__29349\,
            I => \N__29346\
        );

    \I__4959\ : CascadeMux
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__4958\ : CascadeBuf
    port map (
            O => \N__29343\,
            I => \N__29340\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__29340\,
            I => \N__29337\
        );

    \I__4956\ : CascadeBuf
    port map (
            O => \N__29337\,
            I => \N__29334\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__4954\ : CascadeBuf
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__29328\,
            I => \N__29324\
        );

    \I__4952\ : CascadeMux
    port map (
            O => \N__29327\,
            I => \N__29321\
        );

    \I__4951\ : CascadeBuf
    port map (
            O => \N__29324\,
            I => \N__29318\
        );

    \I__4950\ : CascadeBuf
    port map (
            O => \N__29321\,
            I => \N__29315\
        );

    \I__4949\ : CascadeMux
    port map (
            O => \N__29318\,
            I => \N__29312\
        );

    \I__4948\ : CascadeMux
    port map (
            O => \N__29315\,
            I => \N__29309\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29306\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29303\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__29306\,
            I => \N__29300\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29303\,
            I => \N__29297\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__29300\,
            I => \N__29294\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__29297\,
            I => \N__29290\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__29294\,
            I => \N__29287\
        );

    \I__4940\ : CascadeMux
    port map (
            O => \N__29293\,
            I => \N__29284\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__29290\,
            I => \N__29281\
        );

    \I__4938\ : Span4Mux_h
    port map (
            O => \N__29287\,
            I => \N__29278\
        );

    \I__4937\ : InMux
    port map (
            O => \N__29284\,
            I => \N__29275\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__29281\,
            I => \N__29270\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__29278\,
            I => \N__29270\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__29275\,
            I => data_count_0
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__29270\,
            I => data_count_0
        );

    \I__4932\ : CascadeMux
    port map (
            O => \N__29265\,
            I => \N__29262\
        );

    \I__4931\ : CascadeBuf
    port map (
            O => \N__29262\,
            I => \N__29259\
        );

    \I__4930\ : CascadeMux
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__4929\ : CascadeBuf
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__4927\ : CascadeBuf
    port map (
            O => \N__29250\,
            I => \N__29247\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__29247\,
            I => \N__29244\
        );

    \I__4925\ : CascadeBuf
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__29241\,
            I => \N__29238\
        );

    \I__4923\ : CascadeBuf
    port map (
            O => \N__29238\,
            I => \N__29235\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__4921\ : CascadeBuf
    port map (
            O => \N__29232\,
            I => \N__29229\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__29229\,
            I => \N__29226\
        );

    \I__4919\ : CascadeBuf
    port map (
            O => \N__29226\,
            I => \N__29223\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__29223\,
            I => \N__29220\
        );

    \I__4917\ : CascadeBuf
    port map (
            O => \N__29220\,
            I => \N__29216\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__29219\,
            I => \N__29213\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__29216\,
            I => \N__29210\
        );

    \I__4914\ : CascadeBuf
    port map (
            O => \N__29213\,
            I => \N__29207\
        );

    \I__4913\ : CascadeBuf
    port map (
            O => \N__29210\,
            I => \N__29204\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__29207\,
            I => \N__29201\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__29204\,
            I => \N__29198\
        );

    \I__4910\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29195\
        );

    \I__4909\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29192\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29189\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__29192\,
            I => \N__29186\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__29189\,
            I => \N__29183\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__29186\,
            I => \N__29180\
        );

    \I__4904\ : Sp12to4
    port map (
            O => \N__29183\,
            I => \N__29176\
        );

    \I__4903\ : Sp12to4
    port map (
            O => \N__29180\,
            I => \N__29173\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29179\,
            I => \N__29170\
        );

    \I__4901\ : Span12Mux_v
    port map (
            O => \N__29176\,
            I => \N__29165\
        );

    \I__4900\ : Span12Mux_v
    port map (
            O => \N__29173\,
            I => \N__29165\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29170\,
            I => data_count_1
        );

    \I__4898\ : Odrv12
    port map (
            O => \N__29165\,
            I => data_count_1
        );

    \I__4897\ : InMux
    port map (
            O => \N__29160\,
            I => n19586
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__29157\,
            I => \N__29154\
        );

    \I__4895\ : CascadeBuf
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__4893\ : CascadeBuf
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__29145\,
            I => \N__29142\
        );

    \I__4891\ : CascadeBuf
    port map (
            O => \N__29142\,
            I => \N__29139\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__29139\,
            I => \N__29136\
        );

    \I__4889\ : CascadeBuf
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__4888\ : CascadeMux
    port map (
            O => \N__29133\,
            I => \N__29130\
        );

    \I__4887\ : CascadeBuf
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__4886\ : CascadeMux
    port map (
            O => \N__29127\,
            I => \N__29124\
        );

    \I__4885\ : CascadeBuf
    port map (
            O => \N__29124\,
            I => \N__29121\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__29121\,
            I => \N__29118\
        );

    \I__4883\ : CascadeBuf
    port map (
            O => \N__29118\,
            I => \N__29115\
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__29115\,
            I => \N__29112\
        );

    \I__4881\ : CascadeBuf
    port map (
            O => \N__29112\,
            I => \N__29109\
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__29109\,
            I => \N__29105\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__29108\,
            I => \N__29102\
        );

    \I__4878\ : CascadeBuf
    port map (
            O => \N__29105\,
            I => \N__29099\
        );

    \I__4877\ : CascadeBuf
    port map (
            O => \N__29102\,
            I => \N__29096\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__29099\,
            I => \N__29093\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__29096\,
            I => \N__29090\
        );

    \I__4874\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29087\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29084\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__29087\,
            I => \N__29081\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29078\
        );

    \I__4870\ : Span4Mux_v
    port map (
            O => \N__29081\,
            I => \N__29075\
        );

    \I__4869\ : Sp12to4
    port map (
            O => \N__29078\,
            I => \N__29071\
        );

    \I__4868\ : Sp12to4
    port map (
            O => \N__29075\,
            I => \N__29068\
        );

    \I__4867\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29065\
        );

    \I__4866\ : Span12Mux_v
    port map (
            O => \N__29071\,
            I => \N__29062\
        );

    \I__4865\ : Span12Mux_h
    port map (
            O => \N__29068\,
            I => \N__29059\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__29065\,
            I => data_count_2
        );

    \I__4863\ : Odrv12
    port map (
            O => \N__29062\,
            I => data_count_2
        );

    \I__4862\ : Odrv12
    port map (
            O => \N__29059\,
            I => data_count_2
        );

    \I__4861\ : InMux
    port map (
            O => \N__29052\,
            I => n19587
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__29049\,
            I => \N__29046\
        );

    \I__4859\ : CascadeBuf
    port map (
            O => \N__29046\,
            I => \N__29043\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__4857\ : CascadeBuf
    port map (
            O => \N__29040\,
            I => \N__29037\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__29037\,
            I => \N__29034\
        );

    \I__4855\ : CascadeBuf
    port map (
            O => \N__29034\,
            I => \N__29031\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__29031\,
            I => \N__29028\
        );

    \I__4853\ : CascadeBuf
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__29025\,
            I => \N__29022\
        );

    \I__4851\ : CascadeBuf
    port map (
            O => \N__29022\,
            I => \N__29019\
        );

    \I__4850\ : CascadeMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__4849\ : CascadeBuf
    port map (
            O => \N__29016\,
            I => \N__29013\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__29013\,
            I => \N__29010\
        );

    \I__4847\ : CascadeBuf
    port map (
            O => \N__29010\,
            I => \N__29007\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__29007\,
            I => \N__29004\
        );

    \I__4845\ : CascadeBuf
    port map (
            O => \N__29004\,
            I => \N__29001\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__29001\,
            I => \N__28998\
        );

    \I__4843\ : CascadeBuf
    port map (
            O => \N__28998\,
            I => \N__28994\
        );

    \I__4842\ : CascadeMux
    port map (
            O => \N__28997\,
            I => \N__28991\
        );

    \I__4841\ : CascadeMux
    port map (
            O => \N__28994\,
            I => \N__28988\
        );

    \I__4840\ : CascadeBuf
    port map (
            O => \N__28991\,
            I => \N__28985\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28982\
        );

    \I__4838\ : CascadeMux
    port map (
            O => \N__28985\,
            I => \N__28979\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28976\
        );

    \I__4836\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28973\
        );

    \I__4835\ : Span4Mux_v
    port map (
            O => \N__28976\,
            I => \N__28970\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28973\,
            I => \N__28966\
        );

    \I__4833\ : Sp12to4
    port map (
            O => \N__28970\,
            I => \N__28963\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28960\
        );

    \I__4831\ : Span12Mux_v
    port map (
            O => \N__28966\,
            I => \N__28957\
        );

    \I__4830\ : Span12Mux_h
    port map (
            O => \N__28963\,
            I => \N__28954\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28960\,
            I => data_count_3
        );

    \I__4828\ : Odrv12
    port map (
            O => \N__28957\,
            I => data_count_3
        );

    \I__4827\ : Odrv12
    port map (
            O => \N__28954\,
            I => data_count_3
        );

    \I__4826\ : InMux
    port map (
            O => \N__28947\,
            I => n19588
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__4824\ : CascadeBuf
    port map (
            O => \N__28941\,
            I => \N__28938\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__28938\,
            I => \N__28935\
        );

    \I__4822\ : CascadeBuf
    port map (
            O => \N__28935\,
            I => \N__28932\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__28932\,
            I => \N__28929\
        );

    \I__4820\ : CascadeBuf
    port map (
            O => \N__28929\,
            I => \N__28926\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__28926\,
            I => \N__28923\
        );

    \I__4818\ : CascadeBuf
    port map (
            O => \N__28923\,
            I => \N__28920\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__28920\,
            I => \N__28917\
        );

    \I__4816\ : CascadeBuf
    port map (
            O => \N__28917\,
            I => \N__28914\
        );

    \I__4815\ : CascadeMux
    port map (
            O => \N__28914\,
            I => \N__28911\
        );

    \I__4814\ : CascadeBuf
    port map (
            O => \N__28911\,
            I => \N__28908\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__28908\,
            I => \N__28905\
        );

    \I__4812\ : CascadeBuf
    port map (
            O => \N__28905\,
            I => \N__28902\
        );

    \I__4811\ : CascadeMux
    port map (
            O => \N__28902\,
            I => \N__28899\
        );

    \I__4810\ : CascadeBuf
    port map (
            O => \N__28899\,
            I => \N__28895\
        );

    \I__4809\ : CascadeMux
    port map (
            O => \N__28898\,
            I => \N__28892\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__28895\,
            I => \N__28889\
        );

    \I__4807\ : CascadeBuf
    port map (
            O => \N__28892\,
            I => \N__28886\
        );

    \I__4806\ : CascadeBuf
    port map (
            O => \N__28889\,
            I => \N__28883\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__28886\,
            I => \N__28880\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__28883\,
            I => \N__28877\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28874\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28871\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28868\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__28871\,
            I => \N__28865\
        );

    \I__4799\ : Span4Mux_h
    port map (
            O => \N__28868\,
            I => \N__28862\
        );

    \I__4798\ : Span4Mux_v
    port map (
            O => \N__28865\,
            I => \N__28859\
        );

    \I__4797\ : Span4Mux_v
    port map (
            O => \N__28862\,
            I => \N__28855\
        );

    \I__4796\ : Span4Mux_v
    port map (
            O => \N__28859\,
            I => \N__28852\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28849\
        );

    \I__4794\ : Span4Mux_h
    port map (
            O => \N__28855\,
            I => \N__28846\
        );

    \I__4793\ : Sp12to4
    port map (
            O => \N__28852\,
            I => \N__28843\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__28849\,
            I => data_count_4
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__28846\,
            I => data_count_4
        );

    \I__4790\ : Odrv12
    port map (
            O => \N__28843\,
            I => data_count_4
        );

    \I__4789\ : InMux
    port map (
            O => \N__28836\,
            I => n19589
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__28833\,
            I => \N__28830\
        );

    \I__4787\ : CascadeBuf
    port map (
            O => \N__28830\,
            I => \N__28827\
        );

    \I__4786\ : CascadeMux
    port map (
            O => \N__28827\,
            I => \N__28824\
        );

    \I__4785\ : CascadeBuf
    port map (
            O => \N__28824\,
            I => \N__28821\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__28821\,
            I => \N__28818\
        );

    \I__4783\ : CascadeBuf
    port map (
            O => \N__28818\,
            I => \N__28815\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__28815\,
            I => \N__28812\
        );

    \I__4781\ : CascadeBuf
    port map (
            O => \N__28812\,
            I => \N__28809\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__28809\,
            I => \N__28806\
        );

    \I__4779\ : CascadeBuf
    port map (
            O => \N__28806\,
            I => \N__28803\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__28803\,
            I => \N__28800\
        );

    \I__4777\ : CascadeBuf
    port map (
            O => \N__28800\,
            I => \N__28797\
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__28797\,
            I => \N__28794\
        );

    \I__4775\ : CascadeBuf
    port map (
            O => \N__28794\,
            I => \N__28791\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__28791\,
            I => \N__28787\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__28790\,
            I => \N__28784\
        );

    \I__4772\ : CascadeBuf
    port map (
            O => \N__28787\,
            I => \N__28781\
        );

    \I__4771\ : CascadeBuf
    port map (
            O => \N__28784\,
            I => \N__28778\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__28781\,
            I => \N__28775\
        );

    \I__4769\ : CascadeMux
    port map (
            O => \N__28778\,
            I => \N__28772\
        );

    \I__4768\ : CascadeBuf
    port map (
            O => \N__28775\,
            I => \N__28769\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28772\,
            I => \N__28766\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__28769\,
            I => \N__28763\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__28766\,
            I => \N__28760\
        );

    \I__4764\ : InMux
    port map (
            O => \N__28763\,
            I => \N__28757\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__28760\,
            I => \N__28754\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__28757\,
            I => \N__28750\
        );

    \I__4761\ : Span4Mux_v
    port map (
            O => \N__28754\,
            I => \N__28747\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28744\
        );

    \I__4759\ : Sp12to4
    port map (
            O => \N__28750\,
            I => \N__28741\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__28747\,
            I => \N__28738\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__28744\,
            I => \N__28733\
        );

    \I__4756\ : Span12Mux_v
    port map (
            O => \N__28741\,
            I => \N__28733\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__28738\,
            I => data_count_5
        );

    \I__4754\ : Odrv12
    port map (
            O => \N__28733\,
            I => data_count_5
        );

    \I__4753\ : InMux
    port map (
            O => \N__28728\,
            I => n19590
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__28725\,
            I => \N__28722\
        );

    \I__4751\ : CascadeBuf
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__28719\,
            I => \N__28716\
        );

    \I__4749\ : CascadeBuf
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__4747\ : CascadeBuf
    port map (
            O => \N__28710\,
            I => \N__28707\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__28707\,
            I => \N__28704\
        );

    \I__4745\ : CascadeBuf
    port map (
            O => \N__28704\,
            I => \N__28701\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__28701\,
            I => \N__28698\
        );

    \I__4743\ : CascadeBuf
    port map (
            O => \N__28698\,
            I => \N__28695\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__28695\,
            I => \N__28692\
        );

    \I__4741\ : CascadeBuf
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__28689\,
            I => \N__28686\
        );

    \I__4739\ : CascadeBuf
    port map (
            O => \N__28686\,
            I => \N__28682\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__28685\,
            I => \N__28679\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__28682\,
            I => \N__28676\
        );

    \I__4736\ : CascadeBuf
    port map (
            O => \N__28679\,
            I => \N__28673\
        );

    \I__4735\ : CascadeBuf
    port map (
            O => \N__28676\,
            I => \N__28670\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__28673\,
            I => \N__28667\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__28670\,
            I => \N__28664\
        );

    \I__4732\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28661\
        );

    \I__4731\ : CascadeBuf
    port map (
            O => \N__28664\,
            I => \N__28658\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28661\,
            I => \N__28655\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__28658\,
            I => \N__28652\
        );

    \I__4728\ : Span4Mux_v
    port map (
            O => \N__28655\,
            I => \N__28649\
        );

    \I__4727\ : InMux
    port map (
            O => \N__28652\,
            I => \N__28646\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__28649\,
            I => \N__28642\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__28646\,
            I => \N__28639\
        );

    \I__4724\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28636\
        );

    \I__4723\ : Span4Mux_h
    port map (
            O => \N__28642\,
            I => \N__28633\
        );

    \I__4722\ : Span12Mux_v
    port map (
            O => \N__28639\,
            I => \N__28630\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__28636\,
            I => data_count_6
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__28633\,
            I => data_count_6
        );

    \I__4719\ : Odrv12
    port map (
            O => \N__28630\,
            I => data_count_6
        );

    \I__4718\ : InMux
    port map (
            O => \N__28623\,
            I => n19591
        );

    \I__4717\ : InMux
    port map (
            O => \N__28620\,
            I => n19770
        );

    \I__4716\ : InMux
    port map (
            O => \N__28617\,
            I => n19771
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__28614\,
            I => \N__28611\
        );

    \I__4714\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28603\
        );

    \I__4712\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28600\
        );

    \I__4711\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28597\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__28603\,
            I => \N__28594\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__28600\,
            I => \N__28591\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__28597\,
            I => buf_dds1_14
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__28594\,
            I => buf_dds1_14
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__28591\,
            I => buf_dds1_14
        );

    \I__4705\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28581\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__28581\,
            I => \CLK_DDS.tmp_buf_13\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__4702\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__28572\,
            I => \CLK_DDS.tmp_buf_14\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28566\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__28566\,
            I => \CLK_DDS.tmp_buf_0\
        );

    \I__4698\ : CascadeMux
    port map (
            O => \N__28563\,
            I => \N__28560\
        );

    \I__4697\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__28557\,
            I => \CLK_DDS.tmp_buf_1\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__28554\,
            I => \N__28551\
        );

    \I__4694\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28548\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__28548\,
            I => \CLK_DDS.tmp_buf_2\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__28545\,
            I => \N__28542\
        );

    \I__4691\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28539\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__28539\,
            I => \CLK_DDS.tmp_buf_3\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__4688\ : InMux
    port map (
            O => \N__28533\,
            I => \N__28530\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__28530\,
            I => \CLK_DDS.tmp_buf_4\
        );

    \I__4686\ : CascadeMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__4685\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__28521\,
            I => \CLK_DDS.tmp_buf_5\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28518\,
            I => \N__28515\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__28515\,
            I => \CLK_DDS.tmp_buf_6\
        );

    \I__4681\ : InMux
    port map (
            O => \N__28512\,
            I => n19761
        );

    \I__4680\ : InMux
    port map (
            O => \N__28509\,
            I => n19762
        );

    \I__4679\ : InMux
    port map (
            O => \N__28506\,
            I => n19763
        );

    \I__4678\ : InMux
    port map (
            O => \N__28503\,
            I => n19764
        );

    \I__4677\ : InMux
    port map (
            O => \N__28500\,
            I => \bfn_11_11_0_\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28497\,
            I => n19766
        );

    \I__4675\ : InMux
    port map (
            O => \N__28494\,
            I => n19767
        );

    \I__4674\ : InMux
    port map (
            O => \N__28491\,
            I => n19768
        );

    \I__4673\ : InMux
    port map (
            O => \N__28488\,
            I => n19769
        );

    \I__4672\ : InMux
    port map (
            O => \N__28485\,
            I => n19752
        );

    \I__4671\ : InMux
    port map (
            O => \N__28482\,
            I => n19753
        );

    \I__4670\ : InMux
    port map (
            O => \N__28479\,
            I => n19754
        );

    \I__4669\ : InMux
    port map (
            O => \N__28476\,
            I => n19755
        );

    \I__4668\ : InMux
    port map (
            O => \N__28473\,
            I => n19756
        );

    \I__4667\ : InMux
    port map (
            O => \N__28470\,
            I => \bfn_11_10_0_\
        );

    \I__4666\ : InMux
    port map (
            O => \N__28467\,
            I => n19758
        );

    \I__4665\ : InMux
    port map (
            O => \N__28464\,
            I => n19759
        );

    \I__4664\ : InMux
    port map (
            O => \N__28461\,
            I => n19760
        );

    \I__4663\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28448\
        );

    \I__4662\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28448\
        );

    \I__4661\ : InMux
    port map (
            O => \N__28456\,
            I => \N__28448\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28455\,
            I => \N__28445\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__28448\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28445\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__4657\ : CascadeMux
    port map (
            O => \N__28440\,
            I => \N__28435\
        );

    \I__4656\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28430\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28430\
        );

    \I__4654\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28427\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__28430\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__28427\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28406\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28406\
        );

    \I__4648\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28406\
        );

    \I__4647\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28406\
        );

    \I__4646\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28403\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__28406\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__28403\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__4643\ : CascadeMux
    port map (
            O => \N__28398\,
            I => \N__28394\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__28397\,
            I => \N__28391\
        );

    \I__4641\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28388\
        );

    \I__4640\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28384\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__28388\,
            I => \N__28381\
        );

    \I__4638\ : InMux
    port map (
            O => \N__28387\,
            I => \N__28378\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__28384\,
            I => cmd_rdadctmp_11
        );

    \I__4636\ : Odrv12
    port map (
            O => \N__28381\,
            I => cmd_rdadctmp_11
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__28378\,
            I => cmd_rdadctmp_11
        );

    \I__4634\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__28365\,
            I => \N__28362\
        );

    \I__4631\ : Sp12to4
    port map (
            O => \N__28362\,
            I => \N__28357\
        );

    \I__4630\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28352\
        );

    \I__4629\ : InMux
    port map (
            O => \N__28360\,
            I => \N__28352\
        );

    \I__4628\ : Odrv12
    port map (
            O => \N__28357\,
            I => buf_adcdata_vac_3
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__28352\,
            I => buf_adcdata_vac_3
        );

    \I__4626\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28343\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__28346\,
            I => \N__28340\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__28343\,
            I => \N__28337\
        );

    \I__4623\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__4622\ : Span4Mux_v
    port map (
            O => \N__28337\,
            I => \N__28328\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28328\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__28333\,
            I => \N__28325\
        );

    \I__4619\ : Span4Mux_h
    port map (
            O => \N__28328\,
            I => \N__28322\
        );

    \I__4618\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28319\
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__28322\,
            I => cmd_rdadctmp_10_adj_1440
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__28319\,
            I => cmd_rdadctmp_10_adj_1440
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__28314\,
            I => \N__28310\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__28313\,
            I => \N__28307\
        );

    \I__4613\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28299\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28299\
        );

    \I__4611\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28299\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__28299\,
            I => cmd_rdadctmp_11_adj_1439
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__28296\,
            I => \N__28293\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28289\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__28292\,
            I => \N__28286\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__28289\,
            I => \N__28283\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28279\
        );

    \I__4604\ : Span4Mux_h
    port map (
            O => \N__28283\,
            I => \N__28276\
        );

    \I__4603\ : InMux
    port map (
            O => \N__28282\,
            I => \N__28273\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__28279\,
            I => \N__28270\
        );

    \I__4601\ : Span4Mux_h
    port map (
            O => \N__28276\,
            I => \N__28267\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__28273\,
            I => cmd_rdadctmp_12_adj_1438
        );

    \I__4599\ : Odrv12
    port map (
            O => \N__28270\,
            I => cmd_rdadctmp_12_adj_1438
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__28267\,
            I => cmd_rdadctmp_12_adj_1438
        );

    \I__4597\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__28257\,
            I => n22_adj_1640
        );

    \I__4595\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28251\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__28251\,
            I => \N__28248\
        );

    \I__4593\ : Sp12to4
    port map (
            O => \N__28248\,
            I => \N__28245\
        );

    \I__4592\ : Span12Mux_h
    port map (
            O => \N__28245\,
            I => \N__28242\
        );

    \I__4591\ : Odrv12
    port map (
            O => \N__28242\,
            I => buf_data_iac_2
        );

    \I__4590\ : InMux
    port map (
            O => \N__28239\,
            I => \bfn_11_9_0_\
        );

    \I__4589\ : InMux
    port map (
            O => \N__28236\,
            I => n19750
        );

    \I__4588\ : InMux
    port map (
            O => \N__28233\,
            I => n19751
        );

    \I__4587\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28227\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__28227\,
            I => \N__28223\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__28226\,
            I => \N__28220\
        );

    \I__4584\ : Span4Mux_h
    port map (
            O => \N__28223\,
            I => \N__28217\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28214\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__28217\,
            I => buf_adcdata_vdc_2
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__28214\,
            I => buf_adcdata_vdc_2
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__28209\,
            I => \n19_adj_1639_cascade_\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28203\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__28203\,
            I => \N__28200\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__28200\,
            I => \N__28197\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__28197\,
            I => buf_data_iac_5
        );

    \I__4575\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28191\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__28191\,
            I => \N__28188\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__28188\,
            I => \N__28185\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__28185\,
            I => \N__28182\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__28182\,
            I => n22_adj_1630
        );

    \I__4570\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28176\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__28176\,
            I => \N__28173\
        );

    \I__4568\ : Span4Mux_v
    port map (
            O => \N__28173\,
            I => \N__28168\
        );

    \I__4567\ : InMux
    port map (
            O => \N__28172\,
            I => \N__28163\
        );

    \I__4566\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28163\
        );

    \I__4565\ : Sp12to4
    port map (
            O => \N__28168\,
            I => \N__28160\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__28163\,
            I => buf_adcdata_iac_2
        );

    \I__4563\ : Odrv12
    port map (
            O => \N__28160\,
            I => buf_adcdata_iac_2
        );

    \I__4562\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28148\
        );

    \I__4561\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28148\
        );

    \I__4560\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28145\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__28148\,
            I => cmd_rdadctmp_9
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__28145\,
            I => cmd_rdadctmp_9
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__28140\,
            I => \N__28135\
        );

    \I__4556\ : InMux
    port map (
            O => \N__28139\,
            I => \N__28128\
        );

    \I__4555\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28128\
        );

    \I__4554\ : InMux
    port map (
            O => \N__28135\,
            I => \N__28128\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__28128\,
            I => cmd_rdadctmp_10
        );

    \I__4552\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28119\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__28124\,
            I => \N__28109\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__28123\,
            I => \N__28105\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__28122\,
            I => \N__28100\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28094\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__28118\,
            I => \N__28088\
        );

    \I__4546\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28083\
        );

    \I__4545\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28083\
        );

    \I__4544\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28076\
        );

    \I__4543\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28076\
        );

    \I__4542\ : InMux
    port map (
            O => \N__28113\,
            I => \N__28076\
        );

    \I__4541\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28073\
        );

    \I__4540\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28070\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__28108\,
            I => \N__28067\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28056\
        );

    \I__4537\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28056\
        );

    \I__4536\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28056\
        );

    \I__4535\ : InMux
    port map (
            O => \N__28100\,
            I => \N__28051\
        );

    \I__4534\ : InMux
    port map (
            O => \N__28099\,
            I => \N__28051\
        );

    \I__4533\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28048\
        );

    \I__4532\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28042\
        );

    \I__4531\ : Span4Mux_h
    port map (
            O => \N__28094\,
            I => \N__28039\
        );

    \I__4530\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28036\
        );

    \I__4529\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28031\
        );

    \I__4528\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28028\
        );

    \I__4527\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28025\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__28083\,
            I => \N__28020\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__28076\,
            I => \N__28020\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__28073\,
            I => \N__28017\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__28070\,
            I => \N__28014\
        );

    \I__4522\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28009\
        );

    \I__4521\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28009\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__28065\,
            I => \N__28006\
        );

    \I__4519\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28002\
        );

    \I__4518\ : InMux
    port map (
            O => \N__28063\,
            I => \N__27999\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__28056\,
            I => \N__27996\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__28051\,
            I => \N__27991\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__28048\,
            I => \N__27991\
        );

    \I__4514\ : InMux
    port map (
            O => \N__28047\,
            I => \N__27984\
        );

    \I__4513\ : InMux
    port map (
            O => \N__28046\,
            I => \N__27984\
        );

    \I__4512\ : InMux
    port map (
            O => \N__28045\,
            I => \N__27984\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__28042\,
            I => \N__27979\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__28039\,
            I => \N__27979\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__27976\
        );

    \I__4508\ : InMux
    port map (
            O => \N__28035\,
            I => \N__27970\
        );

    \I__4507\ : InMux
    port map (
            O => \N__28034\,
            I => \N__27970\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__28031\,
            I => \N__27959\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__28028\,
            I => \N__27959\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__28025\,
            I => \N__27959\
        );

    \I__4503\ : Span4Mux_v
    port map (
            O => \N__28020\,
            I => \N__27959\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__28017\,
            I => \N__27959\
        );

    \I__4501\ : Sp12to4
    port map (
            O => \N__28014\,
            I => \N__27954\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__28009\,
            I => \N__27954\
        );

    \I__4499\ : InMux
    port map (
            O => \N__28006\,
            I => \N__27949\
        );

    \I__4498\ : InMux
    port map (
            O => \N__28005\,
            I => \N__27949\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__28002\,
            I => \N__27946\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__27999\,
            I => \N__27943\
        );

    \I__4495\ : Span4Mux_v
    port map (
            O => \N__27996\,
            I => \N__27938\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__27991\,
            I => \N__27938\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27931\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__27979\,
            I => \N__27931\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__27976\,
            I => \N__27931\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27928\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__27970\,
            I => \N__27923\
        );

    \I__4488\ : Span4Mux_v
    port map (
            O => \N__27959\,
            I => \N__27923\
        );

    \I__4487\ : Span12Mux_v
    port map (
            O => \N__27954\,
            I => \N__27920\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__27949\,
            I => \N__27911\
        );

    \I__4485\ : Span4Mux_h
    port map (
            O => \N__27946\,
            I => \N__27911\
        );

    \I__4484\ : Span4Mux_v
    port map (
            O => \N__27943\,
            I => \N__27911\
        );

    \I__4483\ : Span4Mux_v
    port map (
            O => \N__27938\,
            I => \N__27911\
        );

    \I__4482\ : Span4Mux_v
    port map (
            O => \N__27931\,
            I => \N__27908\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27928\,
            I => n12498
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__27923\,
            I => n12498
        );

    \I__4479\ : Odrv12
    port map (
            O => \N__27920\,
            I => n12498
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__27911\,
            I => n12498
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__27908\,
            I => n12498
        );

    \I__4476\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27894\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27894\,
            I => \N__27891\
        );

    \I__4474\ : Span4Mux_h
    port map (
            O => \N__27891\,
            I => \N__27888\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__27888\,
            I => \N__27883\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27878\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27878\
        );

    \I__4470\ : Span4Mux_h
    port map (
            O => \N__27883\,
            I => \N__27875\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__27878\,
            I => buf_adcdata_vac_2
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__27875\,
            I => buf_adcdata_vac_2
        );

    \I__4467\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27867\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27867\,
            I => \N__27863\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__27866\,
            I => \N__27860\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__27863\,
            I => \N__27857\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27854\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__27857\,
            I => buf_adcdata_vdc_3
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__27854\,
            I => buf_adcdata_vdc_3
        );

    \I__4460\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27846\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__27846\,
            I => \ADC_VDC.n21952\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27843\,
            I => \bfn_11_5_0_\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27840\,
            I => n19746
        );

    \I__4456\ : InMux
    port map (
            O => \N__27837\,
            I => n19747
        );

    \I__4455\ : InMux
    port map (
            O => \N__27834\,
            I => n19748
        );

    \I__4454\ : InMux
    port map (
            O => \N__27831\,
            I => n19749
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__27828\,
            I => \N__27825\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27817\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27817\
        );

    \I__4450\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27814\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27811\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__27817\,
            I => \N__27803\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27814\,
            I => \N__27803\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__27811\,
            I => \N__27803\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27800\
        );

    \I__4444\ : Span4Mux_v
    port map (
            O => \N__27803\,
            I => \N__27795\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__27800\,
            I => \N__27795\
        );

    \I__4442\ : Span4Mux_v
    port map (
            O => \N__27795\,
            I => \N__27792\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__27792\,
            I => \N__27789\
        );

    \I__4440\ : Sp12to4
    port map (
            O => \N__27789\,
            I => \N__27786\
        );

    \I__4439\ : Span12Mux_h
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__4438\ : Odrv12
    port map (
            O => \N__27783\,
            I => \ICE_SPI_SCLK\
        );

    \I__4437\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27777\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27777\,
            I => \comm_spi.n14596\
        );

    \I__4435\ : SRMux
    port map (
            O => \N__27774\,
            I => \N__27771\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27771\,
            I => \N__27768\
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__27768\,
            I => \comm_spi.iclk_N_762\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27762\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__27762\,
            I => n22255
        );

    \I__4430\ : SRMux
    port map (
            O => \N__27759\,
            I => \N__27753\
        );

    \I__4429\ : SRMux
    port map (
            O => \N__27758\,
            I => \N__27750\
        );

    \I__4428\ : SRMux
    port map (
            O => \N__27757\,
            I => \N__27745\
        );

    \I__4427\ : SRMux
    port map (
            O => \N__27756\,
            I => \N__27742\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27753\,
            I => \N__27737\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__27750\,
            I => \N__27737\
        );

    \I__4424\ : SRMux
    port map (
            O => \N__27749\,
            I => \N__27734\
        );

    \I__4423\ : SRMux
    port map (
            O => \N__27748\,
            I => \N__27731\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__27745\,
            I => \N__27726\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__27742\,
            I => \N__27723\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__27737\,
            I => \N__27716\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27716\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__27731\,
            I => \N__27716\
        );

    \I__4417\ : SRMux
    port map (
            O => \N__27730\,
            I => \N__27713\
        );

    \I__4416\ : SRMux
    port map (
            O => \N__27729\,
            I => \N__27710\
        );

    \I__4415\ : Span4Mux_v
    port map (
            O => \N__27726\,
            I => \N__27703\
        );

    \I__4414\ : Span4Mux_h
    port map (
            O => \N__27723\,
            I => \N__27700\
        );

    \I__4413\ : Span4Mux_v
    port map (
            O => \N__27716\,
            I => \N__27693\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__27713\,
            I => \N__27693\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27693\
        );

    \I__4410\ : SRMux
    port map (
            O => \N__27709\,
            I => \N__27690\
        );

    \I__4409\ : SRMux
    port map (
            O => \N__27708\,
            I => \N__27687\
        );

    \I__4408\ : SRMux
    port map (
            O => \N__27707\,
            I => \N__27684\
        );

    \I__4407\ : SRMux
    port map (
            O => \N__27706\,
            I => \N__27681\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__27703\,
            I => \N__27678\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__27700\,
            I => \N__27675\
        );

    \I__4404\ : Span4Mux_v
    port map (
            O => \N__27693\,
            I => \N__27668\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__27690\,
            I => \N__27668\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__27687\,
            I => \N__27668\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27663\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__27681\,
            I => \N__27663\
        );

    \I__4399\ : Span4Mux_v
    port map (
            O => \N__27678\,
            I => \N__27660\
        );

    \I__4398\ : Span4Mux_v
    port map (
            O => \N__27675\,
            I => \N__27657\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__27668\,
            I => \N__27652\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__27663\,
            I => \N__27652\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__27660\,
            I => \N__27649\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__27657\,
            I => \N__27646\
        );

    \I__4393\ : Sp12to4
    port map (
            O => \N__27652\,
            I => \N__27643\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__27649\,
            I => \iac_raw_buf_N_734\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__27646\,
            I => \iac_raw_buf_N_734\
        );

    \I__4390\ : Odrv12
    port map (
            O => \N__27643\,
            I => \iac_raw_buf_N_734\
        );

    \I__4389\ : IoInMux
    port map (
            O => \N__27636\,
            I => \N__27633\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__27633\,
            I => \N__27630\
        );

    \I__4387\ : Span4Mux_s1_v
    port map (
            O => \N__27630\,
            I => \N__27626\
        );

    \I__4386\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27622\
        );

    \I__4385\ : Sp12to4
    port map (
            O => \N__27626\,
            I => \N__27619\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__27625\,
            I => \N__27616\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__27622\,
            I => \N__27613\
        );

    \I__4382\ : Span12Mux_h
    port map (
            O => \N__27619\,
            I => \N__27610\
        );

    \I__4381\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27607\
        );

    \I__4380\ : Span4Mux_h
    port map (
            O => \N__27613\,
            I => \N__27604\
        );

    \I__4379\ : Odrv12
    port map (
            O => \N__27610\,
            I => \IAC_OSR0\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__27607\,
            I => \IAC_OSR0\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__27604\,
            I => \IAC_OSR0\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__27597\,
            I => \n12367_cascade_\
        );

    \I__4375\ : CascadeMux
    port map (
            O => \N__27594\,
            I => \n16563_cascade_\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__27591\,
            I => \N__27587\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__27590\,
            I => \N__27583\
        );

    \I__4372\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27580\
        );

    \I__4371\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27577\
        );

    \I__4370\ : InMux
    port map (
            O => \N__27583\,
            I => \N__27574\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__27580\,
            I => \N__27571\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__27577\,
            I => \N__27568\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27565\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__27571\,
            I => cmd_rdadctmp_27
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__27568\,
            I => cmd_rdadctmp_27
        );

    \I__4364\ : Odrv4
    port map (
            O => \N__27565\,
            I => cmd_rdadctmp_27
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__27558\,
            I => \N__27555\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27555\,
            I => \N__27552\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__27552\,
            I => \N__27547\
        );

    \I__4360\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27544\
        );

    \I__4359\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27541\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__27547\,
            I => cmd_rdadctmp_28
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27544\,
            I => cmd_rdadctmp_28
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__27541\,
            I => cmd_rdadctmp_28
        );

    \I__4355\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27531\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27531\,
            I => \N__27528\
        );

    \I__4353\ : Span4Mux_v
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__4352\ : Span4Mux_h
    port map (
            O => \N__27525\,
            I => \N__27522\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__27522\,
            I => n19_adj_1527
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__27519\,
            I => \n22279_cascade_\
        );

    \I__4349\ : InMux
    port map (
            O => \N__27516\,
            I => \N__27513\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__27513\,
            I => n17_adj_1526
        );

    \I__4347\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27507\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__27507\,
            I => \N__27504\
        );

    \I__4345\ : Odrv12
    port map (
            O => \N__27504\,
            I => n23_adj_1529
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__27501\,
            I => \n22363_cascade_\
        );

    \I__4343\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27495\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27492\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__27492\,
            I => n21285
        );

    \I__4340\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__27486\,
            I => n22282
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__27483\,
            I => \n22366_cascade_\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27476\
        );

    \I__4336\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27472\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27469\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27466\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__27472\,
            I => buf_dds1_15
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__27469\,
            I => buf_dds1_15
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__27466\,
            I => buf_dds1_15
        );

    \I__4330\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27456\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__27456\,
            I => n16_adj_1525
        );

    \I__4328\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27450\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__27450\,
            I => \N__27445\
        );

    \I__4326\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27442\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__27448\,
            I => \N__27435\
        );

    \I__4324\ : Span4Mux_v
    port map (
            O => \N__27445\,
            I => \N__27425\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27425\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27422\
        );

    \I__4321\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27419\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27416\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27413\
        );

    \I__4318\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27410\
        );

    \I__4317\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27405\
        );

    \I__4316\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27405\
        );

    \I__4315\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27398\
        );

    \I__4314\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27398\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27398\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__27425\,
            I => \N__27395\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__27422\,
            I => \N__27392\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__27419\,
            I => adc_state_1_adj_1417
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__27416\,
            I => adc_state_1_adj_1417
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27413\,
            I => adc_state_1_adj_1417
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__27410\,
            I => adc_state_1_adj_1417
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__27405\,
            I => adc_state_1_adj_1417
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__27398\,
            I => adc_state_1_adj_1417
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__27395\,
            I => adc_state_1_adj_1417
        );

    \I__4303\ : Odrv12
    port map (
            O => \N__27392\,
            I => adc_state_1_adj_1417
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__27375\,
            I => \N__27370\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__27374\,
            I => \N__27367\
        );

    \I__4300\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27364\
        );

    \I__4299\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27361\
        );

    \I__4298\ : InMux
    port map (
            O => \N__27367\,
            I => \N__27358\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__27364\,
            I => \N__27355\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__27361\,
            I => cmd_rdadctmp_24
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__27358\,
            I => cmd_rdadctmp_24
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__27355\,
            I => cmd_rdadctmp_24
        );

    \I__4293\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27340\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27337\
        );

    \I__4290\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27334\
        );

    \I__4289\ : Span12Mux_v
    port map (
            O => \N__27340\,
            I => \N__27331\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27328\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__27334\,
            I => buf_adcdata_iac_16
        );

    \I__4286\ : Odrv12
    port map (
            O => \N__27331\,
            I => buf_adcdata_iac_16
        );

    \I__4285\ : Odrv4
    port map (
            O => \N__27328\,
            I => buf_adcdata_iac_16
        );

    \I__4284\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27317\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__27320\,
            I => \N__27314\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__27317\,
            I => \N__27310\
        );

    \I__4281\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27305\
        );

    \I__4280\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27305\
        );

    \I__4279\ : Odrv12
    port map (
            O => \N__27310\,
            I => cmd_rdadctmp_26
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__27305\,
            I => cmd_rdadctmp_26
        );

    \I__4277\ : InMux
    port map (
            O => \N__27300\,
            I => \N__27291\
        );

    \I__4276\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27284\
        );

    \I__4275\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27284\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27284\
        );

    \I__4273\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27281\
        );

    \I__4272\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27276\
        );

    \I__4271\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27276\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__27291\,
            I => \N__27273\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__27284\,
            I => \N__27268\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__27281\,
            I => \N__27268\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__27276\,
            I => \N__27265\
        );

    \I__4266\ : Span4Mux_h
    port map (
            O => \N__27273\,
            I => \N__27259\
        );

    \I__4265\ : Span4Mux_v
    port map (
            O => \N__27268\,
            I => \N__27259\
        );

    \I__4264\ : Span4Mux_h
    port map (
            O => \N__27265\,
            I => \N__27256\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27253\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__27259\,
            I => n12395
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__27256\,
            I => n12395
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27253\,
            I => n12395
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__27246\,
            I => \N__27243\
        );

    \I__4258\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__27240\,
            I => \CLK_DDS.tmp_buf_11\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__4255\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__27231\,
            I => \CLK_DDS.tmp_buf_12\
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__27228\,
            I => \N__27224\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__27227\,
            I => \N__27221\
        );

    \I__4251\ : InMux
    port map (
            O => \N__27224\,
            I => \N__27218\
        );

    \I__4250\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27215\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__27218\,
            I => tmp_buf_15_adj_1455
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27215\,
            I => tmp_buf_15_adj_1455
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4246\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__27204\,
            I => \CLK_DDS.tmp_buf_7\
        );

    \I__4244\ : InMux
    port map (
            O => \N__27201\,
            I => \N__27196\
        );

    \I__4243\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27193\
        );

    \I__4242\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27190\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__27196\,
            I => \N__27187\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__27193\,
            I => buf_dds1_8
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__27190\,
            I => buf_dds1_8
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__27187\,
            I => buf_dds1_8
        );

    \I__4237\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27177\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__27177\,
            I => \N__27172\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27169\
        );

    \I__4234\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27166\
        );

    \I__4233\ : Span4Mux_h
    port map (
            O => \N__27172\,
            I => \N__27163\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__27169\,
            I => buf_dds1_13
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__27166\,
            I => buf_dds1_13
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__27163\,
            I => buf_dds1_13
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__27156\,
            I => \n11347_cascade_\
        );

    \I__4228\ : CEMux
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__27150\,
            I => n11919
        );

    \I__4226\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__27144\,
            I => buf_control_7
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__4223\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27135\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__27135\,
            I => \CLK_DDS.tmp_buf_10\
        );

    \I__4221\ : IoInMux
    port map (
            O => \N__27132\,
            I => \N__27129\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__4219\ : IoSpan4Mux
    port map (
            O => \N__27126\,
            I => \N__27123\
        );

    \I__4218\ : IoSpan4Mux
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__4217\ : Sp12to4
    port map (
            O => \N__27120\,
            I => \N__27116\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__27119\,
            I => \N__27113\
        );

    \I__4215\ : Span12Mux_s7_v
    port map (
            O => \N__27116\,
            I => \N__27110\
        );

    \I__4214\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27107\
        );

    \I__4213\ : Odrv12
    port map (
            O => \N__27110\,
            I => \DDS_SCK1\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__27107\,
            I => \DDS_SCK1\
        );

    \I__4211\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27098\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__27101\,
            I => \N__27095\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27092\
        );

    \I__4208\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27089\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__27092\,
            I => buf_adcdata_vdc_18
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__27089\,
            I => buf_adcdata_vdc_18
        );

    \I__4205\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27081\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__27081\,
            I => \N__27077\
        );

    \I__4203\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27073\
        );

    \I__4202\ : Span12Mux_h
    port map (
            O => \N__27077\,
            I => \N__27070\
        );

    \I__4201\ : InMux
    port map (
            O => \N__27076\,
            I => \N__27067\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__27073\,
            I => buf_adcdata_vac_18
        );

    \I__4199\ : Odrv12
    port map (
            O => \N__27070\,
            I => buf_adcdata_vac_18
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__27067\,
            I => buf_adcdata_vac_18
        );

    \I__4197\ : InMux
    port map (
            O => \N__27060\,
            I => \N__27057\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__27057\,
            I => \N__27054\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__27054\,
            I => \N__27051\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__27051\,
            I => \N__27048\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__27048\,
            I => n21081
        );

    \I__4192\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27041\
        );

    \I__4191\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27038\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__27041\,
            I => cmd_rdadctmp_6
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__27038\,
            I => cmd_rdadctmp_6
        );

    \I__4188\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27030\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__27027\
        );

    \I__4186\ : Span4Mux_v
    port map (
            O => \N__27027\,
            I => \N__27023\
        );

    \I__4185\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27020\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__27023\,
            I => cmd_rdadctmp_4
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__27020\,
            I => cmd_rdadctmp_4
        );

    \I__4182\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27009\
        );

    \I__4181\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27009\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__27009\,
            I => cmd_rdadctmp_5
        );

    \I__4179\ : InMux
    port map (
            O => \N__27006\,
            I => \N__27003\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__27000\
        );

    \I__4177\ : Span12Mux_h
    port map (
            O => \N__27000\,
            I => \N__26997\
        );

    \I__4176\ : Span12Mux_v
    port map (
            O => \N__26997\,
            I => \N__26994\
        );

    \I__4175\ : Odrv12
    port map (
            O => \N__26994\,
            I => \THERMOSTAT\
        );

    \I__4174\ : InMux
    port map (
            O => \N__26991\,
            I => \N__26988\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__26988\,
            I => \N__26985\
        );

    \I__4172\ : Span4Mux_h
    port map (
            O => \N__26985\,
            I => \N__26982\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__26982\,
            I => \N__26979\
        );

    \I__4170\ : Span4Mux_h
    port map (
            O => \N__26979\,
            I => \N__26976\
        );

    \I__4169\ : Odrv4
    port map (
            O => \N__26976\,
            I => buf_data_iac_0
        );

    \I__4168\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26970\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26970\,
            I => \N__26967\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__26967\,
            I => \N__26963\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__26966\,
            I => \N__26960\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__26963\,
            I => \N__26956\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26953\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26950\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__26956\,
            I => \N__26947\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__26953\,
            I => buf_adcdata_iac_0
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26950\,
            I => buf_adcdata_iac_0
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__26947\,
            I => buf_adcdata_iac_0
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26934\,
            I => \N__26931\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__26931\,
            I => \N__26927\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__26930\,
            I => \N__26924\
        );

    \I__4152\ : Span4Mux_v
    port map (
            O => \N__26927\,
            I => \N__26920\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26917\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26914\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__26920\,
            I => cmd_rdadctmp_8_adj_1442
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26917\,
            I => cmd_rdadctmp_8_adj_1442
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__26914\,
            I => cmd_rdadctmp_8_adj_1442
        );

    \I__4146\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26901\
        );

    \I__4144\ : Span4Mux_v
    port map (
            O => \N__26901\,
            I => \N__26898\
        );

    \I__4143\ : Span4Mux_h
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__26895\,
            I => \N__26890\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26885\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26885\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__26890\,
            I => buf_adcdata_vac_0
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26885\,
            I => buf_adcdata_vac_0
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__26880\,
            I => \N__26876\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26871\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26876\,
            I => \N__26871\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26871\,
            I => \N__26868\
        );

    \I__4133\ : Span4Mux_h
    port map (
            O => \N__26868\,
            I => \N__26864\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26867\,
            I => \N__26861\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__26864\,
            I => cmd_rdadctmp_8
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26861\,
            I => cmd_rdadctmp_8
        );

    \I__4129\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__26853\,
            I => \N__26826\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26821\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26821\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26816\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26849\,
            I => \N__26798\
        );

    \I__4123\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26798\
        );

    \I__4122\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26798\
        );

    \I__4121\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26798\
        );

    \I__4120\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26798\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26798\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26798\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26798\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26789\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26789\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26789\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26789\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__26837\,
            I => \N__26786\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26836\,
            I => \N__26779\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26773\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26773\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26768\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26768\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26757\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26754\
        );

    \I__4104\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26751\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__26826\,
            I => \N__26744\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26821\,
            I => \N__26744\
        );

    \I__4101\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26739\
        );

    \I__4100\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26739\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__26816\,
            I => \N__26736\
        );

    \I__4098\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26732\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__26798\,
            I => \N__26727\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__26789\,
            I => \N__26727\
        );

    \I__4095\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26717\
        );

    \I__4094\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26717\
        );

    \I__4093\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26717\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26714\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26711\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__26779\,
            I => \N__26708\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26705\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26773\,
            I => \N__26700\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26768\,
            I => \N__26700\
        );

    \I__4086\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26693\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26693\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26693\
        );

    \I__4083\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26686\
        );

    \I__4082\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26686\
        );

    \I__4081\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26686\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26681\
        );

    \I__4079\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26681\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__26757\,
            I => \N__26674\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26674\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26674\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26669\
        );

    \I__4074\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26669\
        );

    \I__4073\ : Span4Mux_v
    port map (
            O => \N__26744\,
            I => \N__26662\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__26739\,
            I => \N__26662\
        );

    \I__4071\ : Span4Mux_h
    port map (
            O => \N__26736\,
            I => \N__26662\
        );

    \I__4070\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26659\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26656\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__26727\,
            I => \N__26653\
        );

    \I__4067\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26648\
        );

    \I__4066\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26648\
        );

    \I__4065\ : InMux
    port map (
            O => \N__26724\,
            I => \N__26645\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26642\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__26714\,
            I => \N__26637\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__26711\,
            I => \N__26637\
        );

    \I__4061\ : Span4Mux_v
    port map (
            O => \N__26708\,
            I => \N__26622\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__26705\,
            I => \N__26622\
        );

    \I__4059\ : Span4Mux_v
    port map (
            O => \N__26700\,
            I => \N__26622\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__26693\,
            I => \N__26622\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__26686\,
            I => \N__26622\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__26681\,
            I => \N__26622\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__26674\,
            I => \N__26622\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__26669\,
            I => \N__26615\
        );

    \I__4053\ : Span4Mux_h
    port map (
            O => \N__26662\,
            I => \N__26615\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__26659\,
            I => \N__26615\
        );

    \I__4051\ : Odrv12
    port map (
            O => \N__26656\,
            I => adc_state_2_adj_1481
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__26653\,
            I => adc_state_2_adj_1481
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__26648\,
            I => adc_state_2_adj_1481
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__26645\,
            I => adc_state_2_adj_1481
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__26642\,
            I => adc_state_2_adj_1481
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__26637\,
            I => adc_state_2_adj_1481
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__26622\,
            I => adc_state_2_adj_1481
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__26615\,
            I => adc_state_2_adj_1481
        );

    \I__4043\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26586\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__26597\,
            I => \N__26581\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26577\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26572\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26572\
        );

    \I__4038\ : InMux
    port map (
            O => \N__26593\,
            I => \N__26569\
        );

    \I__4037\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26566\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__26591\,
            I => \N__26562\
        );

    \I__4035\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26554\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26554\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__26586\,
            I => \N__26551\
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__26585\,
            I => \N__26548\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__26584\,
            I => \N__26545\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26536\
        );

    \I__4029\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26536\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__26577\,
            I => \N__26530\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__26572\,
            I => \N__26527\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26569\,
            I => \N__26522\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__26566\,
            I => \N__26522\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26513\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26513\
        );

    \I__4022\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26513\
        );

    \I__4021\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26513\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26559\,
            I => \N__26510\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__26554\,
            I => \N__26505\
        );

    \I__4018\ : Span4Mux_h
    port map (
            O => \N__26551\,
            I => \N__26505\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26498\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26545\,
            I => \N__26498\
        );

    \I__4015\ : InMux
    port map (
            O => \N__26544\,
            I => \N__26498\
        );

    \I__4014\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26493\
        );

    \I__4013\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26493\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26490\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__26536\,
            I => \N__26487\
        );

    \I__4010\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26482\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26534\,
            I => \N__26482\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26479\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__26530\,
            I => \N__26470\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__26527\,
            I => \N__26470\
        );

    \I__4005\ : Span4Mux_v
    port map (
            O => \N__26522\,
            I => \N__26470\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__26513\,
            I => \N__26470\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26510\,
            I => \N__26463\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__26505\,
            I => \N__26463\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__26498\,
            I => \N__26463\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26493\,
            I => \RTD.adc_state_1\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__26490\,
            I => \RTD.adc_state_1\
        );

    \I__3998\ : Odrv4
    port map (
            O => \N__26487\,
            I => \RTD.adc_state_1\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__26482\,
            I => \RTD.adc_state_1\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__26479\,
            I => \RTD.adc_state_1\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__26470\,
            I => \RTD.adc_state_1\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__26463\,
            I => \RTD.adc_state_1\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__26448\,
            I => \N__26444\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__26447\,
            I => \N__26438\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26428\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__26443\,
            I => \N__26422\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__26442\,
            I => \N__26416\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__26441\,
            I => \N__26412\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26409\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26404\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26404\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26401\
        );

    \I__3983\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26392\
        );

    \I__3982\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26392\
        );

    \I__3981\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26392\
        );

    \I__3980\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26392\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__26428\,
            I => \N__26386\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__26427\,
            I => \N__26382\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26373\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26373\
        );

    \I__3975\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26373\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__26421\,
            I => \N__26370\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26363\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26363\
        );

    \I__3971\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26363\
        );

    \I__3970\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26360\
        );

    \I__3969\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26357\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__26409\,
            I => \N__26350\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26350\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__26401\,
            I => \N__26350\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__26392\,
            I => \N__26347\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__26391\,
            I => \N__26344\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26339\
        );

    \I__3962\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26339\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__26386\,
            I => \N__26336\
        );

    \I__3960\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26333\
        );

    \I__3959\ : InMux
    port map (
            O => \N__26382\,
            I => \N__26328\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26328\
        );

    \I__3957\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26325\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__26373\,
            I => \N__26322\
        );

    \I__3955\ : InMux
    port map (
            O => \N__26370\,
            I => \N__26319\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__26363\,
            I => \N__26316\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26311\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26357\,
            I => \N__26311\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__26350\,
            I => \N__26306\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__26347\,
            I => \N__26306\
        );

    \I__3949\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26303\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26298\
        );

    \I__3947\ : Sp12to4
    port map (
            O => \N__26336\,
            I => \N__26298\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__26333\,
            I => \RTD.adc_state_3\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__26328\,
            I => \RTD.adc_state_3\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__26325\,
            I => \RTD.adc_state_3\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__26322\,
            I => \RTD.adc_state_3\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__26319\,
            I => \RTD.adc_state_3\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__26316\,
            I => \RTD.adc_state_3\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__26311\,
            I => \RTD.adc_state_3\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__26306\,
            I => \RTD.adc_state_3\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__26303\,
            I => \RTD.adc_state_3\
        );

    \I__3937\ : Odrv12
    port map (
            O => \N__26298\,
            I => \RTD.adc_state_3\
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__26277\,
            I => \N__26274\
        );

    \I__3935\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26254\
        );

    \I__3934\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26248\
        );

    \I__3933\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26245\
        );

    \I__3932\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26242\
        );

    \I__3931\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26235\
        );

    \I__3930\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26235\
        );

    \I__3929\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26235\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26225\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26225\
        );

    \I__3926\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26225\
        );

    \I__3925\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26222\
        );

    \I__3924\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26219\
        );

    \I__3923\ : InMux
    port map (
            O => \N__26262\,
            I => \N__26214\
        );

    \I__3922\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26214\
        );

    \I__3921\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26207\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26207\
        );

    \I__3919\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26207\
        );

    \I__3918\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26196\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26193\
        );

    \I__3916\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26190\
        );

    \I__3915\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26184\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26251\,
            I => \N__26181\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__26248\,
            I => \N__26174\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__26245\,
            I => \N__26174\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__26242\,
            I => \N__26174\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__26235\,
            I => \N__26171\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26164\
        );

    \I__3908\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26164\
        );

    \I__3907\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26164\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26161\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26158\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__26219\,
            I => \N__26151\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__26214\,
            I => \N__26151\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__26207\,
            I => \N__26151\
        );

    \I__3901\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26134\
        );

    \I__3900\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26134\
        );

    \I__3899\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26134\
        );

    \I__3898\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26134\
        );

    \I__3897\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26134\
        );

    \I__3896\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26134\
        );

    \I__3895\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26134\
        );

    \I__3894\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26134\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__26196\,
            I => \N__26131\
        );

    \I__3892\ : Span4Mux_h
    port map (
            O => \N__26193\,
            I => \N__26126\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__26190\,
            I => \N__26126\
        );

    \I__3890\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26119\
        );

    \I__3889\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26119\
        );

    \I__3888\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26119\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__26184\,
            I => \N__26112\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26181\,
            I => \N__26112\
        );

    \I__3885\ : Span4Mux_v
    port map (
            O => \N__26174\,
            I => \N__26112\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__26171\,
            I => \N__26101\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__26164\,
            I => \N__26101\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__26161\,
            I => \N__26101\
        );

    \I__3881\ : Span4Mux_h
    port map (
            O => \N__26158\,
            I => \N__26101\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__26151\,
            I => \N__26101\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__26134\,
            I => \RTD.adc_state_0\
        );

    \I__3878\ : Odrv12
    port map (
            O => \N__26131\,
            I => \RTD.adc_state_0\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__26126\,
            I => \RTD.adc_state_0\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__26119\,
            I => \RTD.adc_state_0\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__26112\,
            I => \RTD.adc_state_0\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__26101\,
            I => \RTD.adc_state_0\
        );

    \I__3873\ : SRMux
    port map (
            O => \N__26088\,
            I => \N__26085\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__26085\,
            I => \N__26082\
        );

    \I__3871\ : Sp12to4
    port map (
            O => \N__26082\,
            I => \N__26079\
        );

    \I__3870\ : Odrv12
    port map (
            O => \N__26079\,
            I => \RTD.n15065\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__26076\,
            I => \n13087_cascade_\
        );

    \I__3868\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26070\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26067\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__26067\,
            I => \N__26063\
        );

    \I__3865\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26060\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__26063\,
            I => cmd_rdadcbuf_26
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__26060\,
            I => cmd_rdadcbuf_26
        );

    \I__3862\ : InMux
    port map (
            O => \N__26055\,
            I => \N__26052\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__26052\,
            I => \N__26048\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__26051\,
            I => \N__26044\
        );

    \I__3859\ : Span4Mux_h
    port map (
            O => \N__26048\,
            I => \N__26041\
        );

    \I__3858\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26038\
        );

    \I__3857\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26035\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__26041\,
            I => cmd_rdadctmp_22_adj_1457
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__26038\,
            I => cmd_rdadctmp_22_adj_1457
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__26035\,
            I => cmd_rdadctmp_22_adj_1457
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__26028\,
            I => \N__26025\
        );

    \I__3852\ : InMux
    port map (
            O => \N__26025\,
            I => \N__26021\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__26024\,
            I => \N__26018\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__26021\,
            I => \N__26015\
        );

    \I__3849\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26012\
        );

    \I__3848\ : Span4Mux_h
    port map (
            O => \N__26015\,
            I => \N__26009\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__26012\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__26009\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__3845\ : CEMux
    port map (
            O => \N__26004\,
            I => \N__26001\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__26001\,
            I => \N__25998\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__25998\,
            I => \N__25995\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__25995\,
            I => \ADC_VDC.n12899\
        );

    \I__3841\ : SRMux
    port map (
            O => \N__25992\,
            I => \N__25989\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__25989\,
            I => \N__25986\
        );

    \I__3839\ : Odrv12
    port map (
            O => \N__25986\,
            I => \ADC_VDC.n20656\
        );

    \I__3838\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25980\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__25980\,
            I => \comm_spi.n22860\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__25977\,
            I => \comm_spi.n22860_cascade_\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25971\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__25971\,
            I => \N__25968\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__25968\,
            I => \comm_spi.n14597\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25961\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__25964\,
            I => \N__25958\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__25961\,
            I => \N__25955\
        );

    \I__3829\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25952\
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__25955\,
            I => buf_adcdata_vdc_0
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__25952\,
            I => buf_adcdata_vdc_0
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__25947\,
            I => \n19_adj_1484_cascade_\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__25944\,
            I => \n22_adj_1483_cascade_\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__25941\,
            I => \N__25937\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__25940\,
            I => \N__25933\
        );

    \I__3822\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25930\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__25936\,
            I => \N__25926\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25923\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25930\,
            I => \N__25919\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25914\
        );

    \I__3817\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25914\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25923\,
            I => \N__25911\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__25922\,
            I => \N__25908\
        );

    \I__3814\ : Span4Mux_v
    port map (
            O => \N__25919\,
            I => \N__25905\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__25914\,
            I => \N__25902\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__25911\,
            I => \N__25899\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25896\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__25905\,
            I => \N__25891\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__25902\,
            I => \N__25891\
        );

    \I__3808\ : Sp12to4
    port map (
            O => \N__25899\,
            I => \N__25884\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__25896\,
            I => \N__25884\
        );

    \I__3806\ : Sp12to4
    port map (
            O => \N__25891\,
            I => \N__25884\
        );

    \I__3805\ : Span12Mux_h
    port map (
            O => \N__25884\,
            I => \N__25881\
        );

    \I__3804\ : Odrv12
    port map (
            O => \N__25881\,
            I => \IAC_DRDY\
        );

    \I__3803\ : CEMux
    port map (
            O => \N__25878\,
            I => \N__25874\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25871\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__25874\,
            I => \N__25868\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25871\,
            I => \N__25865\
        );

    \I__3799\ : Span4Mux_h
    port map (
            O => \N__25868\,
            I => \N__25862\
        );

    \I__3798\ : Span4Mux_h
    port map (
            O => \N__25865\,
            I => \N__25859\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__25862\,
            I => \ADC_IAC.n12473\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__25859\,
            I => \ADC_IAC.n12473\
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__25854\,
            I => \ADC_VDC.n11676_cascade_\
        );

    \I__3794\ : IoInMux
    port map (
            O => \N__25851\,
            I => \N__25848\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25848\,
            I => \N__25845\
        );

    \I__3792\ : IoSpan4Mux
    port map (
            O => \N__25845\,
            I => \N__25842\
        );

    \I__3791\ : Span4Mux_s3_h
    port map (
            O => \N__25842\,
            I => \N__25839\
        );

    \I__3790\ : Span4Mux_h
    port map (
            O => \N__25839\,
            I => \N__25836\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__25836\,
            I => \N__25832\
        );

    \I__3788\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25829\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__25832\,
            I => \VDC_SCLK\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25829\,
            I => \VDC_SCLK\
        );

    \I__3785\ : SRMux
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25818\
        );

    \I__3783\ : Span4Mux_h
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__25815\,
            I => \comm_spi.iclk_N_763\
        );

    \I__3781\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__25809\,
            I => \N__25806\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__25803\,
            I => \N__25799\
        );

    \I__3777\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25796\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__25799\,
            I => cmd_rdadcbuf_33
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__25796\,
            I => cmd_rdadcbuf_33
        );

    \I__3774\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25788\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__25788\,
            I => \N__25785\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__25785\,
            I => \N__25781\
        );

    \I__3771\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25778\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__25781\,
            I => cmd_rdadcbuf_11
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25778\,
            I => cmd_rdadcbuf_11
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__25773\,
            I => \N__25770\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25767\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__25767\,
            I => \N__25764\
        );

    \I__3765\ : Span4Mux_v
    port map (
            O => \N__25764\,
            I => \N__25760\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25757\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__25760\,
            I => cmd_rdadcbuf_21
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__25757\,
            I => cmd_rdadcbuf_21
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__25752\,
            I => \N__25737\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25751\,
            I => \N__25720\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25750\,
            I => \N__25720\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25720\
        );

    \I__3757\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25720\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25720\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25720\
        );

    \I__3754\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25720\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25709\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25709\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25709\
        );

    \I__3750\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25709\
        );

    \I__3749\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25709\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25702\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25702\
        );

    \I__3746\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25702\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25720\,
            I => \N__25698\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25695\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__25702\,
            I => \N__25692\
        );

    \I__3742\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25689\
        );

    \I__3741\ : Span4Mux_v
    port map (
            O => \N__25698\,
            I => \N__25679\
        );

    \I__3740\ : Span4Mux_h
    port map (
            O => \N__25695\,
            I => \N__25676\
        );

    \I__3739\ : Span4Mux_h
    port map (
            O => \N__25692\,
            I => \N__25673\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25689\,
            I => \N__25670\
        );

    \I__3737\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25665\
        );

    \I__3736\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25665\
        );

    \I__3735\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25660\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25660\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25653\
        );

    \I__3732\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25653\
        );

    \I__3731\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25653\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__25679\,
            I => n13087
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__25676\,
            I => n13087
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__25673\,
            I => n13087
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__25670\,
            I => n13087
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__25665\,
            I => n13087
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__25660\,
            I => n13087
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__25653\,
            I => n13087
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__25638\,
            I => \ADC_IAC.n20960_cascade_\
        );

    \I__3722\ : CEMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__3720\ : Span4Mux_h
    port map (
            O => \N__25629\,
            I => \N__25626\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__25626\,
            I => \ADC_IAC.n20961\
        );

    \I__3718\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25619\
        );

    \I__3717\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25616\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__25619\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__25616\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__3714\ : InMux
    port map (
            O => \N__25611\,
            I => \N__25607\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25604\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__25607\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__25604\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__25599\,
            I => \N__25595\
        );

    \I__3709\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25592\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__25592\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25589\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25580\
        );

    \I__3704\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25577\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__25580\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__25577\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25568\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25565\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__25568\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__25565\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__3697\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25556\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25553\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__25556\,
            I => \N__25550\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__25553\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__25550\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__25545\,
            I => \ADC_IAC.n21295_cascade_\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25539\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__25539\,
            I => \ADC_IAC.n21294\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25532\
        );

    \I__3688\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25529\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__25532\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__25529\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__3685\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25520\
        );

    \I__3684\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25517\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__25520\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__25517\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__25512\,
            I => \N__25508\
        );

    \I__3680\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25505\
        );

    \I__3679\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25502\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__25505\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__25502\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__3676\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25493\
        );

    \I__3675\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25490\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__25493\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__25490\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25481\
        );

    \I__3671\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25478\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__25481\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25478\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__3668\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25469\
        );

    \I__3667\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25466\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__25469\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__25466\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__25461\,
            I => \ADC_VAC.n21029_cascade_\
        );

    \I__3663\ : InMux
    port map (
            O => \N__25458\,
            I => \N__25454\
        );

    \I__3662\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25451\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__25454\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__25451\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__3659\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__25440\,
            I => \ADC_VAC.n21043\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__25437\,
            I => \N__25433\
        );

    \I__3655\ : InMux
    port map (
            O => \N__25436\,
            I => \N__25430\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25427\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25430\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__25427\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__3651\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25418\
        );

    \I__3650\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25415\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__25418\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25415\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__3647\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__25407\,
            I => \ADC_IAC.n16\
        );

    \I__3645\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25399\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25396\
        );

    \I__3643\ : CascadeMux
    port map (
            O => \N__25402\,
            I => \N__25393\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__25399\,
            I => \N__25386\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__25396\,
            I => \N__25386\
        );

    \I__3640\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25383\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25380\
        );

    \I__3638\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25377\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__25386\,
            I => \N__25374\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25383\,
            I => acadc_trig
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__25380\,
            I => acadc_trig
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__25377\,
            I => acadc_trig
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__25374\,
            I => acadc_trig
        );

    \I__3632\ : IoInMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__3630\ : Span4Mux_s1_h
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__3629\ : Sp12to4
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__3628\ : Span12Mux_s11_v
    port map (
            O => \N__25353\,
            I => \N__25348\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25343\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25351\,
            I => \N__25343\
        );

    \I__3625\ : Odrv12
    port map (
            O => \N__25348\,
            I => \VAC_FLT1\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__25343\,
            I => \VAC_FLT1\
        );

    \I__3623\ : InMux
    port map (
            O => \N__25338\,
            I => \bfn_9_16_0_\
        );

    \I__3622\ : InMux
    port map (
            O => \N__25335\,
            I => \ADC_VAC.n19656\
        );

    \I__3621\ : InMux
    port map (
            O => \N__25332\,
            I => \ADC_VAC.n19657\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25329\,
            I => \ADC_VAC.n19658\
        );

    \I__3619\ : InMux
    port map (
            O => \N__25326\,
            I => \ADC_VAC.n19659\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__25323\,
            I => \N__25320\
        );

    \I__3617\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25317\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25313\
        );

    \I__3615\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25310\
        );

    \I__3614\ : Sp12to4
    port map (
            O => \N__25313\,
            I => \N__25307\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__25310\,
            I => \N__25302\
        );

    \I__3612\ : Span12Mux_s10_v
    port map (
            O => \N__25307\,
            I => \N__25302\
        );

    \I__3611\ : Odrv12
    port map (
            O => \N__25302\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__3610\ : InMux
    port map (
            O => \N__25299\,
            I => \ADC_VAC.n19660\
        );

    \I__3609\ : InMux
    port map (
            O => \N__25296\,
            I => \ADC_VAC.n19661\
        );

    \I__3608\ : InMux
    port map (
            O => \N__25293\,
            I => \ADC_VAC.n19662\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25287\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__25287\,
            I => \N__25283\
        );

    \I__3605\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25279\
        );

    \I__3604\ : Span4Mux_v
    port map (
            O => \N__25283\,
            I => \N__25276\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__25282\,
            I => \N__25273\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__25279\,
            I => \N__25270\
        );

    \I__3601\ : Sp12to4
    port map (
            O => \N__25276\,
            I => \N__25267\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25264\
        );

    \I__3599\ : Span4Mux_v
    port map (
            O => \N__25270\,
            I => \N__25261\
        );

    \I__3598\ : Span12Mux_h
    port map (
            O => \N__25267\,
            I => \N__25258\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__25264\,
            I => buf_adcdata_vac_19
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__25261\,
            I => buf_adcdata_vac_19
        );

    \I__3595\ : Odrv12
    port map (
            O => \N__25258\,
            I => buf_adcdata_vac_19
        );

    \I__3594\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__25245\,
            I => n22435
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25236\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__25236\,
            I => \N__25232\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__25235\,
            I => \N__25229\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__25232\,
            I => \N__25226\
        );

    \I__3586\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25223\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__25226\,
            I => buf_adcdata_vdc_19
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__25223\,
            I => buf_adcdata_vdc_19
        );

    \I__3583\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25212\
        );

    \I__3582\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25212\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__25212\,
            I => \N__25209\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__25209\,
            I => cmd_rdadctmp_31
        );

    \I__3579\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25202\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__25205\,
            I => \N__25198\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__25202\,
            I => \N__25195\
        );

    \I__3576\ : InMux
    port map (
            O => \N__25201\,
            I => \N__25190\
        );

    \I__3575\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25190\
        );

    \I__3574\ : Odrv4
    port map (
            O => \N__25195\,
            I => cmd_rdadctmp_29
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__25190\,
            I => cmd_rdadctmp_29
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__25185\,
            I => \N__25180\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__25184\,
            I => \N__25177\
        );

    \I__3570\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25172\
        );

    \I__3569\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25172\
        );

    \I__3568\ : InMux
    port map (
            O => \N__25177\,
            I => \N__25169\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__25172\,
            I => cmd_rdadctmp_30
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__25169\,
            I => cmd_rdadctmp_30
        );

    \I__3565\ : InMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__25158\,
            I => \N__25154\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__25157\,
            I => \N__25151\
        );

    \I__3561\ : Sp12to4
    port map (
            O => \N__25154\,
            I => \N__25147\
        );

    \I__3560\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25144\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25150\,
            I => \N__25141\
        );

    \I__3558\ : Span12Mux_v
    port map (
            O => \N__25147\,
            I => \N__25138\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__25144\,
            I => buf_adcdata_iac_23
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__25141\,
            I => buf_adcdata_iac_23
        );

    \I__3555\ : Odrv12
    port map (
            O => \N__25138\,
            I => buf_adcdata_iac_23
        );

    \I__3554\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__25128\,
            I => \N__25123\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__25127\,
            I => \N__25120\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25117\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__25123\,
            I => \N__25114\
        );

    \I__3549\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25111\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__25117\,
            I => cmd_rdadctmp_23
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__25114\,
            I => cmd_rdadctmp_23
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__25111\,
            I => cmd_rdadctmp_23
        );

    \I__3545\ : InMux
    port map (
            O => \N__25104\,
            I => \N__25101\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__25101\,
            I => n22417
        );

    \I__3543\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25092\
        );

    \I__3541\ : Span4Mux_v
    port map (
            O => \N__25092\,
            I => \N__25087\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__25091\,
            I => \N__25084\
        );

    \I__3539\ : InMux
    port map (
            O => \N__25090\,
            I => \N__25081\
        );

    \I__3538\ : Sp12to4
    port map (
            O => \N__25087\,
            I => \N__25078\
        );

    \I__3537\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25075\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25072\
        );

    \I__3535\ : Span12Mux_h
    port map (
            O => \N__25078\,
            I => \N__25069\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__25075\,
            I => buf_adcdata_vac_20
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__25072\,
            I => buf_adcdata_vac_20
        );

    \I__3532\ : Odrv12
    port map (
            O => \N__25069\,
            I => buf_adcdata_vac_20
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__3530\ : InMux
    port map (
            O => \N__25059\,
            I => \N__25055\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__25058\,
            I => \N__25052\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__25055\,
            I => \N__25049\
        );

    \I__3527\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25046\
        );

    \I__3526\ : Odrv12
    port map (
            O => \N__25049\,
            I => buf_adcdata_vdc_20
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__25046\,
            I => buf_adcdata_vdc_20
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__3523\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25031\
        );

    \I__3522\ : InMux
    port map (
            O => \N__25037\,
            I => \N__25031\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__25036\,
            I => \N__25028\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__25025\
        );

    \I__3519\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25022\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__25025\,
            I => cmd_rdadctmp_20
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__25022\,
            I => cmd_rdadctmp_20
        );

    \I__3516\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__25014\,
            I => n21139
        );

    \I__3514\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__25008\,
            I => n22291
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__25005\,
            I => \n21138_cascade_\
        );

    \I__3511\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24999\,
            I => \N__24994\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__24998\,
            I => \N__24991\
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__24997\,
            I => \N__24988\
        );

    \I__3507\ : Span12Mux_s9_v
    port map (
            O => \N__24994\,
            I => \N__24985\
        );

    \I__3506\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24982\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24988\,
            I => \N__24979\
        );

    \I__3504\ : Span12Mux_h
    port map (
            O => \N__24985\,
            I => \N__24976\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__24982\,
            I => buf_adcdata_iac_21
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24979\,
            I => buf_adcdata_iac_21
        );

    \I__3501\ : Odrv12
    port map (
            O => \N__24976\,
            I => buf_adcdata_iac_21
        );

    \I__3500\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__24966\,
            I => \N__24962\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__24965\,
            I => \N__24959\
        );

    \I__3497\ : Span4Mux_v
    port map (
            O => \N__24962\,
            I => \N__24956\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24953\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__24956\,
            I => buf_adcdata_vdc_13
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24953\,
            I => buf_adcdata_vdc_13
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__24948\,
            I => \N__24943\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__24947\,
            I => \N__24940\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24937\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24932\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24932\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__24937\,
            I => cmd_rdadctmp_21_adj_1429
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__24932\,
            I => cmd_rdadctmp_21_adj_1429
        );

    \I__3486\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24924\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24921\
        );

    \I__3484\ : Span12Mux_v
    port map (
            O => \N__24921\,
            I => \N__24918\
        );

    \I__3483\ : Span12Mux_h
    port map (
            O => \N__24918\,
            I => \N__24913\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24917\,
            I => \N__24908\
        );

    \I__3481\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24908\
        );

    \I__3480\ : Odrv12
    port map (
            O => \N__24913\,
            I => buf_adcdata_vac_13
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__24908\,
            I => buf_adcdata_vac_13
        );

    \I__3478\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24898\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__24902\,
            I => \N__24895\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24892\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__24898\,
            I => \N__24889\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24895\,
            I => \N__24886\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24892\,
            I => cmd_rdadctmp_22_adj_1428
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__24889\,
            I => cmd_rdadctmp_22_adj_1428
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__24886\,
            I => cmd_rdadctmp_22_adj_1428
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__24879\,
            I => \N__24874\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24871\
        );

    \I__3468\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24866\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24874\,
            I => \N__24866\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__24871\,
            I => cmd_rdadctmp_20_adj_1430
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__24866\,
            I => cmd_rdadctmp_20_adj_1430
        );

    \I__3464\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24858\,
            I => \N__24855\
        );

    \I__3462\ : Span12Mux_v
    port map (
            O => \N__24855\,
            I => \N__24851\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24847\
        );

    \I__3460\ : Span12Mux_h
    port map (
            O => \N__24851\,
            I => \N__24844\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24850\,
            I => \N__24841\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24847\,
            I => buf_adcdata_vac_12
        );

    \I__3457\ : Odrv12
    port map (
            O => \N__24844\,
            I => buf_adcdata_vac_12
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__24841\,
            I => buf_adcdata_vac_12
        );

    \I__3455\ : InMux
    port map (
            O => \N__24834\,
            I => \N__24830\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24827\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__24830\,
            I => \N__24823\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__24827\,
            I => \N__24820\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24817\
        );

    \I__3450\ : Span12Mux_s11_h
    port map (
            O => \N__24823\,
            I => \N__24814\
        );

    \I__3449\ : Span4Mux_h
    port map (
            O => \N__24820\,
            I => \N__24811\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24817\,
            I => buf_adcdata_iac_7
        );

    \I__3447\ : Odrv12
    port map (
            O => \N__24814\,
            I => buf_adcdata_iac_7
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24811\,
            I => buf_adcdata_iac_7
        );

    \I__3445\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__24798\,
            I => n19_adj_1623
        );

    \I__3442\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__3439\ : Span4Mux_h
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__24783\,
            I => buf_data_iac_7
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__24780\,
            I => \n22_adj_1624_cascade_\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24767\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24767\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24775\,
            I => \N__24767\
        );

    \I__3433\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24764\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__24767\,
            I => \N__24758\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__24764\,
            I => \N__24758\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24755\
        );

    \I__3429\ : Span4Mux_v
    port map (
            O => \N__24758\,
            I => \N__24752\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__24755\,
            I => bit_cnt_0_adj_1456
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__24752\,
            I => bit_cnt_0_adj_1456
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__24747\,
            I => \N__24744\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24740\
        );

    \I__3424\ : CascadeMux
    port map (
            O => \N__24743\,
            I => \N__24737\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24740\,
            I => \N__24734\
        );

    \I__3422\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24731\
        );

    \I__3421\ : Odrv12
    port map (
            O => \N__24734\,
            I => cmd_rdadctmp_7
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__24731\,
            I => cmd_rdadctmp_7
        );

    \I__3419\ : IoInMux
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24723\,
            I => \N__24720\
        );

    \I__3417\ : IoSpan4Mux
    port map (
            O => \N__24720\,
            I => \N__24717\
        );

    \I__3416\ : Span4Mux_s3_v
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__3413\ : Span4Mux_v
    port map (
            O => \N__24708\,
            I => \N__24704\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24707\,
            I => \N__24701\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__24704\,
            I => \DDS_MOSI1\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24701\,
            I => \DDS_MOSI1\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__24696\,
            I => \N__24693\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24688\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24685\
        );

    \I__3406\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24682\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__24688\,
            I => \N__24679\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__24685\,
            I => \N__24675\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__24682\,
            I => \N__24672\
        );

    \I__3402\ : Span4Mux_v
    port map (
            O => \N__24679\,
            I => \N__24668\
        );

    \I__3401\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24665\
        );

    \I__3400\ : Span4Mux_h
    port map (
            O => \N__24675\,
            I => \N__24662\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__24672\,
            I => \N__24659\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24656\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__24668\,
            I => \N__24651\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24665\,
            I => \N__24651\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__24662\,
            I => \N__24646\
        );

    \I__3394\ : Span4Mux_h
    port map (
            O => \N__24659\,
            I => \N__24646\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__24656\,
            I => \N__24641\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__24651\,
            I => \N__24641\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__24646\,
            I => \buf_cfgRTD_3\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__24641\,
            I => \buf_cfgRTD_3\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__3388\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24630\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__24630\,
            I => \N__24626\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__24629\,
            I => \N__24623\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__24626\,
            I => \N__24620\
        );

    \I__3384\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24617\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__24620\,
            I => \buf_readRTD_11\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__24617\,
            I => \buf_readRTD_11\
        );

    \I__3381\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24609\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24605\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__24608\,
            I => \N__24602\
        );

    \I__3378\ : Span4Mux_v
    port map (
            O => \N__24605\,
            I => \N__24599\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24596\
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__24599\,
            I => buf_adcdata_vdc_12
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__24596\,
            I => buf_adcdata_vdc_12
        );

    \I__3374\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24588\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__24588\,
            I => n19_adj_1511
        );

    \I__3372\ : InMux
    port map (
            O => \N__24585\,
            I => \N__24581\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24578\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__24581\,
            I => cmd_rdadcbuf_32
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__24578\,
            I => cmd_rdadcbuf_32
        );

    \I__3368\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24570\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24566\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__24569\,
            I => \N__24563\
        );

    \I__3365\ : Span4Mux_v
    port map (
            O => \N__24566\,
            I => \N__24560\
        );

    \I__3364\ : InMux
    port map (
            O => \N__24563\,
            I => \N__24557\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__24560\,
            I => buf_adcdata_vdc_21
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__24557\,
            I => buf_adcdata_vdc_21
        );

    \I__3361\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24548\
        );

    \I__3360\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24545\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__24548\,
            I => cmd_rdadcbuf_31
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24545\,
            I => cmd_rdadcbuf_31
        );

    \I__3357\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24536\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24533\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24536\,
            I => cmd_rdadcbuf_30
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__24533\,
            I => cmd_rdadcbuf_30
        );

    \I__3353\ : InMux
    port map (
            O => \N__24528\,
            I => \N__24524\
        );

    \I__3352\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24521\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__24524\,
            I => cmd_rdadcbuf_29
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__24521\,
            I => cmd_rdadcbuf_29
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__3348\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24510\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__24510\,
            I => \N__24506\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__24509\,
            I => \N__24502\
        );

    \I__3345\ : Span4Mux_v
    port map (
            O => \N__24506\,
            I => \N__24499\
        );

    \I__3344\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24494\
        );

    \I__3343\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24494\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__24499\,
            I => cmd_rdadctmp_23_adj_1427
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__24494\,
            I => cmd_rdadctmp_23_adj_1427
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__24489\,
            I => \N__24486\
        );

    \I__3339\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24481\
        );

    \I__3338\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24478\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__24484\,
            I => \N__24475\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24472\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24469\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24466\
        );

    \I__3333\ : Span4Mux_v
    port map (
            O => \N__24472\,
            I => \N__24463\
        );

    \I__3332\ : Span4Mux_h
    port map (
            O => \N__24469\,
            I => \N__24460\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__24466\,
            I => cmd_rdadctmp_26_adj_1424
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__24463\,
            I => cmd_rdadctmp_26_adj_1424
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__24460\,
            I => cmd_rdadctmp_26_adj_1424
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__24453\,
            I => \N__24449\
        );

    \I__3327\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24446\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24443\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24446\,
            I => buf_adcdata_vdc_17
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__24443\,
            I => buf_adcdata_vdc_17
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__24438\,
            I => \N__24435\
        );

    \I__3322\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24432\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__24432\,
            I => \N__24429\
        );

    \I__3320\ : Span4Mux_h
    port map (
            O => \N__24429\,
            I => \N__24426\
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__24426\,
            I => n22441
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__24423\,
            I => \N__24420\
        );

    \I__3317\ : InMux
    port map (
            O => \N__24420\,
            I => \N__24417\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__24417\,
            I => \N__24413\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__24416\,
            I => \N__24409\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__24413\,
            I => \N__24406\
        );

    \I__3313\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24403\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24400\
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__24406\,
            I => cmd_rdadctmp_25_adj_1425
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__24403\,
            I => cmd_rdadctmp_25_adj_1425
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__24400\,
            I => cmd_rdadctmp_25_adj_1425
        );

    \I__3308\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__3306\ : Span4Mux_v
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__3304\ : Span4Mux_h
    port map (
            O => \N__24381\,
            I => \N__24376\
        );

    \I__3303\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24371\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24371\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__24376\,
            I => buf_adcdata_vac_17
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24371\,
            I => buf_adcdata_vac_17
        );

    \I__3299\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24362\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24359\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24362\,
            I => cmd_rdadcbuf_24
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__24359\,
            I => cmd_rdadcbuf_24
        );

    \I__3295\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24351\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__24351\,
            I => \N__24347\
        );

    \I__3293\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24344\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__24347\,
            I => cmd_rdadcbuf_17
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__24344\,
            I => cmd_rdadcbuf_17
        );

    \I__3290\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24336\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24336\,
            I => \N__24333\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__24333\,
            I => \N__24329\
        );

    \I__3287\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24326\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__24329\,
            I => buf_adcdata_vdc_6
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__24326\,
            I => buf_adcdata_vdc_6
        );

    \I__3284\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24317\
        );

    \I__3283\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24314\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__24317\,
            I => cmd_rdadcbuf_23
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__24314\,
            I => cmd_rdadcbuf_23
        );

    \I__3280\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24305\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24302\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__24305\,
            I => buf_adcdata_vdc_7
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__24302\,
            I => buf_adcdata_vdc_7
        );

    \I__3276\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24294\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24289\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24293\,
            I => \N__24286\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24283\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__24289\,
            I => \N__24280\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24277\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__24283\,
            I => buf_adcdata_vac_7
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__24280\,
            I => buf_adcdata_vac_7
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__24277\,
            I => buf_adcdata_vac_7
        );

    \I__3267\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24266\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24263\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__24266\,
            I => cmd_rdadcbuf_20
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__24263\,
            I => cmd_rdadcbuf_20
        );

    \I__3263\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24254\
        );

    \I__3262\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24251\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__24254\,
            I => cmd_rdadcbuf_22
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__24251\,
            I => cmd_rdadcbuf_22
        );

    \I__3259\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24242\
        );

    \I__3258\ : InMux
    port map (
            O => \N__24245\,
            I => \N__24239\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__24242\,
            I => cmd_rdadcbuf_28
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__24239\,
            I => cmd_rdadcbuf_28
        );

    \I__3255\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24230\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24227\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24223\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24227\,
            I => \N__24220\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24217\
        );

    \I__3250\ : Span12Mux_h
    port map (
            O => \N__24223\,
            I => \N__24212\
        );

    \I__3249\ : Sp12to4
    port map (
            O => \N__24220\,
            I => \N__24212\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__24217\,
            I => cmd_rdadcbuf_34
        );

    \I__3247\ : Odrv12
    port map (
            O => \N__24212\,
            I => cmd_rdadcbuf_34
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__24207\,
            I => \N__24203\
        );

    \I__3245\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24200\
        );

    \I__3244\ : InMux
    port map (
            O => \N__24203\,
            I => \N__24197\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__24200\,
            I => buf_adcdata_vdc_23
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__24197\,
            I => buf_adcdata_vdc_23
        );

    \I__3241\ : InMux
    port map (
            O => \N__24192\,
            I => \N__24189\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__24189\,
            I => \N__24186\
        );

    \I__3239\ : Span12Mux_s8_h
    port map (
            O => \N__24186\,
            I => \N__24181\
        );

    \I__3238\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24178\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24175\
        );

    \I__3236\ : Span12Mux_h
    port map (
            O => \N__24181\,
            I => \N__24172\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__24178\,
            I => \N__24169\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__24175\,
            I => buf_adcdata_vac_23
        );

    \I__3233\ : Odrv12
    port map (
            O => \N__24172\,
            I => buf_adcdata_vac_23
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__24169\,
            I => buf_adcdata_vac_23
        );

    \I__3231\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24157\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__24161\,
            I => \N__24154\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__24160\,
            I => \N__24151\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__24157\,
            I => \N__24148\
        );

    \I__3227\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24145\
        );

    \I__3226\ : InMux
    port map (
            O => \N__24151\,
            I => \N__24142\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__24148\,
            I => cmd_rdadctmp_5_adj_1474
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__24145\,
            I => cmd_rdadctmp_5_adj_1474
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__24142\,
            I => cmd_rdadctmp_5_adj_1474
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__3221\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24128\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__24131\,
            I => \N__24124\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24121\
        );

    \I__3218\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24118\
        );

    \I__3217\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24115\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__24121\,
            I => cmd_rdadctmp_6_adj_1473
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__24118\,
            I => cmd_rdadctmp_6_adj_1473
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__24115\,
            I => cmd_rdadctmp_6_adj_1473
        );

    \I__3213\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24101\
        );

    \I__3212\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24101\
        );

    \I__3211\ : InMux
    port map (
            O => \N__24106\,
            I => \N__24098\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__24101\,
            I => cmd_rdadctmp_7_adj_1472
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__24098\,
            I => cmd_rdadctmp_7_adj_1472
        );

    \I__3208\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24089\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24086\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__24089\,
            I => cmd_rdadcbuf_15
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__24086\,
            I => cmd_rdadcbuf_15
        );

    \I__3204\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24077\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__24080\,
            I => \N__24074\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__24077\,
            I => \N__24071\
        );

    \I__3201\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24068\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__24071\,
            I => buf_adcdata_vdc_4
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__24068\,
            I => buf_adcdata_vdc_4
        );

    \I__3198\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24058\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__24062\,
            I => \N__24055\
        );

    \I__3196\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24052\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__24058\,
            I => \N__24049\
        );

    \I__3194\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24046\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__24052\,
            I => cmd_rdadctmp_12_adj_1467
        );

    \I__3192\ : Odrv12
    port map (
            O => \N__24049\,
            I => cmd_rdadctmp_12_adj_1467
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__24046\,
            I => cmd_rdadctmp_12_adj_1467
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__24039\,
            I => \N__24034\
        );

    \I__3189\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24031\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__24037\,
            I => \N__24028\
        );

    \I__3187\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24025\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__24031\,
            I => \N__24022\
        );

    \I__3185\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24019\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__24025\,
            I => cmd_rdadctmp_13_adj_1466
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__24022\,
            I => cmd_rdadctmp_13_adj_1466
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__24019\,
            I => cmd_rdadctmp_13_adj_1466
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__24012\,
            I => \N__24007\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__24011\,
            I => \N__24004\
        );

    \I__3179\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24001\
        );

    \I__3178\ : InMux
    port map (
            O => \N__24007\,
            I => \N__23998\
        );

    \I__3177\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23995\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__24001\,
            I => cmd_rdadctmp_9_adj_1470
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__23998\,
            I => cmd_rdadctmp_9_adj_1470
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__23995\,
            I => cmd_rdadctmp_9_adj_1470
        );

    \I__3173\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23984\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__23987\,
            I => \N__23980\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23977\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23974\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23980\,
            I => \N__23971\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__23977\,
            I => cmd_rdadctmp_10_adj_1469
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23974\,
            I => cmd_rdadctmp_10_adj_1469
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__23971\,
            I => cmd_rdadctmp_10_adj_1469
        );

    \I__3165\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23961\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__23961\,
            I => \N__23957\
        );

    \I__3163\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23954\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__23957\,
            I => cmd_rdadcbuf_14
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__23954\,
            I => cmd_rdadcbuf_14
        );

    \I__3160\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23945\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__23948\,
            I => \N__23941\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23938\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23935\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23932\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__23938\,
            I => cmd_rdadctmp_15_adj_1464
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__23935\,
            I => cmd_rdadctmp_15_adj_1464
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__23932\,
            I => cmd_rdadctmp_15_adj_1464
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__23925\,
            I => \N__23922\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23918\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23914\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23918\,
            I => \N__23911\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__23917\,
            I => \N__23908\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23914\,
            I => \N__23903\
        );

    \I__3146\ : Span4Mux_v
    port map (
            O => \N__23911\,
            I => \N__23903\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23900\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__23903\,
            I => cmd_rdadctmp_16_adj_1463
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__23900\,
            I => cmd_rdadctmp_16_adj_1463
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__23895\,
            I => \N__23884\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__23894\,
            I => \N__23881\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__23893\,
            I => \N__23877\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__23892\,
            I => \N__23873\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__23891\,
            I => \N__23870\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__23890\,
            I => \N__23866\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__23889\,
            I => \N__23863\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__23888\,
            I => \N__23857\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23852\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23852\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23841\
        );

    \I__3131\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23841\
        );

    \I__3130\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23841\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23841\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23841\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23820\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23820\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23820\
        );

    \I__3124\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23820\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23820\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23820\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23820\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23820\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__23852\,
            I => \N__23815\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23841\,
            I => \N__23815\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__23840\,
            I => \N__23811\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__23839\,
            I => \N__23808\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__23838\,
            I => \N__23804\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__23837\,
            I => \N__23801\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__23820\,
            I => \N__23797\
        );

    \I__3112\ : Span4Mux_v
    port map (
            O => \N__23815\,
            I => \N__23794\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23787\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23787\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23787\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23784\
        );

    \I__3107\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23777\
        );

    \I__3106\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23777\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23777\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__23797\,
            I => n12871
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__23794\,
            I => n12871
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__23787\,
            I => n12871
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__23784\,
            I => n12871
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__23777\,
            I => n12871
        );

    \I__3099\ : InMux
    port map (
            O => \N__23766\,
            I => \N__23763\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23763\,
            I => \N__23758\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__23762\,
            I => \N__23755\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23752\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__23758\,
            I => \N__23749\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23746\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__23752\,
            I => cmd_rdadctmp_18_adj_1461
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__23749\,
            I => cmd_rdadctmp_18_adj_1461
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23746\,
            I => cmd_rdadctmp_18_adj_1461
        );

    \I__3090\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23731\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__23735\,
            I => \N__23728\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__23734\,
            I => \N__23725\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__23731\,
            I => \N__23722\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23719\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23716\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__23722\,
            I => cmd_rdadctmp_19_adj_1460
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23719\,
            I => cmd_rdadctmp_19_adj_1460
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__23716\,
            I => cmd_rdadctmp_19_adj_1460
        );

    \I__3080\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23706\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__23706\,
            I => \N__23702\
        );

    \I__3078\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23699\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__23702\,
            I => cmd_rdadcbuf_25
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__23699\,
            I => cmd_rdadcbuf_25
        );

    \I__3075\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23691\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23687\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23684\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__23687\,
            I => cmd_rdadcbuf_19
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__23684\,
            I => cmd_rdadcbuf_19
        );

    \I__3070\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23676\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__23673\,
            I => \N__23669\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__23672\,
            I => \N__23666\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__23669\,
            I => \N__23663\
        );

    \I__3065\ : InMux
    port map (
            O => \N__23666\,
            I => \N__23660\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__23663\,
            I => buf_adcdata_vdc_8
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__23660\,
            I => buf_adcdata_vdc_8
        );

    \I__3062\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23651\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23648\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__23651\,
            I => cmd_rdadcbuf_12
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__23648\,
            I => cmd_rdadcbuf_12
        );

    \I__3058\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23639\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23636\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__23639\,
            I => cmd_rdadcbuf_13
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__23636\,
            I => cmd_rdadcbuf_13
        );

    \I__3054\ : InMux
    port map (
            O => \N__23631\,
            I => \N__23627\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__23630\,
            I => \N__23623\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__23627\,
            I => \N__23620\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__23626\,
            I => \N__23617\
        );

    \I__3050\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23614\
        );

    \I__3049\ : Span4Mux_v
    port map (
            O => \N__23620\,
            I => \N__23611\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23608\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__23614\,
            I => cmd_rdadctmp_14_adj_1465
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__23611\,
            I => cmd_rdadctmp_14_adj_1465
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__23608\,
            I => cmd_rdadctmp_14_adj_1465
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__23601\,
            I => \N__23596\
        );

    \I__3043\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23593\
        );

    \I__3042\ : InMux
    port map (
            O => \N__23599\,
            I => \N__23590\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23587\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__23593\,
            I => cmd_rdadctmp_3_adj_1476
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__23590\,
            I => cmd_rdadctmp_3_adj_1476
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__23587\,
            I => cmd_rdadctmp_3_adj_1476
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__23580\,
            I => \N__23575\
        );

    \I__3036\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23572\
        );

    \I__3035\ : InMux
    port map (
            O => \N__23578\,
            I => \N__23569\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23566\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__23572\,
            I => cmd_rdadctmp_4_adj_1475
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__23569\,
            I => cmd_rdadctmp_4_adj_1475
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__23566\,
            I => cmd_rdadctmp_4_adj_1475
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__23559\,
            I => \N__23554\
        );

    \I__3029\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23551\
        );

    \I__3028\ : InMux
    port map (
            O => \N__23557\,
            I => \N__23548\
        );

    \I__3027\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23545\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__23551\,
            I => cmd_rdadctmp_8_adj_1471
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__23548\,
            I => cmd_rdadctmp_8_adj_1471
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__23545\,
            I => cmd_rdadctmp_8_adj_1471
        );

    \I__3023\ : InMux
    port map (
            O => \N__23538\,
            I => \N__23534\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23531\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__23534\,
            I => cmd_rdadcbuf_18
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__23531\,
            I => cmd_rdadcbuf_18
        );

    \I__3019\ : InMux
    port map (
            O => \N__23526\,
            I => \ADC_IAC.n19654\
        );

    \I__3018\ : InMux
    port map (
            O => \N__23523\,
            I => \ADC_IAC.n19655\
        );

    \I__3017\ : SRMux
    port map (
            O => \N__23520\,
            I => \N__23517\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__23517\,
            I => \N__23514\
        );

    \I__3015\ : Sp12to4
    port map (
            O => \N__23514\,
            I => \N__23511\
        );

    \I__3014\ : Odrv12
    port map (
            O => \N__23511\,
            I => \ADC_IAC.n14806\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__23508\,
            I => \ADC_IAC.n17_cascade_\
        );

    \I__3012\ : CEMux
    port map (
            O => \N__23505\,
            I => \N__23502\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__23502\,
            I => \ADC_IAC.n12\
        );

    \I__3010\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23495\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23498\,
            I => \N__23492\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__23495\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__23492\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__3006\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23483\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23480\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__23483\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__23480\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__23475\,
            I => \N__23471\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23468\
        );

    \I__3000\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23465\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__23468\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__23465\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__2997\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23456\
        );

    \I__2996\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23453\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__23456\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__23453\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__2993\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23445\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__23445\,
            I => \ADC_VDC.n20\
        );

    \I__2991\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23438\
        );

    \I__2990\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23435\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__23438\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__23435\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__2987\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23426\
        );

    \I__2986\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23423\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__23426\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23423\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__23418\,
            I => \N__23414\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23411\
        );

    \I__2981\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23408\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__23411\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__23408\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__2978\ : InMux
    port map (
            O => \N__23403\,
            I => \N__23399\
        );

    \I__2977\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23396\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__23399\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__23396\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__2974\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__23388\,
            I => \ADC_VDC.n21\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__23382\,
            I => \N__23379\
        );

    \I__2970\ : Span4Mux_h
    port map (
            O => \N__23379\,
            I => \N__23375\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23372\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__23375\,
            I => cmd_rdadcbuf_27
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__23372\,
            I => cmd_rdadcbuf_27
        );

    \I__2966\ : InMux
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__23364\,
            I => \N__23360\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__23363\,
            I => \N__23357\
        );

    \I__2963\ : Sp12to4
    port map (
            O => \N__23360\,
            I => \N__23354\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23351\
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__23354\,
            I => buf_adcdata_vdc_16
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__23351\,
            I => buf_adcdata_vdc_16
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__23346\,
            I => \N__23343\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23340\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__23340\,
            I => \N__23335\
        );

    \I__2956\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23330\
        );

    \I__2955\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23330\
        );

    \I__2954\ : Span4Mux_v
    port map (
            O => \N__23335\,
            I => \N__23327\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__23330\,
            I => cmd_rdadctmp_18
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__23327\,
            I => cmd_rdadctmp_18
        );

    \I__2951\ : IoInMux
    port map (
            O => \N__23322\,
            I => \N__23319\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__23319\,
            I => \N__23316\
        );

    \I__2949\ : IoSpan4Mux
    port map (
            O => \N__23316\,
            I => \N__23313\
        );

    \I__2948\ : Span4Mux_s3_v
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__2947\ : Sp12to4
    port map (
            O => \N__23310\,
            I => \N__23307\
        );

    \I__2946\ : Span12Mux_s10_v
    port map (
            O => \N__23307\,
            I => \N__23303\
        );

    \I__2945\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23300\
        );

    \I__2944\ : Odrv12
    port map (
            O => \N__23303\,
            I => \IAC_SCLK\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__23300\,
            I => \IAC_SCLK\
        );

    \I__2942\ : InMux
    port map (
            O => \N__23295\,
            I => \bfn_8_17_0_\
        );

    \I__2941\ : InMux
    port map (
            O => \N__23292\,
            I => \ADC_IAC.n19649\
        );

    \I__2940\ : InMux
    port map (
            O => \N__23289\,
            I => \ADC_IAC.n19650\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23286\,
            I => \ADC_IAC.n19651\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23283\,
            I => \ADC_IAC.n19652\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23280\,
            I => \ADC_IAC.n19653\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__23277\,
            I => \N__23273\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23270\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23267\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__23270\,
            I => \buf_readRTD_8\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__23267\,
            I => \buf_readRTD_8\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__23262\,
            I => \N__23258\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23254\
        );

    \I__2929\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23251\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__23257\,
            I => \N__23248\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__23254\,
            I => \N__23245\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23242\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23239\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__23245\,
            I => \N__23236\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__23242\,
            I => \N__23233\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__23239\,
            I => \N__23230\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__23236\,
            I => \N__23227\
        );

    \I__2920\ : Span4Mux_v
    port map (
            O => \N__23233\,
            I => \N__23224\
        );

    \I__2919\ : Span4Mux_h
    port map (
            O => \N__23230\,
            I => \N__23221\
        );

    \I__2918\ : Span4Mux_v
    port map (
            O => \N__23227\,
            I => \N__23216\
        );

    \I__2917\ : Span4Mux_h
    port map (
            O => \N__23224\,
            I => \N__23213\
        );

    \I__2916\ : Span4Mux_v
    port map (
            O => \N__23221\,
            I => \N__23210\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23205\
        );

    \I__2914\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23205\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__23216\,
            I => \buf_cfgRTD_0\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__23213\,
            I => \buf_cfgRTD_0\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__23210\,
            I => \buf_cfgRTD_0\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__23205\,
            I => \buf_cfgRTD_0\
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__23196\,
            I => \N__23193\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23190\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__23190\,
            I => n21202
        );

    \I__2906\ : IoInMux
    port map (
            O => \N__23187\,
            I => \N__23184\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__23184\,
            I => \N__23181\
        );

    \I__2904\ : Span4Mux_s0_h
    port map (
            O => \N__23181\,
            I => \N__23178\
        );

    \I__2903\ : Sp12to4
    port map (
            O => \N__23178\,
            I => \N__23175\
        );

    \I__2902\ : Span12Mux_s11_v
    port map (
            O => \N__23175\,
            I => \N__23170\
        );

    \I__2901\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23167\
        );

    \I__2900\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23164\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__23170\,
            I => \VAC_OSR1\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__23167\,
            I => \VAC_OSR1\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__23164\,
            I => \VAC_OSR1\
        );

    \I__2896\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23153\
        );

    \I__2895\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23150\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__23153\,
            I => \N__23147\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__23150\,
            I => \N__23144\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__23147\,
            I => \N__23140\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__23144\,
            I => \N__23137\
        );

    \I__2890\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23134\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__23140\,
            I => cmd_rdadctmp_16
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__23137\,
            I => cmd_rdadctmp_16
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__23134\,
            I => cmd_rdadctmp_16
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__23127\,
            I => \N__23124\
        );

    \I__2885\ : InMux
    port map (
            O => \N__23124\,
            I => \N__23117\
        );

    \I__2884\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23117\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__23122\,
            I => \N__23114\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23111\
        );

    \I__2881\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23108\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__23111\,
            I => cmd_rdadctmp_17
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__23108\,
            I => cmd_rdadctmp_17
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__23103\,
            I => \N__23096\
        );

    \I__2877\ : InMux
    port map (
            O => \N__23102\,
            I => \N__23093\
        );

    \I__2876\ : InMux
    port map (
            O => \N__23101\,
            I => \N__23090\
        );

    \I__2875\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23087\
        );

    \I__2874\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23084\
        );

    \I__2873\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23081\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__23072\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__23090\,
            I => \N__23072\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__23087\,
            I => \N__23072\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23072\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__23081\,
            I => \N__23069\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__23072\,
            I => \N__23066\
        );

    \I__2866\ : Span12Mux_v
    port map (
            O => \N__23069\,
            I => \N__23061\
        );

    \I__2865\ : Sp12to4
    port map (
            O => \N__23066\,
            I => \N__23061\
        );

    \I__2864\ : Odrv12
    port map (
            O => \N__23061\,
            I => \VAC_DRDY\
        );

    \I__2863\ : IoInMux
    port map (
            O => \N__23058\,
            I => \N__23055\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__23055\,
            I => \N__23052\
        );

    \I__2861\ : Span12Mux_s8_h
    port map (
            O => \N__23052\,
            I => \N__23048\
        );

    \I__2860\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23044\
        );

    \I__2859\ : Span12Mux_v
    port map (
            O => \N__23048\,
            I => \N__23041\
        );

    \I__2858\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23038\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__23035\
        );

    \I__2856\ : Odrv12
    port map (
            O => \N__23041\,
            I => \AMPV_POW\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__23038\,
            I => \AMPV_POW\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__23035\,
            I => \AMPV_POW\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__23028\,
            I => \n23_adj_1540_cascade_\
        );

    \I__2852\ : InMux
    port map (
            O => \N__23025\,
            I => \N__23022\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__23022\,
            I => n21123
        );

    \I__2850\ : InMux
    port map (
            O => \N__23019\,
            I => \N__23016\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__23016\,
            I => \N__23013\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__23013\,
            I => \N__23010\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__2846\ : Span12Mux_h
    port map (
            O => \N__23007\,
            I => \N__23004\
        );

    \I__2845\ : Span12Mux_v
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__2844\ : Odrv12
    port map (
            O => \N__23001\,
            I => \EIS_SYNCCLK\
        );

    \I__2843\ : IoInMux
    port map (
            O => \N__22998\,
            I => \N__22995\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__22995\,
            I => \N__22991\
        );

    \I__2841\ : IoInMux
    port map (
            O => \N__22994\,
            I => \N__22988\
        );

    \I__2840\ : IoSpan4Mux
    port map (
            O => \N__22991\,
            I => \N__22985\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22982\
        );

    \I__2838\ : Span4Mux_s2_h
    port map (
            O => \N__22985\,
            I => \N__22979\
        );

    \I__2837\ : IoSpan4Mux
    port map (
            O => \N__22982\,
            I => \N__22976\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__22979\,
            I => \N__22973\
        );

    \I__2835\ : Span4Mux_s2_v
    port map (
            O => \N__22976\,
            I => \N__22970\
        );

    \I__2834\ : Span4Mux_h
    port map (
            O => \N__22973\,
            I => \N__22967\
        );

    \I__2833\ : Sp12to4
    port map (
            O => \N__22970\,
            I => \N__22964\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__22967\,
            I => \N__22961\
        );

    \I__2831\ : Odrv12
    port map (
            O => \N__22964\,
            I => \IAC_CLK\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__22961\,
            I => \IAC_CLK\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__22956\,
            I => \N__22953\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22950\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__2826\ : Span4Mux_h
    port map (
            O => \N__22947\,
            I => \N__22942\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22937\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22937\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__22942\,
            I => cmd_rdadctmp_15
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22937\,
            I => cmd_rdadctmp_15
        );

    \I__2821\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22929\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__2819\ : Span4Mux_h
    port map (
            O => \N__22926\,
            I => \N__22923\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__22923\,
            I => n21082
        );

    \I__2817\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22917\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__22917\,
            I => \N__22914\
        );

    \I__2815\ : Odrv12
    port map (
            O => \N__22914\,
            I => n21201
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__22911\,
            I => \n22315_cascade_\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22905\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__22905\,
            I => n22318
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__22902\,
            I => \N__22899\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22896\,
            I => \N__22892\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__22895\,
            I => \N__22888\
        );

    \I__2807\ : Span4Mux_h
    port map (
            O => \N__22892\,
            I => \N__22885\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22880\
        );

    \I__2805\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22880\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__22885\,
            I => cmd_rdadctmp_22
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__22880\,
            I => cmd_rdadctmp_22
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__22875\,
            I => \N__22871\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__22874\,
            I => \N__22868\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22865\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22862\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__22865\,
            I => cmd_rdadctmp_31_adj_1419
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__22862\,
            I => cmd_rdadctmp_31_adj_1419
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__22857\,
            I => \N__22852\
        );

    \I__2795\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22847\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22847\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22844\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__22847\,
            I => cmd_rdadctmp_30_adj_1420
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22844\,
            I => cmd_rdadctmp_30_adj_1420
        );

    \I__2790\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__22833\,
            I => n22405
        );

    \I__2787\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22827\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22827\,
            I => \N__22824\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__22824\,
            I => \N__22821\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__22821\,
            I => \N__22817\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__22820\,
            I => \N__22814\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__22817\,
            I => \N__22811\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22807\
        );

    \I__2780\ : Span4Mux_h
    port map (
            O => \N__22811\,
            I => \N__22804\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22801\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__22807\,
            I => \N__22798\
        );

    \I__2777\ : Span4Mux_h
    port map (
            O => \N__22804\,
            I => \N__22795\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__22801\,
            I => buf_adcdata_vac_21
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__22798\,
            I => buf_adcdata_vac_21
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__22795\,
            I => buf_adcdata_vac_21
        );

    \I__2773\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22785\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__22785\,
            I => n21097
        );

    \I__2771\ : InMux
    port map (
            O => \N__22782\,
            I => \N__22778\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__22781\,
            I => \N__22774\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__22778\,
            I => \N__22771\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22768\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22765\
        );

    \I__2766\ : Sp12to4
    port map (
            O => \N__22771\,
            I => \N__22760\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__22768\,
            I => \N__22760\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__22765\,
            I => \N__22757\
        );

    \I__2763\ : Span12Mux_v
    port map (
            O => \N__22760\,
            I => \N__22752\
        );

    \I__2762\ : Span4Mux_h
    port map (
            O => \N__22757\,
            I => \N__22749\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22744\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22744\
        );

    \I__2759\ : Odrv12
    port map (
            O => \N__22752\,
            I => \buf_cfgRTD_4\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__22749\,
            I => \buf_cfgRTD_4\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__22744\,
            I => \buf_cfgRTD_4\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22731\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__2753\ : Span4Mux_h
    port map (
            O => \N__22728\,
            I => \N__22724\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__22727\,
            I => \N__22721\
        );

    \I__2751\ : Span4Mux_v
    port map (
            O => \N__22724\,
            I => \N__22718\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22715\
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__22718\,
            I => \buf_readRTD_12\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__22715\,
            I => \buf_readRTD_12\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__22710\,
            I => \N__22707\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22701\
        );

    \I__2744\ : Span4Mux_v
    port map (
            O => \N__22701\,
            I => \N__22697\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \N__22694\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__22697\,
            I => \N__22691\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22688\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__22691\,
            I => \buf_readRTD_4\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__22688\,
            I => \buf_readRTD_4\
        );

    \I__2738\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22676\
        );

    \I__2736\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22672\
        );

    \I__2735\ : Span12Mux_h
    port map (
            O => \N__22676\,
            I => \N__22669\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22666\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__22672\,
            I => buf_adcdata_vac_16
        );

    \I__2732\ : Odrv12
    port map (
            O => \N__22669\,
            I => buf_adcdata_vac_16
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__22666\,
            I => buf_adcdata_vac_16
        );

    \I__2730\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22652\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__22655\,
            I => \N__22649\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__22652\,
            I => \N__22646\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22643\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__22646\,
            I => cmd_rdadctmp_3
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22643\,
            I => cmd_rdadctmp_3
        );

    \I__2723\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22633\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__22637\,
            I => \N__22630\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22627\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__22633\,
            I => \N__22624\
        );

    \I__2719\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22621\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__22627\,
            I => cmd_rdadctmp_27_adj_1423
        );

    \I__2717\ : Odrv12
    port map (
            O => \N__22624\,
            I => cmd_rdadctmp_27_adj_1423
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__22621\,
            I => cmd_rdadctmp_27_adj_1423
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__22614\,
            I => \N__22609\
        );

    \I__2714\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22606\
        );

    \I__2713\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22601\
        );

    \I__2712\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22601\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__22606\,
            I => cmd_rdadctmp_28_adj_1422
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__22601\,
            I => cmd_rdadctmp_28_adj_1422
        );

    \I__2709\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22592\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__22595\,
            I => \N__22589\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22592\,
            I => \N__22586\
        );

    \I__2706\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22582\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__22586\,
            I => \N__22579\
        );

    \I__2704\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22576\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__22582\,
            I => cmd_rdadctmp_29_adj_1421
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__22579\,
            I => cmd_rdadctmp_29_adj_1421
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__22576\,
            I => cmd_rdadctmp_29_adj_1421
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__22569\,
            I => \N__22566\
        );

    \I__2699\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22563\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__22563\,
            I => \N__22559\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__22562\,
            I => \N__22556\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__22559\,
            I => \N__22553\
        );

    \I__2695\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22550\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__22553\,
            I => cmd_rdadctmp_7_adj_1443
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__22550\,
            I => cmd_rdadctmp_7_adj_1443
        );

    \I__2692\ : InMux
    port map (
            O => \N__22545\,
            I => \ADC_VDC.n19688\
        );

    \I__2691\ : InMux
    port map (
            O => \N__22542\,
            I => \ADC_VDC.n19689\
        );

    \I__2690\ : InMux
    port map (
            O => \N__22539\,
            I => \ADC_VDC.n19690\
        );

    \I__2689\ : InMux
    port map (
            O => \N__22536\,
            I => \ADC_VDC.n19691\
        );

    \I__2688\ : InMux
    port map (
            O => \N__22533\,
            I => \ADC_VDC.n19692\
        );

    \I__2687\ : InMux
    port map (
            O => \N__22530\,
            I => \ADC_VDC.n19693\
        );

    \I__2686\ : InMux
    port map (
            O => \N__22527\,
            I => \bfn_8_10_0_\
        );

    \I__2685\ : InMux
    port map (
            O => \N__22524\,
            I => \ADC_VDC.n19695\
        );

    \I__2684\ : CEMux
    port map (
            O => \N__22521\,
            I => \N__22516\
        );

    \I__2683\ : CEMux
    port map (
            O => \N__22520\,
            I => \N__22510\
        );

    \I__2682\ : CEMux
    port map (
            O => \N__22519\,
            I => \N__22507\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__22516\,
            I => \N__22503\
        );

    \I__2680\ : CEMux
    port map (
            O => \N__22515\,
            I => \N__22500\
        );

    \I__2679\ : CEMux
    port map (
            O => \N__22514\,
            I => \N__22497\
        );

    \I__2678\ : CEMux
    port map (
            O => \N__22513\,
            I => \N__22494\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__22510\,
            I => \N__22489\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__22507\,
            I => \N__22489\
        );

    \I__2675\ : CEMux
    port map (
            O => \N__22506\,
            I => \N__22486\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__22503\,
            I => \N__22483\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__22500\,
            I => \N__22480\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__22497\,
            I => \N__22477\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22474\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__22489\,
            I => \N__22467\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22467\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__22483\,
            I => \N__22467\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__22480\,
            I => \N__22462\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__22477\,
            I => \N__22462\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__22474\,
            I => \ADC_VDC.n13010\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__22467\,
            I => \ADC_VDC.n13010\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__22462\,
            I => \ADC_VDC.n13010\
        );

    \I__2662\ : SRMux
    port map (
            O => \N__22455\,
            I => \N__22448\
        );

    \I__2661\ : SRMux
    port map (
            O => \N__22454\,
            I => \N__22444\
        );

    \I__2660\ : SRMux
    port map (
            O => \N__22453\,
            I => \N__22440\
        );

    \I__2659\ : SRMux
    port map (
            O => \N__22452\,
            I => \N__22437\
        );

    \I__2658\ : SRMux
    port map (
            O => \N__22451\,
            I => \N__22434\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__22448\,
            I => \N__22431\
        );

    \I__2656\ : SRMux
    port map (
            O => \N__22447\,
            I => \N__22428\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__22444\,
            I => \N__22425\
        );

    \I__2654\ : SRMux
    port map (
            O => \N__22443\,
            I => \N__22422\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__22440\,
            I => \N__22419\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22416\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__22434\,
            I => \N__22413\
        );

    \I__2650\ : Span4Mux_v
    port map (
            O => \N__22431\,
            I => \N__22408\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22428\,
            I => \N__22408\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__22425\,
            I => \N__22401\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__22422\,
            I => \N__22401\
        );

    \I__2646\ : Span4Mux_h
    port map (
            O => \N__22419\,
            I => \N__22401\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__22416\,
            I => \N__22398\
        );

    \I__2644\ : Odrv12
    port map (
            O => \N__22413\,
            I => \ADC_VDC.n14915\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__22408\,
            I => \ADC_VDC.n14915\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__22401\,
            I => \ADC_VDC.n14915\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__22398\,
            I => \ADC_VDC.n14915\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22389\,
            I => \ADC_VDC.n19696\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22383\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22380\
        );

    \I__2637\ : Odrv12
    port map (
            O => \N__22380\,
            I => \ADC_VDC.cmd_rdadcbuf_35_N_1138_34\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__22377\,
            I => \N__22372\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22367\
        );

    \I__2634\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22367\
        );

    \I__2633\ : InMux
    port map (
            O => \N__22372\,
            I => \N__22364\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__22367\,
            I => cmd_rdadctmp_17_adj_1462
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__22364\,
            I => cmd_rdadctmp_17_adj_1462
        );

    \I__2630\ : InMux
    port map (
            O => \N__22359\,
            I => \ADC_VDC.n19679\
        );

    \I__2629\ : InMux
    port map (
            O => \N__22356\,
            I => \ADC_VDC.n19680\
        );

    \I__2628\ : InMux
    port map (
            O => \N__22353\,
            I => \ADC_VDC.n19681\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__22350\,
            I => \N__22346\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__22349\,
            I => \N__22342\
        );

    \I__2625\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22339\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22336\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22333\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__22339\,
            I => cmd_rdadctmp_20_adj_1459
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__22336\,
            I => cmd_rdadctmp_20_adj_1459
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__22333\,
            I => cmd_rdadctmp_20_adj_1459
        );

    \I__2619\ : InMux
    port map (
            O => \N__22326\,
            I => \ADC_VDC.n19682\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__22323\,
            I => \N__22318\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22313\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22313\
        );

    \I__2615\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22310\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__22313\,
            I => cmd_rdadctmp_21_adj_1458
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__22310\,
            I => cmd_rdadctmp_21_adj_1458
        );

    \I__2612\ : InMux
    port map (
            O => \N__22305\,
            I => \ADC_VDC.n19683\
        );

    \I__2611\ : InMux
    port map (
            O => \N__22302\,
            I => \ADC_VDC.n19684\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22299\,
            I => \ADC_VDC.n19685\
        );

    \I__2609\ : InMux
    port map (
            O => \N__22296\,
            I => \bfn_8_9_0_\
        );

    \I__2608\ : InMux
    port map (
            O => \N__22293\,
            I => \ADC_VDC.n19687\
        );

    \I__2607\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22287\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__22287\,
            I => \ADC_VDC.cmd_rdadcbuf_9\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22284\,
            I => \ADC_VDC.n19671\
        );

    \I__2604\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22278\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__22278\,
            I => \ADC_VDC.cmd_rdadcbuf_10\
        );

    \I__2602\ : InMux
    port map (
            O => \N__22275\,
            I => \ADC_VDC.n19672\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__22272\,
            I => \N__22268\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__22271\,
            I => \N__22264\
        );

    \I__2599\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22259\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22259\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22256\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__22259\,
            I => cmd_rdadctmp_11_adj_1468
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__22256\,
            I => cmd_rdadctmp_11_adj_1468
        );

    \I__2594\ : InMux
    port map (
            O => \N__22251\,
            I => \ADC_VDC.n19673\
        );

    \I__2593\ : InMux
    port map (
            O => \N__22248\,
            I => \ADC_VDC.n19674\
        );

    \I__2592\ : InMux
    port map (
            O => \N__22245\,
            I => \ADC_VDC.n19675\
        );

    \I__2591\ : InMux
    port map (
            O => \N__22242\,
            I => \ADC_VDC.n19676\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22239\,
            I => \ADC_VDC.n19677\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22233\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__22233\,
            I => \N__22229\
        );

    \I__2587\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22226\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__22229\,
            I => cmd_rdadcbuf_16
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__22226\,
            I => cmd_rdadcbuf_16
        );

    \I__2584\ : InMux
    port map (
            O => \N__22221\,
            I => \bfn_8_8_0_\
        );

    \I__2583\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22215\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__22215\,
            I => \ADC_VDC.cmd_rdadcbuf_0\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__22212\,
            I => \N__22207\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22202\
        );

    \I__2579\ : InMux
    port map (
            O => \N__22210\,
            I => \N__22202\
        );

    \I__2578\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22199\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__22202\,
            I => cmd_rdadctmp_1_adj_1478
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__22199\,
            I => cmd_rdadctmp_1_adj_1478
        );

    \I__2575\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22191\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__22191\,
            I => \ADC_VDC.cmd_rdadcbuf_1\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22188\,
            I => \ADC_VDC.n19663\
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__22185\,
            I => \N__22180\
        );

    \I__2571\ : InMux
    port map (
            O => \N__22184\,
            I => \N__22175\
        );

    \I__2570\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22175\
        );

    \I__2569\ : InMux
    port map (
            O => \N__22180\,
            I => \N__22172\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__22175\,
            I => cmd_rdadctmp_2_adj_1477
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__22172\,
            I => cmd_rdadctmp_2_adj_1477
        );

    \I__2566\ : InMux
    port map (
            O => \N__22167\,
            I => \N__22164\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__22164\,
            I => \ADC_VDC.cmd_rdadcbuf_2\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22161\,
            I => \ADC_VDC.n19664\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22155\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__22155\,
            I => \ADC_VDC.cmd_rdadcbuf_3\
        );

    \I__2561\ : InMux
    port map (
            O => \N__22152\,
            I => \ADC_VDC.n19665\
        );

    \I__2560\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22146\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__22146\,
            I => \ADC_VDC.cmd_rdadcbuf_4\
        );

    \I__2558\ : InMux
    port map (
            O => \N__22143\,
            I => \ADC_VDC.n19666\
        );

    \I__2557\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__22137\,
            I => \ADC_VDC.cmd_rdadcbuf_5\
        );

    \I__2555\ : InMux
    port map (
            O => \N__22134\,
            I => \ADC_VDC.n19667\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22128\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__22128\,
            I => \ADC_VDC.cmd_rdadcbuf_6\
        );

    \I__2552\ : InMux
    port map (
            O => \N__22125\,
            I => \ADC_VDC.n19668\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__2550\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__22116\,
            I => \ADC_VDC.cmd_rdadcbuf_7\
        );

    \I__2548\ : InMux
    port map (
            O => \N__22113\,
            I => \ADC_VDC.n19669\
        );

    \I__2547\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__22107\,
            I => \ADC_VDC.cmd_rdadcbuf_8\
        );

    \I__2545\ : InMux
    port map (
            O => \N__22104\,
            I => \bfn_8_7_0_\
        );

    \I__2544\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22097\
        );

    \I__2543\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22094\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__22097\,
            I => \N__22091\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__22094\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__22091\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__2539\ : InMux
    port map (
            O => \N__22086\,
            I => \ADC_VDC.n19707\
        );

    \I__2538\ : InMux
    port map (
            O => \N__22083\,
            I => \ADC_VDC.n19708\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__22080\,
            I => \ADC_VDC.n13010_cascade_\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__22077\,
            I => \n12871_cascade_\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__22074\,
            I => \N__22069\
        );

    \I__2534\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22064\
        );

    \I__2533\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22064\
        );

    \I__2532\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22061\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__22064\,
            I => cmd_rdadctmp_0_adj_1479
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__22061\,
            I => cmd_rdadctmp_0_adj_1479
        );

    \I__2529\ : InMux
    port map (
            O => \N__22056\,
            I => \ADC_VDC.n19698\
        );

    \I__2528\ : InMux
    port map (
            O => \N__22053\,
            I => \ADC_VDC.n19699\
        );

    \I__2527\ : InMux
    port map (
            O => \N__22050\,
            I => \ADC_VDC.n19700\
        );

    \I__2526\ : InMux
    port map (
            O => \N__22047\,
            I => \ADC_VDC.n19701\
        );

    \I__2525\ : InMux
    port map (
            O => \N__22044\,
            I => \ADC_VDC.n19702\
        );

    \I__2524\ : InMux
    port map (
            O => \N__22041\,
            I => \ADC_VDC.n19703\
        );

    \I__2523\ : InMux
    port map (
            O => \N__22038\,
            I => \ADC_VDC.n19704\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__22035\,
            I => \N__22032\
        );

    \I__2521\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22028\
        );

    \I__2520\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22025\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22022\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__22025\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__22022\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__2516\ : InMux
    port map (
            O => \N__22017\,
            I => \bfn_8_4_0_\
        );

    \I__2515\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22010\
        );

    \I__2514\ : InMux
    port map (
            O => \N__22013\,
            I => \N__22007\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__22004\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__22007\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__22004\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__2510\ : InMux
    port map (
            O => \N__21999\,
            I => \ADC_VDC.n19706\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__21996\,
            I => \ADC_VDC.n19_cascade_\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__21993\,
            I => \ADC_VDC.n18563_cascade_\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__21987\,
            I => \ADC_VDC.n18563\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__21984\,
            I => \ADC_VDC.n21384_cascade_\
        );

    \I__2504\ : CEMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__21975\,
            I => \ADC_VDC.n13034\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21968\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21965\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21968\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__21965\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21960\,
            I => \bfn_8_3_0_\
        );

    \I__2496\ : IoInMux
    port map (
            O => \N__21957\,
            I => \N__21954\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21954\,
            I => \N__21951\
        );

    \I__2494\ : IoSpan4Mux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__2493\ : Span4Mux_s3_h
    port map (
            O => \N__21948\,
            I => \N__21944\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__21947\,
            I => \N__21941\
        );

    \I__2491\ : Span4Mux_h
    port map (
            O => \N__21944\,
            I => \N__21938\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21935\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__21938\,
            I => \VAC_SCLK\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__21935\,
            I => \VAC_SCLK\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__21927\,
            I => \N__21923\
        );

    \I__2485\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21920\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__21923\,
            I => cmd_rdadctmp_5_adj_1445
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__21920\,
            I => cmd_rdadctmp_5_adj_1445
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__21915\,
            I => \N__21911\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21906\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21906\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21906\,
            I => cmd_rdadctmp_6_adj_1444
        );

    \I__2478\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21900\,
            I => \ADC_VAC.n21312\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__21897\,
            I => \ADC_VAC.n20958_cascade_\
        );

    \I__2475\ : CEMux
    port map (
            O => \N__21894\,
            I => \N__21891\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21891\,
            I => \N__21888\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__21888\,
            I => \N__21885\
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__21885\,
            I => \ADC_VAC.n20959\
        );

    \I__2471\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21878\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__21881\,
            I => \N__21874\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__21878\,
            I => \N__21871\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__21877\,
            I => \N__21868\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21865\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__21871\,
            I => \N__21862\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21859\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__21865\,
            I => \N__21856\
        );

    \I__2463\ : Span4Mux_h
    port map (
            O => \N__21862\,
            I => \N__21851\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__21859\,
            I => \N__21851\
        );

    \I__2461\ : Span4Mux_v
    port map (
            O => \N__21856\,
            I => \N__21848\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__21851\,
            I => \N__21845\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__21848\,
            I => \N__21840\
        );

    \I__2458\ : Sp12to4
    port map (
            O => \N__21845\,
            I => \N__21837\
        );

    \I__2457\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21834\
        );

    \I__2456\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21831\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__21840\,
            I => \buf_cfgRTD_2\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__21837\,
            I => \buf_cfgRTD_2\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__21834\,
            I => \buf_cfgRTD_2\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__21831\,
            I => \buf_cfgRTD_2\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__21822\,
            I => \N__21818\
        );

    \I__2450\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21815\
        );

    \I__2449\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21812\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N__21808\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N__21805\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__21811\,
            I => \N__21802\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__21808\,
            I => \N__21797\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__21805\,
            I => \N__21797\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21794\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__21797\,
            I => \N__21790\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__21794\,
            I => \N__21786\
        );

    \I__2440\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21783\
        );

    \I__2439\ : Span4Mux_h
    port map (
            O => \N__21790\,
            I => \N__21780\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21777\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__21786\,
            I => \N__21772\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__21783\,
            I => \N__21772\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__21780\,
            I => \buf_cfgRTD_5\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21777\,
            I => \buf_cfgRTD_5\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__21772\,
            I => \buf_cfgRTD_5\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21760\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__21764\,
            I => \N__21757\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__21763\,
            I => \N__21754\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__21760\,
            I => \N__21751\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21746\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21746\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__21751\,
            I => cmd_rdadctmp_24_adj_1426
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__21746\,
            I => cmd_rdadctmp_24_adj_1426
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__21741\,
            I => \n22321_cascade_\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21730\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21725\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21733\,
            I => \N__21725\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__21730\,
            I => read_buf_8
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__21725\,
            I => read_buf_8
        );

    \I__2417\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21713\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21713\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21705\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__21713\,
            I => \N__21698\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21693\
        );

    \I__2412\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21693\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21688\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21688\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21685\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__21705\,
            I => \N__21680\
        );

    \I__2407\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21671\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21671\
        );

    \I__2405\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21671\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21671\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__21698\,
            I => \N__21663\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__21693\,
            I => \N__21663\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__21688\,
            I => \N__21663\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21685\,
            I => \N__21660\
        );

    \I__2399\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21655\
        );

    \I__2398\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21655\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__21680\,
            I => \N__21650\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__21671\,
            I => \N__21650\
        );

    \I__2395\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21647\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__21663\,
            I => \N__21640\
        );

    \I__2393\ : Span4Mux_h
    port map (
            O => \N__21660\,
            I => \N__21640\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21655\,
            I => \N__21640\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__21650\,
            I => \N__21634\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__21647\,
            I => \N__21634\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__21640\,
            I => \N__21631\
        );

    \I__2388\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21628\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__21634\,
            I => \N__21625\
        );

    \I__2386\ : Span4Mux_h
    port map (
            O => \N__21631\,
            I => \N__21622\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__21628\,
            I => \N__21619\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__21625\,
            I => n11714
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__21622\,
            I => n11714
        );

    \I__2382\ : Odrv12
    port map (
            O => \N__21619\,
            I => n11714
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__21612\,
            I => \N__21608\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__21611\,
            I => \N__21605\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21602\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21599\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__21602\,
            I => \N__21596\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21593\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__21596\,
            I => \N__21589\
        );

    \I__2374\ : Span4Mux_h
    port map (
            O => \N__21593\,
            I => \N__21586\
        );

    \I__2373\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21583\
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__21589\,
            I => cmd_rdadctmp_13_adj_1437
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__21586\,
            I => cmd_rdadctmp_13_adj_1437
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__21583\,
            I => cmd_rdadctmp_13_adj_1437
        );

    \I__2369\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21570\
        );

    \I__2367\ : Span12Mux_s11_h
    port map (
            O => \N__21570\,
            I => \N__21565\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21562\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21559\
        );

    \I__2364\ : Span12Mux_v
    port map (
            O => \N__21565\,
            I => \N__21556\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21553\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__21559\,
            I => buf_adcdata_vac_8
        );

    \I__2361\ : Odrv12
    port map (
            O => \N__21556\,
            I => buf_adcdata_vac_8
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__21553\,
            I => buf_adcdata_vac_8
        );

    \I__2359\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21543\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21543\,
            I => \N__21539\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__21542\,
            I => \N__21535\
        );

    \I__2356\ : Span4Mux_h
    port map (
            O => \N__21539\,
            I => \N__21532\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21529\
        );

    \I__2354\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21526\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__21532\,
            I => \N__21523\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21520\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__21526\,
            I => buf_adcdata_vac_6
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__21523\,
            I => buf_adcdata_vac_6
        );

    \I__2349\ : Odrv12
    port map (
            O => \N__21520\,
            I => buf_adcdata_vac_6
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__21513\,
            I => \N__21509\
        );

    \I__2347\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21501\
        );

    \I__2346\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21501\
        );

    \I__2345\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21501\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__21501\,
            I => cmd_rdadctmp_14_adj_1436
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__21498\,
            I => \N__21495\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21489\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21489\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__21489\,
            I => \N__21486\
        );

    \I__2339\ : Span4Mux_h
    port map (
            O => \N__21486\,
            I => \N__21482\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21479\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__21482\,
            I => cmd_rdadctmp_15_adj_1435
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__21479\,
            I => cmd_rdadctmp_15_adj_1435
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__21474\,
            I => \N__21470\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__21473\,
            I => \N__21466\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21459\
        );

    \I__2332\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21459\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21459\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__21459\,
            I => cmd_rdadctmp_16_adj_1434
        );

    \I__2329\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21453\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__21453\,
            I => \N__21450\
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__21450\,
            I => buf_data_iac_4
        );

    \I__2326\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21444\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__21444\,
            I => n22_adj_1633
        );

    \I__2324\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21437\
        );

    \I__2323\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21434\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__21437\,
            I => bit_cnt_3
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21434\,
            I => bit_cnt_3
        );

    \I__2320\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21426\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21426\,
            I => n21456
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__21423\,
            I => \N__21417\
        );

    \I__2317\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21410\
        );

    \I__2316\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21410\
        );

    \I__2315\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21410\
        );

    \I__2314\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21407\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__21410\,
            I => bit_cnt_1
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__21407\,
            I => bit_cnt_1
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__21402\,
            I => \N__21399\
        );

    \I__2310\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21392\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21392\
        );

    \I__2308\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21389\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__21392\,
            I => bit_cnt_2
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__21389\,
            I => bit_cnt_2
        );

    \I__2305\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21381\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__21381\,
            I => n8_adj_1602
        );

    \I__2303\ : CEMux
    port map (
            O => \N__21378\,
            I => \N__21374\
        );

    \I__2302\ : CEMux
    port map (
            O => \N__21377\,
            I => \N__21371\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__21374\,
            I => \N__21368\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21365\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__21368\,
            I => \N__21362\
        );

    \I__2298\ : Odrv12
    port map (
            O => \N__21365\,
            I => \CLK_DDS.n9\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__21362\,
            I => \CLK_DDS.n9\
        );

    \I__2296\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21354\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__21354\,
            I => n19_adj_1626
        );

    \I__2294\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__21348\,
            I => n20867
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__21345\,
            I => \n20867_cascade_\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21339\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__21339\,
            I => \N__21336\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__21333\,
            I => \N__21330\
        );

    \I__2287\ : IoSpan4Mux
    port map (
            O => \N__21330\,
            I => \N__21327\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__21327\,
            I => \IAC_MISO\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__21324\,
            I => \n12498_cascade_\
        );

    \I__2284\ : InMux
    port map (
            O => \N__21321\,
            I => \N__21315\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21315\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__21315\,
            I => cmd_rdadctmp_0
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__21312\,
            I => \N__21308\
        );

    \I__2280\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21303\
        );

    \I__2279\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21303\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__21303\,
            I => cmd_rdadctmp_1
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__21300\,
            I => \N__21296\
        );

    \I__2276\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21293\
        );

    \I__2275\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21290\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21293\,
            I => \N__21287\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__21290\,
            I => cmd_rdadctmp_2
        );

    \I__2272\ : Odrv12
    port map (
            O => \N__21287\,
            I => cmd_rdadctmp_2
        );

    \I__2271\ : IoInMux
    port map (
            O => \N__21282\,
            I => \N__21279\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__21279\,
            I => \N__21276\
        );

    \I__2269\ : Span4Mux_s3_v
    port map (
            O => \N__21276\,
            I => \N__21273\
        );

    \I__2268\ : Span4Mux_h
    port map (
            O => \N__21273\,
            I => \N__21270\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__21270\,
            I => \N__21267\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__21267\,
            I => \AC_ADC_SYNC\
        );

    \I__2265\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21260\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__21263\,
            I => \N__21257\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__21260\,
            I => \N__21254\
        );

    \I__2262\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21251\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__21254\,
            I => buf_adcdata_vdc_5
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__21251\,
            I => buf_adcdata_vdc_5
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__21246\,
            I => \N__21242\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__21245\,
            I => \N__21239\
        );

    \I__2257\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21234\
        );

    \I__2256\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21234\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21234\,
            I => cmd_rdadctmp_4_adj_1446
        );

    \I__2254\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21228\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__21228\,
            I => n20864
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__21225\,
            I => \n20864_cascade_\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__21222\,
            I => \ADC_VAC.n17_cascade_\
        );

    \I__2250\ : CEMux
    port map (
            O => \N__21219\,
            I => \N__21216\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__21216\,
            I => \ADC_VAC.n12\
        );

    \I__2248\ : IoInMux
    port map (
            O => \N__21213\,
            I => \N__21210\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__2246\ : IoSpan4Mux
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__2245\ : Span4Mux_s2_v
    port map (
            O => \N__21204\,
            I => \N__21200\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__21203\,
            I => \N__21197\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__21200\,
            I => \N__21194\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21191\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__21194\,
            I => \IAC_CS\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__21191\,
            I => \IAC_CS\
        );

    \I__2239\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21183\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__21183\,
            I => n14_adj_1612
        );

    \I__2237\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21175\
        );

    \I__2236\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21172\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__21178\,
            I => \N__21169\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__21175\,
            I => \N__21166\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__21172\,
            I => \N__21163\
        );

    \I__2232\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21160\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__21166\,
            I => \N__21157\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__21163\,
            I => \N__21152\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__21160\,
            I => \N__21152\
        );

    \I__2228\ : Span4Mux_v
    port map (
            O => \N__21157\,
            I => \N__21147\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__21152\,
            I => \N__21144\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21141\
        );

    \I__2225\ : InMux
    port map (
            O => \N__21150\,
            I => \N__21138\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__21147\,
            I => \buf_cfgRTD_1\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__21144\,
            I => \buf_cfgRTD_1\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__21141\,
            I => \buf_cfgRTD_1\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__21138\,
            I => \buf_cfgRTD_1\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__21129\,
            I => \n14_adj_1610_cascade_\
        );

    \I__2219\ : IoInMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__2217\ : Span4Mux_s2_h
    port map (
            O => \N__21120\,
            I => \N__21117\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__21117\,
            I => \N__21113\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__21116\,
            I => \N__21110\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__21113\,
            I => \N__21107\
        );

    \I__2213\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21104\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__21107\,
            I => \VAC_CS\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__21104\,
            I => \VAC_CS\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__2209\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21092\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__21095\,
            I => \N__21089\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__21092\,
            I => \N__21086\
        );

    \I__2206\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21082\
        );

    \I__2205\ : Sp12to4
    port map (
            O => \N__21086\,
            I => \N__21079\
        );

    \I__2204\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21076\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__21082\,
            I => cmd_rdadctmp_14
        );

    \I__2202\ : Odrv12
    port map (
            O => \N__21079\,
            I => cmd_rdadctmp_14
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__21076\,
            I => cmd_rdadctmp_14
        );

    \I__2200\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21065\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__21068\,
            I => \N__21062\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__21065\,
            I => \N__21059\
        );

    \I__2197\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21056\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__21059\,
            I => cmd_rdadctmp_2_adj_1448
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__21056\,
            I => cmd_rdadctmp_2_adj_1448
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__21051\,
            I => \N__21047\
        );

    \I__2193\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21042\
        );

    \I__2192\ : InMux
    port map (
            O => \N__21047\,
            I => \N__21042\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__21042\,
            I => cmd_rdadctmp_3_adj_1447
        );

    \I__2190\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21036\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__21033\,
            I => \N__21028\
        );

    \I__2187\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21025\
        );

    \I__2186\ : InMux
    port map (
            O => \N__21031\,
            I => \N__21022\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__21028\,
            I => read_buf_7
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__21025\,
            I => read_buf_7
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__21022\,
            I => read_buf_7
        );

    \I__2182\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21012\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__21012\,
            I => \N__21008\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__21011\,
            I => \N__21005\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__21008\,
            I => \N__21002\
        );

    \I__2178\ : InMux
    port map (
            O => \N__21005\,
            I => \N__20999\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__21002\,
            I => \buf_readRTD_10\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__20999\,
            I => \buf_readRTD_10\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20980\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20975\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20992\,
            I => \N__20975\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20968\
        );

    \I__2171\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20968\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20968\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20961\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20961\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20961\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20958\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20953\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20953\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__20980\,
            I => \N__20941\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20941\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__20968\,
            I => \N__20941\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__20961\,
            I => \N__20941\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__20958\,
            I => \N__20936\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20936\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20931\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20931\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20928\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__20941\,
            I => \N__20925\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__20936\,
            I => \N__20922\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20931\,
            I => n1_adj_1606
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__20928\,
            I => n1_adj_1606
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__20925\,
            I => n1_adj_1606
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__20922\,
            I => n1_adj_1606
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__20913\,
            I => \N__20908\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__20912\,
            I => \N__20905\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__20911\,
            I => \N__20900\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20888\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20905\,
            I => \N__20888\
        );

    \I__2143\ : InMux
    port map (
            O => \N__20904\,
            I => \N__20883\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20883\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20880\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20899\,
            I => \N__20871\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20871\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20871\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20871\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20864\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20864\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20864\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__20888\,
            I => \N__20855\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__20883\,
            I => \N__20855\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20852\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20871\,
            I => \N__20847\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20864\,
            I => \N__20847\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20842\
        );

    \I__2127\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20842\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20837\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20860\,
            I => \N__20837\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__20855\,
            I => \N__20834\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__20852\,
            I => \N__20829\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__20847\,
            I => \N__20829\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__20842\,
            I => n13293
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20837\,
            I => n13293
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__20834\,
            I => n13293
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__20829\,
            I => n13293
        );

    \I__2117\ : InMux
    port map (
            O => \N__20820\,
            I => \N__20817\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__20817\,
            I => \N__20812\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20807\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20815\,
            I => \N__20807\
        );

    \I__2113\ : Odrv12
    port map (
            O => \N__20812\,
            I => read_buf_10
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__20807\,
            I => read_buf_10
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \N__20797\
        );

    \I__2110\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20794\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20791\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20788\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__20794\,
            I => read_buf_11
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20791\,
            I => read_buf_11
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__20788\,
            I => read_buf_11
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__20781\,
            I => \N__20776\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20773\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20768\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20768\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20773\,
            I => read_buf_13
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__20768\,
            I => read_buf_13
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__20763\,
            I => \N__20759\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__20762\,
            I => \N__20756\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20753\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20750\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20753\,
            I => \buf_readRTD_13\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20750\,
            I => \buf_readRTD_13\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__20745\,
            I => \N__20741\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__20744\,
            I => \N__20737\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20734\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20729\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20737\,
            I => \N__20729\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__20734\,
            I => read_buf_9
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20729\,
            I => read_buf_9
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__20724\,
            I => \N__20721\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20717\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20714\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20717\,
            I => \buf_readRTD_9\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20714\,
            I => \buf_readRTD_9\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__20709\,
            I => \N__20705\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__20708\,
            I => \N__20702\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20690\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20690\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20690\
        );

    \I__2075\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20690\
        );

    \I__2074\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20687\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__20690\,
            I => \RTD.bit_cnt_0\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20687\,
            I => \RTD.bit_cnt_0\
        );

    \I__2071\ : CEMux
    port map (
            O => \N__20682\,
            I => \N__20679\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__20676\,
            I => \N__20673\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__20673\,
            I => \RTD.n11740\
        );

    \I__2067\ : SRMux
    port map (
            O => \N__20670\,
            I => \N__20667\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20667\,
            I => \N__20664\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__20664\,
            I => \CLK_DDS.n16894\
        );

    \I__2064\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20657\
        );

    \I__2063\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20654\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20657\,
            I => read_buf_15
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__20654\,
            I => read_buf_15
        );

    \I__2060\ : InMux
    port map (
            O => \N__20649\,
            I => \N__20645\
        );

    \I__2059\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20641\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__20645\,
            I => \N__20638\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20635\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__20641\,
            I => buf_adcdata_iac_6
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__20638\,
            I => buf_adcdata_iac_6
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__20635\,
            I => buf_adcdata_iac_6
        );

    \I__2053\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20625\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__20625\,
            I => n22_adj_1627
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__2050\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20610\
        );

    \I__2049\ : InMux
    port map (
            O => \N__20618\,
            I => \N__20610\
        );

    \I__2048\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20610\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__20610\,
            I => cmd_rdadctmp_12
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__20607\,
            I => \N__20603\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__20606\,
            I => \N__20600\
        );

    \I__2044\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20596\
        );

    \I__2043\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20591\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20591\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__20596\,
            I => cmd_rdadctmp_13
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__20591\,
            I => cmd_rdadctmp_13
        );

    \I__2039\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20582\
        );

    \I__2038\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20579\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__20582\,
            I => \N__20575\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20579\,
            I => \N__20571\
        );

    \I__2035\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20568\
        );

    \I__2034\ : Span4Mux_h
    port map (
            O => \N__20575\,
            I => \N__20565\
        );

    \I__2033\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20562\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__20571\,
            I => \RTD.n17799\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__20568\,
            I => \RTD.n17799\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__20565\,
            I => \RTD.n17799\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20562\,
            I => \RTD.n17799\
        );

    \I__2028\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20546\
        );

    \I__2027\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20546\
        );

    \I__2026\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20541\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__20546\,
            I => \N__20538\
        );

    \I__2024\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20535\
        );

    \I__2023\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20532\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__20541\,
            I => \N__20529\
        );

    \I__2021\ : Span4Mux_h
    port map (
            O => \N__20538\,
            I => \N__20524\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__20535\,
            I => \N__20524\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__20532\,
            I => \RTD.bit_cnt_3\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__20529\,
            I => \RTD.bit_cnt_3\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__20524\,
            I => \RTD.bit_cnt_3\
        );

    \I__2016\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20507\
        );

    \I__2015\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20507\
        );

    \I__2014\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20507\
        );

    \I__2013\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20504\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__20507\,
            I => \RTD.bit_cnt_1\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__20504\,
            I => \RTD.bit_cnt_1\
        );

    \I__2010\ : InMux
    port map (
            O => \N__20499\,
            I => \N__20492\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20492\
        );

    \I__2008\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20489\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__20492\,
            I => \RTD.bit_cnt_2\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__20489\,
            I => \RTD.bit_cnt_2\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20481\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20481\,
            I => \N__20478\
        );

    \I__2003\ : Span4Mux_h
    port map (
            O => \N__20478\,
            I => \N__20473\
        );

    \I__2002\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20468\
        );

    \I__2001\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20468\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__20473\,
            I => buf_adcdata_vac_5
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__20468\,
            I => buf_adcdata_vac_5
        );

    \I__1998\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20460\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__20460\,
            I => \N__20457\
        );

    \I__1996\ : Span4Mux_h
    port map (
            O => \N__20457\,
            I => \N__20452\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20447\
        );

    \I__1994\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20447\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__20452\,
            I => buf_adcdata_iac_5
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__20447\,
            I => buf_adcdata_iac_5
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__20442\,
            I => \n19_adj_1629_cascade_\
        );

    \I__1990\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20436\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__20433\,
            I => buf_data_iac_6
        );

    \I__1987\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20426\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20422\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__20426\,
            I => \N__20419\
        );

    \I__1984\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20416\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__20422\,
            I => buf_adcdata_vac_4
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__20419\,
            I => buf_adcdata_vac_4
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20416\,
            I => buf_adcdata_vac_4
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__20409\,
            I => \n19_adj_1632_cascade_\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__20403\,
            I => \N__20400\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__20400\,
            I => \N__20395\
        );

    \I__1976\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20390\
        );

    \I__1975\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20390\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__20395\,
            I => buf_adcdata_iac_4
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__20390\,
            I => buf_adcdata_iac_4
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__20385\,
            I => \N__20380\
        );

    \I__1971\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20377\
        );

    \I__1970\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20372\
        );

    \I__1969\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20372\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__20377\,
            I => read_buf_12
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__20372\,
            I => read_buf_12
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__20367\,
            I => \N__20363\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__20366\,
            I => \N__20359\
        );

    \I__1964\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20352\
        );

    \I__1963\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20352\
        );

    \I__1962\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20352\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__20352\,
            I => read_buf_14
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__20349\,
            I => \N__20346\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__20343\,
            I => \N__20340\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__20340\,
            I => \N__20337\
        );

    \I__1956\ : Sp12to4
    port map (
            O => \N__20337\,
            I => \N__20334\
        );

    \I__1955\ : Odrv12
    port map (
            O => \N__20334\,
            I => \VAC_MISO\
        );

    \I__1954\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20328\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20324\
        );

    \I__1952\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20321\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__20324\,
            I => cmd_rdadctmp_0_adj_1450
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__20321\,
            I => cmd_rdadctmp_0_adj_1450
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__20316\,
            I => \N__20312\
        );

    \I__1948\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20307\
        );

    \I__1947\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20307\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__20307\,
            I => cmd_rdadctmp_1_adj_1449
        );

    \I__1945\ : IoInMux
    port map (
            O => \N__20304\,
            I => \N__20301\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__1943\ : IoSpan4Mux
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__1942\ : Span4Mux_s3_v
    port map (
            O => \N__20295\,
            I => \N__20292\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__20289\,
            I => \DDS_CS1\
        );

    \I__1939\ : CEMux
    port map (
            O => \N__20286\,
            I => \N__20283\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__20283\,
            I => \N__20280\
        );

    \I__1937\ : Span4Mux_v
    port map (
            O => \N__20280\,
            I => \N__20277\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__20277\,
            I => \CLK_DDS.n9_adj_1394\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20270\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20267\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20262\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20267\,
            I => \N__20262\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__20262\,
            I => \N__20258\
        );

    \I__1930\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20255\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__20258\,
            I => read_buf_0
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__20255\,
            I => read_buf_0
        );

    \I__1927\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20246\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__20249\,
            I => \N__20242\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20246\,
            I => \N__20239\
        );

    \I__1924\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20234\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20234\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__20239\,
            I => read_buf_1
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__20234\,
            I => read_buf_1
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__20229\,
            I => \N__20224\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20221\
        );

    \I__1918\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20218\
        );

    \I__1917\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20215\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__20221\,
            I => read_buf_5
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__20218\,
            I => read_buf_5
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20215\,
            I => read_buf_5
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__20208\,
            I => \N__20203\
        );

    \I__1912\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20200\
        );

    \I__1911\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20195\
        );

    \I__1910\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20195\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__20200\,
            I => read_buf_6
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__20195\,
            I => read_buf_6
        );

    \I__1907\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20187\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__20187\,
            I => \RTD.cfg_tmp_1\
        );

    \I__1905\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__20181\,
            I => \RTD.cfg_tmp_2\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20175\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__20175\,
            I => \RTD.cfg_tmp_3\
        );

    \I__1901\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20169\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__20169\,
            I => \RTD.cfg_tmp_4\
        );

    \I__1899\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20163\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__20163\,
            I => \RTD.cfg_tmp_5\
        );

    \I__1897\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20157\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__20157\,
            I => \RTD.cfg_tmp_6\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__20154\,
            I => \N__20151\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__20148\,
            I => \N__20145\
        );

    \I__1892\ : Span4Mux_v
    port map (
            O => \N__20145\,
            I => \N__20141\
        );

    \I__1891\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20138\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__20141\,
            I => \RTD.cfg_tmp_7\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__20138\,
            I => \RTD.cfg_tmp_7\
        );

    \I__1888\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20130\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__20130\,
            I => \RTD.cfg_tmp_0\
        );

    \I__1886\ : CEMux
    port map (
            O => \N__20127\,
            I => \N__20124\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__1884\ : Odrv12
    port map (
            O => \N__20121\,
            I => \RTD.n11704\
        );

    \I__1883\ : SRMux
    port map (
            O => \N__20118\,
            I => \N__20115\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__20115\,
            I => \N__20112\
        );

    \I__1881\ : Odrv12
    port map (
            O => \N__20112\,
            I => \RTD.n14999\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20106\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__20106\,
            I => \N__20102\
        );

    \I__1878\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20099\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__20102\,
            I => \N__20096\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__20099\,
            I => \N__20093\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__20096\,
            I => \N__20089\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__20093\,
            I => \N__20086\
        );

    \I__1873\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20083\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__20089\,
            I => read_buf_4
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__20086\,
            I => read_buf_4
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__20083\,
            I => read_buf_4
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__20076\,
            I => \N__20073\
        );

    \I__1868\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20069\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__20072\,
            I => \N__20065\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__20069\,
            I => \N__20062\
        );

    \I__1865\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20057\
        );

    \I__1864\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20057\
        );

    \I__1863\ : Span4Mux_h
    port map (
            O => \N__20062\,
            I => \N__20051\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__20057\,
            I => \N__20051\
        );

    \I__1861\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20048\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__20051\,
            I => \RTD.mode\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__20048\,
            I => \RTD.mode\
        );

    \I__1858\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20038\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__20042\,
            I => \N__20035\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__20041\,
            I => \N__20032\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__20038\,
            I => \N__20029\
        );

    \I__1854\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20026\
        );

    \I__1853\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20023\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__20029\,
            I => \N__20018\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__20026\,
            I => \N__20018\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__20015\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__20018\,
            I => \N__20012\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__20015\,
            I => \N__20009\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__20012\,
            I => \N__20006\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__20009\,
            I => \N__20003\
        );

    \I__1845\ : Sp12to4
    port map (
            O => \N__20006\,
            I => \N__19998\
        );

    \I__1844\ : Sp12to4
    port map (
            O => \N__20003\,
            I => \N__19998\
        );

    \I__1843\ : Odrv12
    port map (
            O => \N__19998\,
            I => \RTD_DRDY\
        );

    \I__1842\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19992\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__19992\,
            I => \N__19986\
        );

    \I__1840\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19983\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19976\
        );

    \I__1838\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19976\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__19986\,
            I => \N__19971\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19983\,
            I => \N__19971\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19966\
        );

    \I__1834\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19966\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__19976\,
            I => \RTD.adress_7_N_1339_7\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__19971\,
            I => \RTD.adress_7_N_1339_7\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__19966\,
            I => \RTD.adress_7_N_1339_7\
        );

    \I__1830\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19956\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__19956\,
            I => \N__19953\
        );

    \I__1828\ : Odrv12
    port map (
            O => \N__19953\,
            I => \RTD.n16638\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__19950\,
            I => \RTD.n16638_cascade_\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__19947\,
            I => \N__19944\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__1823\ : Span4Mux_h
    port map (
            O => \N__19938\,
            I => \N__19934\
        );

    \I__1822\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19931\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__19934\,
            I => \RTD.n20787\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__19931\,
            I => \RTD.n20787\
        );

    \I__1819\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__19923\,
            I => \RTD.n17835\
        );

    \I__1817\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19917\,
            I => \RTD.n7\
        );

    \I__1815\ : CEMux
    port map (
            O => \N__19914\,
            I => \N__19911\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19908\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__19908\,
            I => \N__19904\
        );

    \I__1812\ : CEMux
    port map (
            O => \N__19907\,
            I => \N__19901\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__19904\,
            I => \RTD.n11726\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__19901\,
            I => \RTD.n11726\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19893\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__19893\,
            I => \RTD.n19787\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__19890\,
            I => \RTD.n14_cascade_\
        );

    \I__1806\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19884\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__19884\,
            I => \N__19881\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__19881\,
            I => \N__19877\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19874\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__19877\,
            I => \RTD.n20832\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__19874\,
            I => \RTD.n20832\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__19869\,
            I => \RTD.n11704_cascade_\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__19866\,
            I => \N__19863\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19857\
        );

    \I__1797\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19857\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__19857\,
            I => adress_4
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__19854\,
            I => \RTD.n21362_cascade_\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19847\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19844\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19839\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__19844\,
            I => \N__19836\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19833\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19830\
        );

    \I__1788\ : Span4Mux_h
    port map (
            O => \N__19839\,
            I => \N__19827\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__19836\,
            I => \RTD.n1\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__19833\,
            I => \RTD.n1\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__19830\,
            I => \RTD.n1\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__19827\,
            I => \RTD.n1\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__19818\,
            I => \N__19813\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__19817\,
            I => \N__19809\
        );

    \I__1781\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19805\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19796\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19796\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19809\,
            I => \N__19796\
        );

    \I__1777\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19796\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__19805\,
            I => n14479
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__19796\,
            I => n14479
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19784\
        );

    \I__1772\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19781\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__19784\,
            I => adress_2
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__19781\,
            I => adress_2
        );

    \I__1769\ : CEMux
    port map (
            O => \N__19776\,
            I => \N__19773\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__1767\ : Span4Mux_h
    port map (
            O => \N__19770\,
            I => \N__19762\
        );

    \I__1766\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19759\
        );

    \I__1765\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19750\
        );

    \I__1764\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19750\
        );

    \I__1763\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19750\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19750\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__19762\,
            I => n13165
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__19759\,
            I => n13165
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19750\,
            I => n13165
        );

    \I__1758\ : InMux
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19740\,
            I => \N__19736\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19733\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__19736\,
            I => adress_3
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__19733\,
            I => adress_3
        );

    \I__1753\ : CEMux
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__19725\,
            I => \N__19722\
        );

    \I__1751\ : Odrv12
    port map (
            O => \N__19722\,
            I => \RTD.n11687\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19713\
        );

    \I__1749\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19713\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__19713\,
            I => adress_5
        );

    \I__1747\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19706\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19703\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19698\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19698\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__19698\,
            I => adress_6
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__19695\,
            I => \RTD.n19_cascade_\
        );

    \I__1741\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19689\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__19689\,
            I => \N__19686\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__19686\,
            I => \N__19683\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__19683\,
            I => adress_0
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__19680\,
            I => \n13165_cascade_\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19673\
        );

    \I__1735\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19670\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__19673\,
            I => adress_1
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__19670\,
            I => adress_1
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__19665\,
            I => \n14479_cascade_\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__19662\,
            I => \n1_adj_1606_cascade_\
        );

    \I__1730\ : SRMux
    port map (
            O => \N__19659\,
            I => \N__19655\
        );

    \I__1729\ : SRMux
    port map (
            O => \N__19658\,
            I => \N__19652\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__19655\,
            I => \N__19649\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__19652\,
            I => \N__19646\
        );

    \I__1726\ : Span4Mux_h
    port map (
            O => \N__19649\,
            I => \N__19643\
        );

    \I__1725\ : Span4Mux_v
    port map (
            O => \N__19646\,
            I => \N__19640\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__19643\,
            I => \RTD.n20160\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__19640\,
            I => \RTD.n20160\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19635\,
            I => \N__19631\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__19634\,
            I => \N__19627\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__19631\,
            I => \N__19624\
        );

    \I__1719\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19619\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19619\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__19624\,
            I => read_buf_3
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__19619\,
            I => read_buf_3
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__19614\,
            I => \N__19609\
        );

    \I__1714\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19606\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19601\
        );

    \I__1712\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19601\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__19606\,
            I => read_buf_2
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__19601\,
            I => read_buf_2
        );

    \I__1709\ : IoInMux
    port map (
            O => \N__19596\,
            I => \N__19593\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__19593\,
            I => \N__19590\
        );

    \I__1707\ : Span4Mux_s2_v
    port map (
            O => \N__19590\,
            I => \N__19587\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__19587\,
            I => \N__19584\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__19584\,
            I => \DDS_MCLK1\
        );

    \I__1704\ : IoInMux
    port map (
            O => \N__19581\,
            I => \N__19578\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__19578\,
            I => \N__19575\
        );

    \I__1702\ : Span4Mux_s3_h
    port map (
            O => \N__19575\,
            I => \N__19572\
        );

    \I__1701\ : Sp12to4
    port map (
            O => \N__19572\,
            I => \N__19569\
        );

    \I__1700\ : Span12Mux_s10_v
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__1699\ : Odrv12
    port map (
            O => \N__19566\,
            I => \RTD_CS\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__19563\,
            I => \RTD.n4_cascade_\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19556\
        );

    \I__1696\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19553\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__19556\,
            I => \RTD.cfg_buf_7\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__19553\,
            I => \RTD.cfg_buf_7\
        );

    \I__1693\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19544\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19541\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__19544\,
            I => cfg_buf_1
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__19541\,
            I => cfg_buf_1
        );

    \I__1689\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__19530\,
            I => \RTD.n12\
        );

    \I__1686\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__19524\,
            I => \RTD.n11\
        );

    \I__1684\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19518\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__19518\,
            I => \RTD.n11_adj_1403\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__19515\,
            I => \N__19512\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19509\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__19509\,
            I => \RTD.n32\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__19506\,
            I => \RTD.n32_cascade_\
        );

    \I__1678\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19500\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__19500\,
            I => \RTD.n21555\
        );

    \I__1676\ : InMux
    port map (
            O => \N__19497\,
            I => \N__19494\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__19494\,
            I => \RTD.n6\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__19491\,
            I => \N__19488\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19485\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19485\,
            I => \N__19482\
        );

    \I__1671\ : Span12Mux_s7_h
    port map (
            O => \N__19482\,
            I => \N__19479\
        );

    \I__1670\ : Span12Mux_v
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__1669\ : Odrv12
    port map (
            O => \N__19476\,
            I => \RTD_SDO\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__19473\,
            I => \N__19470\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19467\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__19467\,
            I => \N__19463\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19460\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__19463\,
            I => \RTD.cfg_buf_6\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__19460\,
            I => \RTD.cfg_buf_6\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__19455\,
            I => \N__19452\
        );

    \I__1661\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19448\
        );

    \I__1660\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19445\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__19448\,
            I => cfg_buf_0
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__19445\,
            I => cfg_buf_0
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__19440\,
            I => \RTD.n9_cascade_\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__19437\,
            I => \RTD.adress_7_N_1339_7_cascade_\
        );

    \I__1655\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19430\
        );

    \I__1654\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19427\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__19430\,
            I => \RTD.cfg_buf_5\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__19427\,
            I => \RTD.cfg_buf_5\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19418\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19415\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19418\,
            I => \RTD.cfg_buf_3\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__19415\,
            I => \RTD.cfg_buf_3\
        );

    \I__1647\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19407\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__19407\,
            I => \RTD.n11_adj_1405\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__19404\,
            I => \N__19401\
        );

    \I__1644\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19397\
        );

    \I__1643\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19394\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__19397\,
            I => \RTD.cfg_buf_4\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__19394\,
            I => \RTD.cfg_buf_4\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__19389\,
            I => \N__19386\
        );

    \I__1639\ : InMux
    port map (
            O => \N__19386\,
            I => \N__19382\
        );

    \I__1638\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19379\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__19382\,
            I => \RTD.cfg_buf_2\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__19379\,
            I => \RTD.cfg_buf_2\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19371\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__19371\,
            I => \RTD.n10\
        );

    \I__1633\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19364\
        );

    \I__1632\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19361\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__19364\,
            I => \RTD.adress_7\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__19361\,
            I => \RTD.adress_7\
        );

    \I__1629\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19353\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__19353\,
            I => \N__19350\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__19350\,
            I => \RTD.n7318\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__19347\,
            I => \RTD.n7318_cascade_\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__19344\,
            I => \RTD.n21_cascade_\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__19341\,
            I => \n13176_cascade_\
        );

    \I__1623\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19319\
        );

    \I__1622\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19319\
        );

    \I__1621\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19319\
        );

    \I__1620\ : InMux
    port map (
            O => \N__19335\,
            I => \N__19319\
        );

    \I__1619\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19319\
        );

    \I__1618\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19319\
        );

    \I__1617\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19316\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__19319\,
            I => n18755
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__19316\,
            I => n18755
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__19311\,
            I => \N__19306\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__19310\,
            I => \N__19303\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__19309\,
            I => \N__19298\
        );

    \I__1611\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19282\
        );

    \I__1610\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19282\
        );

    \I__1609\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19282\
        );

    \I__1608\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19282\
        );

    \I__1607\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19282\
        );

    \I__1606\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19282\
        );

    \I__1605\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19277\
        );

    \I__1604\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19277\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__19282\,
            I => n13176
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__19277\,
            I => n13176
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__19272\,
            I => \n18755_cascade_\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19266\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__19266\,
            I => \RTD.n16\
        );

    \I__1598\ : CEMux
    port map (
            O => \N__19263\,
            I => \N__19260\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__19260\,
            I => \N__19257\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__19257\,
            I => \RTD.n8\
        );

    \I__1595\ : IoInMux
    port map (
            O => \N__19254\,
            I => \N__19251\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__1593\ : Span4Mux_s0_h
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__1592\ : Sp12to4
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__1591\ : Span12Mux_v
    port map (
            O => \N__19242\,
            I => \N__19239\
        );

    \I__1590\ : Odrv12
    port map (
            O => \N__19239\,
            I => \RTD_SDI\
        );

    \I__1589\ : CEMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__1587\ : Span4Mux_h
    port map (
            O => \N__19230\,
            I => \N__19227\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__19227\,
            I => \RTD.n11718\
        );

    \I__1585\ : IoInMux
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__1583\ : IoSpan4Mux
    port map (
            O => \N__19218\,
            I => \N__19215\
        );

    \I__1582\ : IoSpan4Mux
    port map (
            O => \N__19215\,
            I => \N__19212\
        );

    \I__1581\ : Span4Mux_s2_h
    port map (
            O => \N__19212\,
            I => \N__19209\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__19209\,
            I => \RTD_SCLK\
        );

    \I__1579\ : IoInMux
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__1577\ : IoSpan4Mux
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__1576\ : IoSpan4Mux
    port map (
            O => \N__19197\,
            I => \N__19194\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__19194\,
            I => \ICE_SYSCLK\
        );

    \I__1574\ : IoInMux
    port map (
            O => \N__19191\,
            I => \N__19188\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__1572\ : IoSpan4Mux
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__1571\ : Span4Mux_s3_v
    port map (
            O => \N__19182\,
            I => \N__19179\
        );

    \I__1570\ : Sp12to4
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__1569\ : Span12Mux_h
    port map (
            O => \N__19176\,
            I => \N__19173\
        );

    \I__1568\ : Odrv12
    port map (
            O => \N__19173\,
            I => \ICE_GPMO_2\
        );

    \INVADC_VDC.genclk.t0on_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i8C_net\,
            I => \N__38755\
        );

    \INVADC_VDC.genclk.t0on_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i0C_net\,
            I => \N__38754\
        );

    \INVADC_VDC.genclk.div_state_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i0C_net\,
            I => \N__38753\
        );

    \INVADC_VDC.genclk.div_state_i1C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i1C_net\,
            I => \N__38749\
        );

    \INVADC_VDC.genclk.t0off_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i8C_net\,
            I => \N__38752\
        );

    \INVADC_VDC.genclk.t0off_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i0C_net\,
            I => \N__38750\
        );

    \INVdata_cntvec_i0_i8C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i8C_net\,
            I => \N__54400\
        );

    \INVdata_cntvec_i0_i0C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i0C_net\,
            I => \N__54388\
        );

    \INVcomm_spi.data_valid_85C\ : INV
    port map (
            O => \INVcomm_spi.data_valid_85C_net\,
            I => \N__54295\
        );

    \INVacadc_skipcnt_i0_i9C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i9C_net\,
            I => \N__54393\
        );

    \INVacadc_skipcnt_i0_i1C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i1C_net\,
            I => \N__54381\
        );

    \INVacadc_skipcnt_i0_i0C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i0C_net\,
            I => \N__54366\
        );

    \INVcomm_spi.imiso_83_12192_12193_setC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12192_12193_setC_net\,
            I => \N__52601\
        );

    \INVdds0_mclk_294C\ : INV
    port map (
            O => \INVdds0_mclk_294C_net\,
            I => \N__38745\
        );

    \INVcomm_spi.MISO_48_12186_12187_setC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12186_12187_setC_net\,
            I => \N__54271\
        );

    \INVcomm_spi.imiso_83_12192_12193_resetC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12192_12193_resetC_net\,
            I => \N__52502\
        );

    \INVdds0_mclkcnt_i7_3772__i0C\ : INV
    port map (
            O => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            I => \N__38739\
        );

    \INVeis_state_i2C\ : INV
    port map (
            O => \INVeis_state_i2C_net\,
            I => \N__54398\
        );

    \INVeis_end_299C\ : INV
    port map (
            O => \INVeis_end_299C_net\,
            I => \N__54359\
        );

    \INVdata_count_i0_i8C\ : INV
    port map (
            O => \INVdata_count_i0_i8C_net\,
            I => \N__54331\
        );

    \INVdata_count_i0_i0C\ : INV
    port map (
            O => \INVdata_count_i0_i0C_net\,
            I => \N__54318\
        );

    \INVcomm_spi.MISO_48_12186_12187_resetC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12186_12187_resetC_net\,
            I => \N__54269\
        );

    \INVeis_state_i0C\ : INV
    port map (
            O => \INVeis_state_i0C_net\,
            I => \N__54384\
        );

    \INVcomm_spi.bit_cnt_3767__i3C\ : INV
    port map (
            O => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            I => \N__52498\
        );

    \INVacadc_trig_300C\ : INV
    port map (
            O => \INVacadc_trig_300C_net\,
            I => \N__54412\
        );

    \INViac_raw_buf_vac_raw_buf_merged2WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            I => \N__54380\
        );

    \INViac_raw_buf_vac_raw_buf_merged7WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            I => \N__54438\
        );

    \INViac_raw_buf_vac_raw_buf_merged1WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            I => \N__54298\
        );

    \INViac_raw_buf_vac_raw_buf_merged6WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            I => \N__54436\
        );

    \INViac_raw_buf_vac_raw_buf_merged0WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            I => \N__54285\
        );

    \INViac_raw_buf_vac_raw_buf_merged5WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            I => \N__54434\
        );

    \INViac_raw_buf_vac_raw_buf_merged9WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            I => \N__54338\
        );

    \INViac_raw_buf_vac_raw_buf_merged4WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            I => \N__54426\
        );

    \INViac_raw_buf_vac_raw_buf_merged8WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            I => \N__54312\
        );

    \INViac_raw_buf_vac_raw_buf_merged10WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            I => \N__54326\
        );

    \INViac_raw_buf_vac_raw_buf_merged3WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            I => \N__54407\
        );

    \INViac_raw_buf_vac_raw_buf_merged11WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            I => \N__54352\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19757,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19765,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \n19610_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19618,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19602,
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19593,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19641,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19632,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_19_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19716\,
            carryinitout => \bfn_19_8_0_\
        );

    \IN_MUX_bfv_22_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_7_0_\
        );

    \IN_MUX_bfv_22_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19731\,
            carryinitout => \bfn_22_8_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_4_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19705\,
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19670\,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19678\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19686\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19694\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RTD.SCLK_51_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010110100110"
        )
    port map (
            in0 => \N__26783\,
            in1 => \N__26596\,
            in2 => \N__26277\,
            in3 => \N__26415\,
            lcout => \RTD_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30472\,
            ce => \N__19263\,
            sr => \_gnd_net_\
        );

    \RTD.i19375_4_lut_4_lut_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111011111"
        )
    port map (
            in0 => \N__26782\,
            in1 => \N__26559\,
            in2 => \N__26441\,
            in3 => \N__26272\,
            lcout => \RTD.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i7_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__19338\,
            in1 => \N__31301\,
            in2 => \N__19311\,
            in3 => \N__19560\,
            lcout => \RTD.cfg_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_40_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010000000"
        )
    port map (
            in0 => \N__26533\,
            in1 => \N__26735\,
            in2 => \N__26391\,
            in3 => \N__26271\,
            lcout => n11714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i4_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__22782\,
            in1 => \N__19302\,
            in2 => \N__19404\,
            in3 => \N__19336\,
            lcout => \RTD.cfg_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i5_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__19337\,
            in1 => \N__21821\,
            in2 => \N__19310\,
            in3 => \N__19434\,
            lcout => \RTD.cfg_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i2_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__21882\,
            in1 => \N__19301\,
            in2 => \N__19389\,
            in3 => \N__19335\,
            lcout => \RTD.cfg_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i1_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__19334\,
            in1 => \N__21180\,
            in2 => \N__19309\,
            in3 => \N__19548\,
            lcout => cfg_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i0_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__23261\,
            in1 => \N__19297\,
            in2 => \N__19455\,
            in3 => \N__19333\,
            lcout => cfg_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30518\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.MOSI_59_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__19367\,
            in1 => \N__26778\,
            in2 => \N__20154\,
            in3 => \N__26273\,
            lcout => \RTD_SDI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30508\,
            ce => \N__19236\,
            sr => \N__19659\
        );

    \RTD.i27_4_lut_4_lut_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000110"
        )
    port map (
            in0 => \N__26724\,
            in1 => \N__26541\,
            in2 => \N__26421\,
            in3 => \N__26252\,
            lcout => \RTD.n11718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i2_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19613\,
            in1 => \N__21639\,
            in2 => \N__46664\,
            in3 => \N__26836\,
            lcout => \buf_readRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i6_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__31378\,
            in1 => \N__19296\,
            in2 => \N__19473\,
            in3 => \N__19332\,
            lcout => \RTD.cfg_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_34_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__26268\,
            in1 => \N__19356\,
            in2 => \N__20041\,
            in3 => \N__19981\,
            lcout => OPEN,
            ltout => \RTD.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_35_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101000"
        )
    port map (
            in0 => \N__20056\,
            in1 => \N__26426\,
            in2 => \N__19344\,
            in3 => \N__26750\,
            lcout => \RTD.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i22_4_lut_4_lut_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010110000000"
        )
    port map (
            in0 => \N__26749\,
            in1 => \N__19851\,
            in2 => \N__26443\,
            in3 => \N__19880\,
            lcout => n13176,
            ltout => \n13176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_3_lut_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26425\,
            in2 => \N__19341\,
            in3 => \N__26269\,
            lcout => n18755,
            ltout => \n18755_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i3_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__24692\,
            in1 => \N__19295\,
            in2 => \N__19272\,
            in3 => \N__19422\,
            lcout => \RTD.cfg_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.mode_53_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__19982\,
            in1 => \N__26270\,
            in2 => \N__19947\,
            in3 => \N__19269\,
            lcout => \RTD.mode\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i7_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__19990\,
            in1 => \N__19710\,
            in2 => \N__26585\,
            in3 => \N__26260\,
            lcout => \RTD.adress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30517\,
            ce => \N__19776\,
            sr => \N__19658\
        );

    \RTD.i1_4_lut_adj_37_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__31386\,
            in1 => \N__19466\,
            in2 => \N__23262\,
            in3 => \N__19451\,
            lcout => OPEN,
            ltout => \RTD.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i7_4_lut_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19536\,
            in1 => \N__19374\,
            in2 => \N__19440\,
            in3 => \N__19410\,
            lcout => \RTD.adress_7_N_1339_7\,
            ltout => \RTD.adress_7_N_1339_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__26258\,
            in1 => \_gnd_net_\,
            in2 => \N__19437\,
            in3 => \N__26544\,
            lcout => \RTD.n20832\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i3_4_lut_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__19433\,
            in1 => \N__24691\,
            in2 => \N__21822\,
            in3 => \N__19421\,
            lcout => \RTD.n11_adj_1405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_4_lut_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__22777\,
            in1 => \N__19400\,
            in2 => \N__21881\,
            in3 => \N__19385\,
            lcout => \RTD.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i0_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111001111"
        )
    port map (
            in0 => \N__19989\,
            in1 => \N__19368\,
            in2 => \N__26584\,
            in3 => \N__26259\,
            lcout => adress_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30517\,
            ce => \N__19776\,
            sr => \N__19658\
        );

    \RTD.adc_state_i2_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__26764\,
            in1 => \N__19850\,
            in2 => \N__26427\,
            in3 => \N__19503\,
            lcout => adc_state_2_adj_1481,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30525\,
            ce => \N__19914\,
            sr => \_gnd_net_\
        );

    \RTD.i4903_2_lut_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26762\,
            in2 => \_gnd_net_\,
            in3 => \N__26534\,
            lcout => \RTD.n7318\,
            ltout => \RTD.n7318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i1_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__26381\,
            in1 => \N__19521\,
            in2 => \N__19347\,
            in3 => \N__26263\,
            lcout => \RTD.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30525\,
            ce => \N__19914\,
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26535\,
            in2 => \_gnd_net_\,
            in3 => \N__20585\,
            lcout => OPEN,
            ltout => \RTD.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i3_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111000000"
        )
    port map (
            in0 => \N__26763\,
            in1 => \N__19527\,
            in2 => \N__19563\,
            in3 => \N__26385\,
            lcout => \RTD.adc_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30525\,
            ce => \N__19914\,
            sr => \_gnd_net_\
        );

    \RTD.i4_4_lut_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__21179\,
            in1 => \N__19559\,
            in2 => \N__31300\,
            in3 => \N__19547\,
            lcout => \RTD.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i22_4_lut_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000110"
        )
    port map (
            in0 => \N__26261\,
            in1 => \N__26726\,
            in2 => \N__20072\,
            in3 => \N__20553\,
            lcout => \RTD.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i24_4_lut_4_lut_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100110"
        )
    port map (
            in0 => \N__26725\,
            in1 => \N__26543\,
            in2 => \N__19515\,
            in3 => \N__26262\,
            lcout => \RTD.n11_adj_1403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_23_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20552\,
            in2 => \_gnd_net_\,
            in3 => \N__20586\,
            lcout => \RTD.n32\,
            ltout => \RTD.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19313_4_lut_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__26380\,
            in1 => \N__19497\,
            in2 => \N__19506\,
            in3 => \N__20068\,
            lcout => \RTD.n21555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_31_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__26251\,
            in1 => \N__26542\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RTD.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i0_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__20261\,
            in1 => \N__20950\,
            in2 => \N__19491\,
            in3 => \N__20861\,
            lcout => read_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_adj_26_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__26419\,
            in1 => \_gnd_net_\,
            in2 => \N__26837\,
            in3 => \N__26267\,
            lcout => n1_adj_1606,
            ltout => \n1_adj_1606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i4_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__20860\,
            in1 => \N__20092\,
            in2 => \N__19662\,
            in3 => \N__19635\,
            lcout => read_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_39_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010010001"
        )
    port map (
            in0 => \N__26784\,
            in1 => \N__26580\,
            in2 => \N__26442\,
            in3 => \N__26266\,
            lcout => n13293,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__26265\,
            in1 => \N__26785\,
            in2 => \N__26597\,
            in3 => \N__26420\,
            lcout => \RTD.n20160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i3_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19612\,
            in1 => \N__20952\,
            in2 => \N__19634\,
            in3 => \N__20863\,
            lcout => read_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i3_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19630\,
            in1 => \N__21670\,
            in2 => \N__50141\,
            in3 => \N__26815\,
            lcout => \buf_readRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i2_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20250\,
            in1 => \N__20951\,
            in2 => \N__19614\,
            in3 => \N__20862\,
            lcout => read_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_main.i19883_1_lut_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38765\,
            lcout => \DDS_MCLK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.CS_52_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001101011111"
        )
    port map (
            in0 => \N__26593\,
            in1 => \N__19959\,
            in2 => \N__26447\,
            in3 => \N__26257\,
            lcout => \RTD_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30416\,
            ce => \N__19728\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34750\,
            in2 => \_gnd_net_\,
            in3 => \N__34529\,
            lcout => dds_state_2_adj_1452,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19332_3_lut_3_lut_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010011001"
        )
    port map (
            in0 => \N__26435\,
            in1 => \N__26829\,
            in2 => \_gnd_net_\,
            in3 => \N__26592\,
            lcout => \RTD.n11687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i4_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33680\,
            in1 => \N__33388\,
            in2 => \N__28296\,
            in3 => \N__20429\,
            lcout => buf_adcdata_vac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i5_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19718\,
            in1 => \N__19812\,
            in2 => \N__19866\,
            in3 => \N__19767\,
            lcout => adress_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i6_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19768\,
            in1 => \N__19719\,
            in2 => \N__19818\,
            in3 => \N__19709\,
            lcout => adress_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i34_4_lut_4_lut_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110011101"
        )
    port map (
            in0 => \N__26594\,
            in1 => \N__26253\,
            in2 => \N__20042\,
            in3 => \N__19991\,
            lcout => OPEN,
            ltout => \RTD.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i35_4_lut_4_lut_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__26830\,
            in1 => \N__26436\,
            in2 => \N__19695\,
            in3 => \N__19843\,
            lcout => n13165,
            ltout => \n13165_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i1_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__19692\,
            in1 => \N__19676\,
            in2 => \N__19680\,
            in3 => \N__19808\,
            lcout => adress_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12067_2_lut_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26437\,
            in2 => \_gnd_net_\,
            in3 => \N__26595\,
            lcout => n14479,
            ltout => \n14479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i2_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__19677\,
            in1 => \N__19787\,
            in2 => \N__19665\,
            in3 => \N__19765\,
            lcout => adress_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i4_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19766\,
            in1 => \N__19743\,
            in2 => \N__19817\,
            in3 => \N__19862\,
            lcout => adress_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_2_lut_3_lut_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__26389\,
            in1 => \N__26760\,
            in2 => \_gnd_net_\,
            in3 => \N__26561\,
            lcout => \RTD.n20787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19242_3_lut_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__26565\,
            in1 => \N__20551\,
            in2 => \_gnd_net_\,
            in3 => \N__20578\,
            lcout => OPEN,
            ltout => \RTD.n21362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__26766\,
            in1 => \N__19842\,
            in2 => \N__19854\,
            in3 => \N__26189\,
            lcout => \RTD.n17835\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i7_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__21684\,
            in1 => \N__21039\,
            in2 => \N__50177\,
            in3 => \N__26767\,
            lcout => \buf_readRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4933_2_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26560\,
            in2 => \_gnd_net_\,
            in3 => \N__26187\,
            lcout => \RTD.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19410_4_lut_4_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101101111000"
        )
    port map (
            in0 => \N__26188\,
            in1 => \N__26765\,
            in2 => \N__26591\,
            in3 => \N__26390\,
            lcout => \RTD.n11740\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i4_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20109\,
            in1 => \N__21683\,
            in2 => \N__22700\,
            in3 => \N__26761\,
            lcout => \buf_readRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i3_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__19816\,
            in1 => \N__19739\,
            in2 => \N__19791\,
            in3 => \N__19769\,
            lcout => adress_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000101010101"
        )
    port map (
            in0 => \N__26234\,
            in1 => \N__26820\,
            in2 => \N__20076\,
            in3 => \N__19896\,
            lcout => \RTD.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_38_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__20043\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19995\,
            lcout => \RTD.n16638\,
            ltout => \RTD.n16638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_adj_24_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__26233\,
            in1 => \_gnd_net_\,
            in2 => \N__19950\,
            in3 => \N__19937\,
            lcout => \RTD.n11726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i0_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__19926\,
            in1 => \N__26434\,
            in2 => \_gnd_net_\,
            in3 => \N__19920\,
            lcout => \RTD.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30468\,
            ce => \N__19907\,
            sr => \_gnd_net_\
        );

    \RTD.i17182_3_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__20545\,
            in1 => \N__26590\,
            in2 => \_gnd_net_\,
            in3 => \N__20574\,
            lcout => \RTD.n19787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i31_3_lut_3_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26589\,
            in1 => \N__26431\,
            in2 => \_gnd_net_\,
            in3 => \N__26232\,
            lcout => OPEN,
            ltout => \RTD.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i30_4_lut_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__26432\,
            in1 => \N__26819\,
            in2 => \N__19890\,
            in3 => \N__19887\,
            lcout => \RTD.n11704\,
            ltout => \RTD.n11704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12586_2_lut_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19869\,
            in3 => \N__26433\,
            lcout => \RTD.n14999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_tmp_i1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__26199\,
            in1 => \N__20133\,
            in2 => \N__21178\,
            in3 => \N__26847\,
            lcout => \RTD.cfg_tmp_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.cfg_tmp_i2_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__26843\,
            in1 => \N__20190\,
            in2 => \N__21877\,
            in3 => \N__26206\,
            lcout => \RTD.cfg_tmp_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.cfg_tmp_i3_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__26200\,
            in1 => \N__20184\,
            in2 => \N__24696\,
            in3 => \N__26848\,
            lcout => \RTD.cfg_tmp_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.cfg_tmp_i4_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__26844\,
            in1 => \N__26204\,
            in2 => \N__22781\,
            in3 => \N__20178\,
            lcout => \RTD.cfg_tmp_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.cfg_tmp_i5_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__26201\,
            in1 => \N__26846\,
            in2 => \N__21811\,
            in3 => \N__20172\,
            lcout => \RTD.cfg_tmp_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.cfg_tmp_i6_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__26845\,
            in1 => \N__26205\,
            in2 => \N__31385\,
            in3 => \N__20166\,
            lcout => \RTD.cfg_tmp_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.cfg_tmp_i7_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__26202\,
            in1 => \N__20160\,
            in2 => \N__31302\,
            in3 => \N__26849\,
            lcout => \RTD.cfg_tmp_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.cfg_tmp_i0_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__26842\,
            in1 => \N__26203\,
            in2 => \N__23257\,
            in3 => \N__20144\,
            lcout => \RTD.cfg_tmp_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30492\,
            ce => \N__20127\,
            sr => \N__20118\
        );

    \RTD.read_buf_i5_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__20893\,
            in1 => \N__20105\,
            in2 => \N__20229\,
            in3 => \N__20985\,
            lcout => read_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26838\,
            in1 => \N__20273\,
            in2 => \N__43439\,
            in3 => \N__21701\,
            lcout => \buf_readRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i1_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__21703\,
            in1 => \N__20245\,
            in2 => \N__37193\,
            in3 => \N__26840\,
            lcout => \buf_readRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20274\,
            in1 => \N__20984\,
            in2 => \N__20249\,
            in3 => \N__20895\,
            lcout => read_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i6_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__21704\,
            in1 => \N__20207\,
            in2 => \N__46304\,
            in3 => \N__26841\,
            lcout => \buf_readRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i12_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__21702\,
            in1 => \N__20383\,
            in2 => \N__22727\,
            in3 => \N__26839\,
            lcout => \buf_readRTD_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i12_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20801\,
            in1 => \N__20983\,
            in2 => \N__20385\,
            in3 => \N__20894\,
            lcout => read_buf_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i14_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__20896\,
            in1 => \N__20779\,
            in2 => \N__20366\,
            in3 => \N__20992\,
            lcout => read_buf_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i7_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__20206\,
            in1 => \N__20988\,
            in2 => \N__20911\,
            in3 => \N__21031\,
            lcout => read_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20227\,
            in1 => \N__21710\,
            in2 => \N__51194\,
            in3 => \N__26833\,
            lcout => \buf_readRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i6_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20228\,
            in1 => \N__20987\,
            in2 => \N__20208\,
            in3 => \N__20899\,
            lcout => read_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i15_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__20897\,
            in1 => \N__20660\,
            in2 => \N__20367\,
            in3 => \N__20993\,
            lcout => read_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i13_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20384\,
            in1 => \N__20986\,
            in2 => \N__20781\,
            in3 => \N__20898\,
            lcout => read_buf_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i14_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20362\,
            in1 => \N__21709\,
            in2 => \N__31403\,
            in3 => \N__26832\,
            lcout => \buf_readRTD_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__20327\,
            in1 => \N__33387\,
            in2 => \N__20349\,
            in3 => \N__31619\,
            lcout => cmd_rdadctmp_0_adj_1450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19764_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21793\,
            in1 => \N__55158\,
            in2 => \N__20763\,
            in3 => \N__57738\,
            lcout => n22405,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i5_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56554\,
            in1 => \N__41891\,
            in2 => \N__43600\,
            in3 => \N__23047\,
            lcout => \AMPV_POW\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i1_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20331\,
            in1 => \N__33389\,
            in2 => \N__20316\,
            in3 => \N__31562\,
            lcout => cmd_rdadctmp_1_adj_1449,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i2_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20315\,
            in1 => \N__33390\,
            in2 => \N__21068\,
            in3 => \N__31563\,
            lcout => cmd_rdadctmp_2_adj_1448,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.CS_28_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__34796\,
            in1 => \N__34567\,
            in2 => \_gnd_net_\,
            in3 => \N__34459\,
            lcout => \DDS_CS1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54275\,
            ce => \N__20286\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.i23_4_lut_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110110011001"
        )
    port map (
            in0 => \N__34710\,
            in1 => \N__34548\,
            in2 => \N__44073\,
            in3 => \N__34458\,
            lcout => \CLK_DDS.n9_adj_1394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i5_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35797\,
            in1 => \N__35625\,
            in2 => \N__20607\,
            in3 => \N__20456\,
            lcout => buf_adcdata_iac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i5_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__20477\,
            in1 => \N__33681\,
            in2 => \N__21612\,
            in3 => \N__33475\,
            lcout => buf_adcdata_vac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i19_3_lut_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21264\,
            in1 => \N__20476\,
            in2 => \_gnd_net_\,
            in3 => \N__57815\,
            lcout => OPEN,
            ltout => \n19_adj_1629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i22_3_lut_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20455\,
            in2 => \N__20442\,
            in3 => \N__53797\,
            lcout => n22_adj_1630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i6_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35624\,
            in1 => \N__35798\,
            in2 => \N__21095\,
            in3 => \N__20648\,
            lcout => buf_adcdata_iac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i30_3_lut_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20439\,
            in1 => \N__20628\,
            in2 => \_gnd_net_\,
            in3 => \N__54765\,
            lcout => n30_adj_1628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i19_3_lut_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24081\,
            in1 => \N__20425\,
            in2 => \_gnd_net_\,
            in3 => \N__57816\,
            lcout => OPEN,
            ltout => \n19_adj_1632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i22_3_lut_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20398\,
            in2 => \N__20409\,
            in3 => \N__53799\,
            lcout => n22_adj_1633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i4_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35802\,
            in1 => \N__35632\,
            in2 => \N__20622\,
            in3 => \N__20399\,
            lcout => buf_adcdata_iac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i22_3_lut_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53798\,
            in1 => \N__20644\,
            in2 => \_gnd_net_\,
            in3 => \N__21357\,
            lcout => n22_adj_1627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i12_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__20617\,
            in1 => \N__28103\,
            in2 => \N__28398\,
            in3 => \N__35633\,
            lcout => cmd_rdadctmp_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i13_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__35631\,
            in1 => \N__20618\,
            in2 => \N__28123\,
            in3 => \N__20599\,
            lcout => cmd_rdadctmp_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i14_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__21085\,
            in1 => \N__28104\,
            in2 => \N__20606\,
            in3 => \N__35634\,
            lcout => cmd_rdadctmp_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i10_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20820\,
            in1 => \N__21708\,
            in2 => \N__21011\,
            in3 => \N__26831\,
            lcout => \buf_readRTD_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i1_3_lut_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__34711\,
            in1 => \N__34536\,
            in2 => \_gnd_net_\,
            in3 => \N__34425\,
            lcout => \CLK_DDS.n16894\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20699\,
            in1 => \N__20514\,
            in2 => \_gnd_net_\,
            in3 => \N__20497\,
            lcout => \RTD.n17799\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.bit_cnt_3771__i3_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__20517\,
            in1 => \N__20544\,
            in2 => \N__20709\,
            in3 => \N__20499\,
            lcout => \RTD.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30449\,
            ce => \N__20682\,
            sr => \N__26088\
        );

    \RTD.bit_cnt_3771__i1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20701\,
            in2 => \_gnd_net_\,
            in3 => \N__20515\,
            lcout => \RTD.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30449\,
            ce => \N__20682\,
            sr => \N__26088\
        );

    \RTD.bit_cnt_3771__i2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20516\,
            in1 => \_gnd_net_\,
            in2 => \N__20708\,
            in3 => \N__20498\,
            lcout => \RTD.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30449\,
            ce => \N__20682\,
            sr => \N__26088\
        );

    \RTD.bit_cnt_3771__i0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20700\,
            lcout => \RTD.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30449\,
            ce => \N__20682\,
            sr => \N__26088\
        );

    \i15340_2_lut_3_lut_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__40120\,
            in1 => \N__51726\,
            in2 => \_gnd_net_\,
            in3 => \N__55516\,
            lcout => n14_adj_1580,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15341_2_lut_3_lut_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__55517\,
            in1 => \N__50319\,
            in2 => \_gnd_net_\,
            in3 => \N__51727\,
            lcout => n14_adj_1551,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i3_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__24777\,
            in1 => \N__21422\,
            in2 => \N__21402\,
            in3 => \N__21441\,
            lcout => bit_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54340\,
            ce => \N__34751\,
            sr => \N__20670\
        );

    \CLK_DDS.bit_cnt_i2_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21421\,
            in1 => \N__21398\,
            in2 => \_gnd_net_\,
            in3 => \N__24776\,
            lcout => bit_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54340\,
            ce => \N__34751\,
            sr => \N__20670\
        );

    \CLK_DDS.bit_cnt_i1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21420\,
            lcout => bit_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54340\,
            ce => \N__34751\,
            sr => \N__20670\
        );

    \ADC_VAC.cmd_rdadctmp_i27_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33450\,
            in1 => \N__24485\,
            in2 => \N__22637\,
            in3 => \N__31592\,
            lcout => cmd_rdadctmp_27_adj_1423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i11_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20816\,
            in1 => \N__20990\,
            in2 => \N__20802\,
            in3 => \N__20904\,
            lcout => read_buf_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i15_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20661\,
            in1 => \N__21712\,
            in2 => \N__31319\,
            in3 => \N__26835\,
            lcout => \buf_readRTD_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i8_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__21733\,
            in1 => \N__20991\,
            in2 => \N__20913\,
            in3 => \N__21032\,
            lcout => read_buf_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i9_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__20903\,
            in1 => \N__21734\,
            in2 => \N__20744\,
            in3 => \N__20994\,
            lcout => read_buf_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18472_3_lut_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21015\,
            in1 => \N__21843\,
            in2 => \_gnd_net_\,
            in3 => \N__57784\,
            lcout => n21082,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i10_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__20815\,
            in1 => \N__20989\,
            in2 => \N__20912\,
            in3 => \N__20740\,
            lcout => read_buf_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i11_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20800\,
            in1 => \N__21711\,
            in2 => \N__24629\,
            in3 => \N__26834\,
            lcout => \buf_readRTD_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i13_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26851\,
            in1 => \N__20780\,
            in2 => \N__20762\,
            in3 => \N__21719\,
            lcout => \buf_readRTD_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21150\,
            in1 => \N__55159\,
            in2 => \N__20724\,
            in3 => \N__57740\,
            lcout => n22441,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i9_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__21720\,
            in1 => \N__20720\,
            in2 => \N__20745\,
            in3 => \N__26852\,
            lcout => \buf_readRTD_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i23_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35535\,
            in1 => \N__22891\,
            in2 => \N__25127\,
            in3 => \N__28046\,
            lcout => cmd_rdadctmp_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i22_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__28045\,
            in1 => \N__35240\,
            in2 => \N__22895\,
            in3 => \N__35538\,
            lcout => cmd_rdadctmp_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i10_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35742\,
            in1 => \N__35537\,
            in2 => \N__23346\,
            in3 => \N__46633\,
            lcout => buf_adcdata_iac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i1_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56555\,
            in1 => \N__27300\,
            in2 => \N__40161\,
            in3 => \N__21151\,
            lcout => \buf_cfgRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35536\,
            in1 => \N__21299\,
            in2 => \N__22655\,
            in3 => \N__28047\,
            lcout => cmd_rdadctmp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__31560\,
            in1 => \N__21050\,
            in2 => \N__21245\,
            in3 => \N__33273\,
            lcout => cmd_rdadctmp_4_adj_1446,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i16_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__35558\,
            in1 => \N__23143\,
            in2 => \N__28065\,
            in3 => \N__22946\,
            lcout => cmd_rdadctmp_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_192_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__33264\,
            in1 => \N__30707\,
            in2 => \N__21116\,
            in3 => \N__27438\,
            lcout => OPEN,
            ltout => \n14_adj_1610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.CS_37_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__23099\,
            in1 => \N__21231\,
            in2 => \N__21129\,
            in3 => \N__33266\,
            lcout => \VAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i15_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22945\,
            in1 => \N__28005\,
            in2 => \N__21099\,
            in3 => \N__35559\,
            lcout => cmd_rdadctmp_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i3_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21069\,
            in1 => \N__33265\,
            in2 => \N__21051\,
            in3 => \N__31559\,
            lcout => cmd_rdadctmp_3_adj_1447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__31561\,
            in1 => \N__21926\,
            in2 => \N__21246\,
            in3 => \N__33274\,
            lcout => cmd_rdadctmp_5_adj_1445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i2_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__33221\,
            in1 => \N__30702\,
            in2 => \_gnd_net_\,
            in3 => \N__27431\,
            lcout => \DTRIG_N_918_adj_1451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54419\,
            ce => \N__21219\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i1_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__33220\,
            in1 => \N__30701\,
            in2 => \_gnd_net_\,
            in3 => \N__27432\,
            lcout => adc_state_1_adj_1417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54419\,
            ce => \N__21219\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_203_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30700\,
            in2 => \_gnd_net_\,
            in3 => \N__27430\,
            lcout => n20864,
            ltout => \n20864_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_3_lut_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23100\,
            in2 => \N__21225\,
            in3 => \N__33219\,
            lcout => n12653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i30_4_lut_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000101"
        )
    port map (
            in0 => \N__30706\,
            in1 => \N__23101\,
            in2 => \N__27448\,
            in3 => \N__25404\,
            lcout => OPEN,
            ltout => \ADC_VAC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19365_2_lut_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21222\,
            in3 => \N__33259\,
            lcout => \ADC_VAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.CS_37_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__35408\,
            in1 => \N__21186\,
            in2 => \N__25936\,
            in3 => \N__21351\,
            lcout => \IAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_195_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001110"
        )
    port map (
            in0 => \N__29883\,
            in1 => \N__29973\,
            in2 => \N__21203\,
            in3 => \N__35407\,
            lcout => n14_adj_1612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_199_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29959\,
            in2 => \_gnd_net_\,
            in3 => \N__29882\,
            lcout => n20867,
            ltout => \n20867_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_3_lut_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25929\,
            in2 => \N__21345\,
            in3 => \N__35406\,
            lcout => n12498,
            ltout => \n12498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__35409\,
            in1 => \N__21342\,
            in2 => \N__21324\,
            in3 => \N__21320\,
            lcout => cmd_rdadctmp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i1_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35410\,
            in1 => \N__21321\,
            in2 => \N__21312\,
            in3 => \N__28035\,
            lcout => cmd_rdadctmp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i2_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__28034\,
            in1 => \N__35411\,
            in2 => \N__21300\,
            in3 => \N__21311\,
            lcout => cmd_rdadctmp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_I_0_1_lut_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40898\,
            lcout => \AC_ADC_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i5_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25701\,
            in1 => \N__48843\,
            in2 => \N__21263\,
            in3 => \N__22236\,
            lcout => buf_adcdata_vdc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34547\,
            in2 => \_gnd_net_\,
            in3 => \N__34453\,
            lcout => dds_state_1_adj_1453,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54287\,
            ce => \N__21377\,
            sr => \N__34772\
        );

    \ADC_VDC.cmd_rdadctmp_i11_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__23988\,
            in1 => \N__22267\,
            in2 => \N__23888\,
            in3 => \N__48586\,
            lcout => cmd_rdadctmp_11_adj_1468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__48583\,
            in1 => \N__24038\,
            in2 => \N__23630\,
            in3 => \N__23861\,
            lcout => cmd_rdadctmp_14_adj_1465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i22_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__22321\,
            in1 => \N__26047\,
            in2 => \N__23891\,
            in3 => \N__48589\,
            lcout => cmd_rdadctmp_22_adj_1457,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__48585\,
            in1 => \N__22322\,
            in2 => \N__22350\,
            in3 => \N__23869\,
            lcout => cmd_rdadctmp_21_adj_1458,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__22345\,
            in1 => \N__23739\,
            in2 => \N__23890\,
            in3 => \N__48588\,
            lcout => cmd_rdadctmp_20_adj_1459,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i12_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48582\,
            in1 => \N__23860\,
            in2 => \N__22272\,
            in3 => \N__24061\,
            lcout => cmd_rdadctmp_12_adj_1467,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i18_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__22376\,
            in1 => \N__23761\,
            in2 => \N__23889\,
            in3 => \N__48587\,
            lcout => cmd_rdadctmp_18_adj_1461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i17_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__48584\,
            in1 => \N__22375\,
            in2 => \N__23925\,
            in3 => \N__23862\,
            lcout => cmd_rdadctmp_17_adj_1462,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i19_3_lut_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24339\,
            in1 => \N__21538\,
            in2 => \_gnd_net_\,
            in3 => \N__57747\,
            lcout => n19_adj_1626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i13_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__33490\,
            in1 => \N__21592\,
            in2 => \N__28292\,
            in3 => \N__31683\,
            lcout => cmd_rdadctmp_13_adj_1437,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i7_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33650\,
            in1 => \N__33492\,
            in2 => \N__21498\,
            in3 => \N__24292\,
            lcout => buf_adcdata_vac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i16_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33491\,
            in1 => \N__21494\,
            in2 => \N__21473\,
            in3 => \N__31684\,
            lcout => cmd_rdadctmp_16_adj_1434,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i17_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__31685\,
            in1 => \N__21469\,
            in2 => \N__31711\,
            in3 => \N__33493\,
            lcout => cmd_rdadctmp_17_adj_1433,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i8_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33489\,
            in1 => \N__33651\,
            in2 => \N__21474\,
            in3 => \N__21568\,
            lcout => buf_adcdata_vac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i30_3_lut_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21456\,
            in1 => \N__21447\,
            in2 => \_gnd_net_\,
            in3 => \N__54753\,
            lcout => n30_adj_1634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010100000101"
        )
    port map (
            in0 => \N__34437\,
            in1 => \N__21384\,
            in2 => \N__34752\,
            in3 => \N__21429\,
            lcout => dds_state_0_adj_1454,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54315\,
            ce => \N__21378\,
            sr => \_gnd_net_\
        );

    \SecClk_292_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39168\,
            in2 => \_gnd_net_\,
            in3 => \N__31137\,
            lcout => \TEST_LED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18974_2_lut_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24774\,
            in2 => \_gnd_net_\,
            in3 => \N__21440\,
            lcout => n21456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i3_3_lut_4_lut_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34595\,
            in1 => \N__34423\,
            in2 => \N__21423\,
            in3 => \N__21397\,
            lcout => n8_adj_1602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i19392_4_lut_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__34594\,
            in1 => \N__34424\,
            in2 => \N__44069\,
            in3 => \N__34706\,
            lcout => \CLK_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i19_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33620\,
            in1 => \N__33307\,
            in2 => \N__25282\,
            in3 => \N__22636\,
            lcout => buf_adcdata_vac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i29_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__31670\,
            in1 => \N__22585\,
            in2 => \N__33375\,
            in3 => \N__22613\,
            lcout => cmd_rdadctmp_29_adj_1421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i14_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21508\,
            in1 => \N__33308\,
            in2 => \N__21611\,
            in3 => \N__31668\,
            lcout => cmd_rdadctmp_14_adj_1436,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_0_i19_3_lut_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23679\,
            in1 => \N__21569\,
            in2 => \_gnd_net_\,
            in3 => \N__57572\,
            lcout => n19_adj_1486,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i6_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33306\,
            in1 => \N__33621\,
            in2 => \N__21542\,
            in3 => \N__21512\,
            lcout => buf_adcdata_vac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21485\,
            in1 => \N__33309\,
            in2 => \N__21513\,
            in3 => \N__31669\,
            lcout => cmd_rdadctmp_15_adj_1435,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i16_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33603\,
            in1 => \N__33486\,
            in2 => \N__21764\,
            in3 => \N__22679\,
            lcout => buf_adcdata_vac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i23_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__24903\,
            in1 => \N__33487\,
            in2 => \N__24509\,
            in3 => \N__31628\,
            lcout => cmd_rdadctmp_23_adj_1427,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i24_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__24505\,
            in1 => \N__33488\,
            in2 => \N__21763\,
            in3 => \N__31629\,
            lcout => cmd_rdadctmp_24_adj_1426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i30_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__22596\,
            in1 => \N__33374\,
            in2 => \N__22857\,
            in3 => \N__31660\,
            lcout => cmd_rdadctmp_30_adj_1420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56558\,
            in1 => \N__27298\,
            in2 => \N__44229\,
            in3 => \N__24671\,
            lcout => \buf_cfgRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i2_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__27297\,
            in1 => \N__56559\,
            in2 => \N__44793\,
            in3 => \N__21844\,
            lcout => \buf_cfgRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56557\,
            in1 => \N__27299\,
            in2 => \N__43605\,
            in3 => \N__21789\,
            lcout => \buf_cfgRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i20_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__31994\,
            in1 => \N__28063\,
            in2 => \N__25036\,
            in3 => \N__35520\,
            lcout => cmd_rdadctmp_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i25_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21765\,
            in1 => \N__33373\,
            in2 => \N__24416\,
            in3 => \N__31659\,
            lcout => cmd_rdadctmp_25_adj_1425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19694_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23025\,
            in1 => \N__54748\,
            in2 => \N__35196\,
            in3 => \N__53780\,
            lcout => OPEN,
            ltout => \n22321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22321_bdd_4_lut_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__54749\,
            in1 => \N__22788\,
            in2 => \N__21741\,
            in3 => \N__22908\,
            lcout => n22324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i8_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__21738\,
            in1 => \N__21718\,
            in2 => \N__23277\,
            in3 => \N__26856\,
            lcout => \buf_readRTD_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i7_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__31565\,
            in1 => \N__21914\,
            in2 => \N__22562\,
            in3 => \N__33272\,
            lcout => cmd_rdadctmp_7_adj_1443,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i15_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__35719\,
            in1 => \N__35459\,
            in2 => \N__52177\,
            in3 => \N__25126\,
            lcout => buf_adcdata_iac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.SCLK_35_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000101100000"
        )
    port map (
            in0 => \N__27439\,
            in1 => \N__33267\,
            in2 => \N__21947\,
            in3 => \N__30708\,
            lcout => \VAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i6_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21930\,
            in1 => \N__33268\,
            in2 => \N__21915\,
            in3 => \N__31564\,
            lcout => cmd_rdadctmp_6_adj_1444,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i0_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__30713\,
            in1 => \N__27440\,
            in2 => \N__33343\,
            in3 => \N__21903\,
            lcout => adc_state_0_adj_1418,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54410\,
            ce => \N__21894\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29993\,
            in2 => \_gnd_net_\,
            in3 => \N__29902\,
            lcout => n20858,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i12393_2_lut_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__29994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25877\,
            lcout => \ADC_IAC.n14806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19093_4_lut_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__33260\,
            in1 => \N__27434\,
            in2 => \N__25323\,
            in3 => \N__25446\,
            lcout => \ADC_VAC.n21312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__33245\,
            in1 => \N__23102\,
            in2 => \N__30720\,
            in3 => \N__25403\,
            lcout => OPEN,
            ltout => \ADC_VAC.n20958_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_adj_4_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21897\,
            in3 => \N__27433\,
            lcout => \ADC_VAC.n20959\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i17_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__23156\,
            in1 => \N__27975\,
            in2 => \N__23122\,
            in3 => \N__35405\,
            lcout => cmd_rdadctmp_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54428\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i2_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35403\,
            in2 => \N__29995\,
            in3 => \N__29901\,
            lcout => \DTRIG_N_918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54432\,
            ce => \N__23505\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i1_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__29900\,
            in1 => \N__29974\,
            in2 => \_gnd_net_\,
            in3 => \N__35404\,
            lcout => adc_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54432\,
            ce => \N__23505\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_3_lut_4_lut_4_lut_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110000000"
        )
    port map (
            in0 => \N__47385\,
            in1 => \N__48847\,
            in2 => \N__48357\,
            in3 => \N__48568\,
            lcout => \ADC_VDC.n13034\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7_4_lut_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22014\,
            in1 => \N__21971\,
            in2 => \N__22035\,
            in3 => \N__22101\,
            lcout => OPEN,
            ltout => \ADC_VDC.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i11_3_lut_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23448\,
            in2 => \N__21996\,
            in3 => \N__23391\,
            lcout => \ADC_VDC.n18563\,
            ltout => \ADC_VDC.n18563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16137_3_lut_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48350\,
            in2 => \N__21993\,
            in3 => \N__47384\,
            lcout => \ADC_VDC.n18566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19290_3_lut_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__24226\,
            in1 => \_gnd_net_\,
            in2 => \N__48871\,
            in3 => \N__21990\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i34_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__48354\,
            in1 => \N__22386\,
            in2 => \N__21984\,
            in3 => \N__48569\,
            lcout => cmd_rdadcbuf_34,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53325\,
            ce => \N__21981\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.avg_cnt_i0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21972\,
            in2 => \_gnd_net_\,
            in3 => \N__21960\,
            lcout => \ADC_VDC.avg_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \ADC_VDC.n19698\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23417\,
            in2 => \_gnd_net_\,
            in3 => \N__22056\,
            lcout => \ADC_VDC.avg_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19698\,
            carryout => \ADC_VDC.n19699\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i2_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23430\,
            in2 => \_gnd_net_\,
            in3 => \N__22053\,
            lcout => \ADC_VDC.avg_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19699\,
            carryout => \ADC_VDC.n19700\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i3_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23474\,
            in2 => \_gnd_net_\,
            in3 => \N__22050\,
            lcout => \ADC_VDC.avg_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19700\,
            carryout => \ADC_VDC.n19701\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i4_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23499\,
            in2 => \_gnd_net_\,
            in3 => \N__22047\,
            lcout => \ADC_VDC.avg_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19701\,
            carryout => \ADC_VDC.n19702\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i5_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23460\,
            in2 => \_gnd_net_\,
            in3 => \N__22044\,
            lcout => \ADC_VDC.avg_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19702\,
            carryout => \ADC_VDC.n19703\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i6_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23403\,
            in2 => \_gnd_net_\,
            in3 => \N__22041\,
            lcout => \ADC_VDC.avg_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19703\,
            carryout => \ADC_VDC.n19704\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i7_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23487\,
            in2 => \_gnd_net_\,
            in3 => \N__22038\,
            lcout => \ADC_VDC.avg_cnt_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19704\,
            carryout => \ADC_VDC.n19705\,
            clk => \N__53319\,
            ce => \N__22506\,
            sr => \N__22443\
        );

    \ADC_VDC.avg_cnt_i8_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22031\,
            in2 => \_gnd_net_\,
            in3 => \N__22017\,
            lcout => \ADC_VDC.avg_cnt_8\,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \ADC_VDC.n19706\,
            clk => \N__53320\,
            ce => \N__22514\,
            sr => \N__22452\
        );

    \ADC_VDC.avg_cnt_i9_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22013\,
            in2 => \_gnd_net_\,
            in3 => \N__21999\,
            lcout => \ADC_VDC.avg_cnt_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19706\,
            carryout => \ADC_VDC.n19707\,
            clk => \N__53320\,
            ce => \N__22514\,
            sr => \N__22452\
        );

    \ADC_VDC.avg_cnt_i10_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22100\,
            in2 => \_gnd_net_\,
            in3 => \N__22086\,
            lcout => \ADC_VDC.avg_cnt_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19707\,
            carryout => \ADC_VDC.n19708\,
            clk => \N__53320\,
            ce => \N__22514\,
            sr => \N__22452\
        );

    \ADC_VDC.avg_cnt_i11_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23442\,
            in2 => \_gnd_net_\,
            in3 => \N__22083\,
            lcout => \ADC_VDC.avg_cnt_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53320\,
            ce => \N__22514\,
            sr => \N__22452\
        );

    \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__22184\,
            in1 => \N__23599\,
            in2 => \N__23838\,
            in3 => \N__48562\,
            lcout => cmd_rdadctmp_3_adj_1476,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010101000"
        )
    port map (
            in0 => \N__48556\,
            in1 => \N__48347\,
            in2 => \N__48869\,
            in3 => \N__47364\,
            lcout => \ADC_VDC.n13010\,
            ltout => \ADC_VDC.n13010_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i12541_2_lut_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22080\,
            in3 => \N__48557\,
            lcout => \ADC_VDC.n14915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__48558\,
            in1 => \N__48348\,
            in2 => \N__48870\,
            in3 => \N__47365\,
            lcout => n12871,
            ltout => \n12871_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i2_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__22183\,
            in1 => \N__22211\,
            in2 => \N__22077\,
            in3 => \N__48561\,
            lcout => cmd_rdadctmp_2_adj_1477,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__22073\,
            in1 => \N__22210\,
            in2 => \N__23837\,
            in3 => \N__48560\,
            lcout => cmd_rdadctmp_1_adj_1478,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48559\,
            in1 => \N__23800\,
            in2 => \N__47426\,
            in3 => \N__22072\,
            lcout => cmd_rdadctmp_0_adj_1479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22218\,
            in2 => \N__22074\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.cmd_rdadcbuf_0\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \ADC_VDC.n19663\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22194\,
            in2 => \N__22212\,
            in3 => \N__22188\,
            lcout => \ADC_VDC.cmd_rdadcbuf_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19663\,
            carryout => \ADC_VDC.n19664\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22167\,
            in2 => \N__22185\,
            in3 => \N__22161\,
            lcout => \ADC_VDC.cmd_rdadcbuf_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19664\,
            carryout => \ADC_VDC.n19665\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22158\,
            in2 => \N__23601\,
            in3 => \N__22152\,
            lcout => \ADC_VDC.cmd_rdadcbuf_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19665\,
            carryout => \ADC_VDC.n19666\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22149\,
            in2 => \N__23580\,
            in3 => \N__22143\,
            lcout => \ADC_VDC.cmd_rdadcbuf_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19666\,
            carryout => \ADC_VDC.n19667\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22140\,
            in2 => \N__24160\,
            in3 => \N__22134\,
            lcout => \ADC_VDC.cmd_rdadcbuf_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19667\,
            carryout => \ADC_VDC.n19668\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22131\,
            in2 => \N__24131\,
            in3 => \N__22125\,
            lcout => \ADC_VDC.cmd_rdadcbuf_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19668\,
            carryout => \ADC_VDC.n19669\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24106\,
            in2 => \N__22122\,
            in3 => \N__22113\,
            lcout => \ADC_VDC.cmd_rdadcbuf_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19669\,
            carryout => \ADC_VDC.n19670\,
            clk => \N__53256\,
            ce => \N__22521\,
            sr => \N__22453\
        );

    \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22110\,
            in2 => \N__23559\,
            in3 => \N__22104\,
            lcout => \ADC_VDC.cmd_rdadcbuf_8\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \ADC_VDC.n19671\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22290\,
            in2 => \N__24011\,
            in3 => \N__22284\,
            lcout => \ADC_VDC.cmd_rdadcbuf_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19671\,
            carryout => \ADC_VDC.n19672\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22281\,
            in2 => \N__23987\,
            in3 => \N__22275\,
            lcout => \ADC_VDC.cmd_rdadcbuf_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19672\,
            carryout => \ADC_VDC.n19673\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25784\,
            in2 => \N__22271\,
            in3 => \N__22251\,
            lcout => cmd_rdadcbuf_11,
            ltout => OPEN,
            carryin => \ADC_VDC.n19673\,
            carryout => \ADC_VDC.n19674\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23654\,
            in2 => \N__24062\,
            in3 => \N__22248\,
            lcout => cmd_rdadcbuf_12,
            ltout => OPEN,
            carryin => \ADC_VDC.n19674\,
            carryout => \ADC_VDC.n19675\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23642\,
            in2 => \N__24037\,
            in3 => \N__22245\,
            lcout => cmd_rdadcbuf_13,
            ltout => OPEN,
            carryin => \ADC_VDC.n19675\,
            carryout => \ADC_VDC.n19676\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23960\,
            in2 => \N__23626\,
            in3 => \N__22242\,
            lcout => cmd_rdadcbuf_14,
            ltout => OPEN,
            carryin => \ADC_VDC.n19676\,
            carryout => \ADC_VDC.n19677\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24092\,
            in2 => \N__23948\,
            in3 => \N__22239\,
            lcout => cmd_rdadcbuf_15,
            ltout => OPEN,
            carryin => \ADC_VDC.n19677\,
            carryout => \ADC_VDC.n19678\,
            clk => \N__53278\,
            ce => \N__22513\,
            sr => \N__22447\
        );

    \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22232\,
            in2 => \N__23917\,
            in3 => \N__22221\,
            lcout => cmd_rdadcbuf_16,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \ADC_VDC.n19679\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24350\,
            in2 => \N__22377\,
            in3 => \N__22359\,
            lcout => cmd_rdadcbuf_17,
            ltout => OPEN,
            carryin => \ADC_VDC.n19679\,
            carryout => \ADC_VDC.n19680\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23537\,
            in2 => \N__23762\,
            in3 => \N__22356\,
            lcout => cmd_rdadcbuf_18,
            ltout => OPEN,
            carryin => \ADC_VDC.n19680\,
            carryout => \ADC_VDC.n19681\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23690\,
            in2 => \N__23734\,
            in3 => \N__22353\,
            lcout => cmd_rdadcbuf_19,
            ltout => OPEN,
            carryin => \ADC_VDC.n19681\,
            carryout => \ADC_VDC.n19682\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24269\,
            in2 => \N__22349\,
            in3 => \N__22326\,
            lcout => cmd_rdadcbuf_20,
            ltout => OPEN,
            carryin => \ADC_VDC.n19682\,
            carryout => \ADC_VDC.n19683\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25763\,
            in2 => \N__22323\,
            in3 => \N__22305\,
            lcout => cmd_rdadcbuf_21,
            ltout => OPEN,
            carryin => \ADC_VDC.n19683\,
            carryout => \ADC_VDC.n19684\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24257\,
            in2 => \N__26051\,
            in3 => \N__22302\,
            lcout => cmd_rdadcbuf_22,
            ltout => OPEN,
            carryin => \ADC_VDC.n19684\,
            carryout => \ADC_VDC.n19685\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24320\,
            in2 => \N__26028\,
            in3 => \N__22299\,
            lcout => cmd_rdadcbuf_23,
            ltout => OPEN,
            carryin => \ADC_VDC.n19685\,
            carryout => \ADC_VDC.n19686\,
            clk => \N__53276\,
            ce => \N__22519\,
            sr => \N__22454\
        );

    \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24365\,
            in2 => \_gnd_net_\,
            in3 => \N__22296\,
            lcout => cmd_rdadcbuf_24,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \ADC_VDC.n19687\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23705\,
            in2 => \_gnd_net_\,
            in3 => \N__22293\,
            lcout => cmd_rdadcbuf_25,
            ltout => OPEN,
            carryin => \ADC_VDC.n19687\,
            carryout => \ADC_VDC.n19688\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26066\,
            in2 => \_gnd_net_\,
            in3 => \N__22545\,
            lcout => cmd_rdadcbuf_26,
            ltout => OPEN,
            carryin => \ADC_VDC.n19688\,
            carryout => \ADC_VDC.n19689\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23378\,
            in2 => \_gnd_net_\,
            in3 => \N__22542\,
            lcout => cmd_rdadcbuf_27,
            ltout => OPEN,
            carryin => \ADC_VDC.n19689\,
            carryout => \ADC_VDC.n19690\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24245\,
            in2 => \_gnd_net_\,
            in3 => \N__22539\,
            lcout => cmd_rdadcbuf_28,
            ltout => OPEN,
            carryin => \ADC_VDC.n19690\,
            carryout => \ADC_VDC.n19691\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24527\,
            in2 => \_gnd_net_\,
            in3 => \N__22536\,
            lcout => cmd_rdadcbuf_29,
            ltout => OPEN,
            carryin => \ADC_VDC.n19691\,
            carryout => \ADC_VDC.n19692\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24539\,
            in2 => \_gnd_net_\,
            in3 => \N__22533\,
            lcout => cmd_rdadcbuf_30,
            ltout => OPEN,
            carryin => \ADC_VDC.n19692\,
            carryout => \ADC_VDC.n19693\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24551\,
            in2 => \_gnd_net_\,
            in3 => \N__22530\,
            lcout => cmd_rdadcbuf_31,
            ltout => OPEN,
            carryin => \ADC_VDC.n19693\,
            carryout => \ADC_VDC.n19694\,
            clk => \N__53301\,
            ce => \N__22515\,
            sr => \N__22451\
        );

    \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24584\,
            in2 => \_gnd_net_\,
            in3 => \N__22527\,
            lcout => cmd_rdadcbuf_32,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \ADC_VDC.n19695\,
            clk => \N__53318\,
            ce => \N__22520\,
            sr => \N__22455\
        );

    \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25802\,
            in2 => \_gnd_net_\,
            in3 => \N__22524\,
            lcout => cmd_rdadcbuf_33,
            ltout => OPEN,
            carryin => \ADC_VDC.n19695\,
            carryout => \ADC_VDC.n19696\,
            clk => \N__53318\,
            ce => \N__22520\,
            sr => \N__22455\
        );

    \ADC_VDC.add_23_36_lut_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24233\,
            in2 => \_gnd_net_\,
            in3 => \N__22389\,
            lcout => \ADC_VDC.cmd_rdadcbuf_35_N_1138_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18591_3_lut_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23367\,
            in1 => \N__22675\,
            in2 => \_gnd_net_\,
            in3 => \N__57777\,
            lcout => n21201,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i4_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__22659\,
            in1 => \N__28097\,
            in2 => \N__35585\,
            in3 => \N__27026\,
            lcout => cmd_rdadctmp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i23_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33377\,
            in1 => \N__33649\,
            in2 => \N__22875\,
            in3 => \N__24184\,
            lcout => buf_adcdata_vac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i20_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33647\,
            in1 => \N__33379\,
            in2 => \N__25091\,
            in3 => \N__22612\,
            lcout => buf_adcdata_vac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i28_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__33378\,
            in1 => \N__31671\,
            in2 => \N__22614\,
            in3 => \N__22638\,
            lcout => cmd_rdadctmp_28_adj_1422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i21_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33376\,
            in1 => \N__33648\,
            in2 => \N__22595\,
            in3 => \N__22810\,
            lcout => buf_adcdata_vac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i8_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__31672\,
            in1 => \N__26923\,
            in2 => \N__22569\,
            in3 => \N__33380\,
            lcout => cmd_rdadctmp_8_adj_1442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i22_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__31656\,
            in1 => \N__24946\,
            in2 => \N__24902\,
            in3 => \N__33484\,
            lcout => cmd_rdadctmp_22_adj_1428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i10_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33481\,
            in1 => \N__33734\,
            in2 => \N__28333\,
            in3 => \N__31655\,
            lcout => cmd_rdadctmp_10_adj_1440,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i31_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__31658\,
            in1 => \N__22855\,
            in2 => \N__22874\,
            in3 => \N__33485\,
            lcout => cmd_rdadctmp_31_adj_1419,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i26_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33482\,
            in1 => \N__24412\,
            in2 => \N__24484\,
            in3 => \N__31657\,
            lcout => cmd_rdadctmp_26_adj_1424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i22_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33657\,
            in1 => \N__33483\,
            in2 => \N__40429\,
            in3 => \N__22856\,
            lcout => buf_adcdata_vac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22405_bdd_4_lut_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__22839\,
            in1 => \N__55170\,
            in2 => \N__22820\,
            in3 => \N__24573\,
            lcout => n21097,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i4_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56560\,
            in1 => \N__27296\,
            in2 => \N__41496\,
            in3 => \N__22756\,
            lcout => \buf_cfgRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18529_3_lut_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57794\,
            in1 => \N__27344\,
            in2 => \_gnd_net_\,
            in3 => \N__27629\,
            lcout => n21139,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19778_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__22755\,
            in1 => \N__57795\,
            in2 => \N__22737\,
            in3 => \N__55171\,
            lcout => n22417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i7_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56561\,
            in1 => \N__44862\,
            in2 => \N__45362\,
            in3 => \N__31885\,
            lcout => \VAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19621_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__24591\,
            in1 => \N__55172\,
            in2 => \N__22710\,
            in3 => \N__53786\,
            lcout => n22231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i25_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35551\,
            in1 => \N__27373\,
            in2 => \N__31964\,
            in3 => \N__28112\,
            lcout => cmd_rdadctmp_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_5_i23_3_lut_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23051\,
            in1 => \N__57786\,
            in2 => \_gnd_net_\,
            in3 => \N__32247\,
            lcout => OPEN,
            ltout => \n23_adj_1540_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18513_4_lut_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__57787\,
            in1 => \N__55162\,
            in2 => \N__23028\,
            in3 => \N__33948\,
            lcout => n21123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \EIS_SYNCCLK_I_0_1_lut_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23019\,
            lcout => \IAC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i7_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35531\,
            in1 => \N__35756\,
            in2 => \N__22956\,
            in3 => \N__24826\,
            lcout => buf_adcdata_iac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19704_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011010000"
        )
    port map (
            in0 => \N__53779\,
            in1 => \N__22932\,
            in2 => \N__55213\,
            in3 => \N__27060\,
            lcout => n22327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19689_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__22920\,
            in1 => \N__55164\,
            in2 => \N__23196\,
            in3 => \N__53778\,
            lcout => n22291,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19729_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__55163\,
            in1 => \N__23173\,
            in2 => \N__24997\,
            in3 => \N__57788\,
            lcout => OPEN,
            ltout => \n22315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22315_bdd_4_lut_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__41630\,
            in1 => \N__27180\,
            in2 => \N__22911\,
            in3 => \N__55165\,
            lcout => n22318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i14_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35806\,
            in1 => \N__35458\,
            in2 => \N__22902\,
            in3 => \N__47032\,
            lcout => buf_adcdata_iac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_80_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30721\,
            in2 => \_gnd_net_\,
            in3 => \N__27449\,
            lcout => n20853,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i6_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__27295\,
            in1 => \N__45357\,
            in2 => \N__56568\,
            in3 => \N__31352\,
            lcout => \buf_cfgRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i0_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__23220\,
            in1 => \N__56563\,
            in2 => \N__43829\,
            in3 => \N__27294\,
            lcout => \buf_cfgRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18592_3_lut_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57785\,
            in1 => \N__23276\,
            in2 => \_gnd_net_\,
            in3 => \N__23219\,
            lcout => n21202,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i6_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56562\,
            in1 => \N__44861\,
            in2 => \N__43601\,
            in3 => \N__23174\,
            lcout => \VAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i8_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__35492\,
            in1 => \N__35702\,
            in2 => \N__43504\,
            in3 => \N__23157\,
            lcout => buf_adcdata_iac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i9_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35701\,
            in1 => \N__35495\,
            in2 => \N__23127\,
            in3 => \N__37159\,
            lcout => buf_adcdata_iac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i18_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__35493\,
            in1 => \N__23123\,
            in2 => \N__28118\,
            in3 => \N__23338\,
            lcout => cmd_rdadctmp_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_adj_5_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000100"
        )
    port map (
            in0 => \N__33218\,
            in1 => \N__30709\,
            in2 => \N__23103\,
            in3 => \N__27441\,
            lcout => \ADC_VAC.n12594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i19_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35494\,
            in1 => \N__23339\,
            in2 => \N__31993\,
            in3 => \N__28091\,
            lcout => cmd_rdadctmp_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.SCLK_35_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111000000010"
        )
    port map (
            in0 => \N__30002\,
            in1 => \N__35496\,
            in2 => \N__29916\,
            in3 => \N__23306\,
            lcout => \IAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15343_2_lut_3_lut_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__47794\,
            in1 => \N__51994\,
            in2 => \_gnd_net_\,
            in3 => \N__55560\,
            lcout => n14_adj_1553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.bit_cnt_i0_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25422\,
            in2 => \_gnd_net_\,
            in3 => \N__23295\,
            lcout => \ADC_IAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \ADC_IAC.n19649\,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.bit_cnt_i1_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25571\,
            in2 => \_gnd_net_\,
            in3 => \N__23292\,
            lcout => \ADC_IAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19649\,
            carryout => \ADC_IAC.n19650\,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.bit_cnt_i2_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25623\,
            in2 => \_gnd_net_\,
            in3 => \N__23289\,
            lcout => \ADC_IAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19650\,
            carryout => \ADC_IAC.n19651\,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.bit_cnt_i3_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25598\,
            in2 => \_gnd_net_\,
            in3 => \N__23286\,
            lcout => \ADC_IAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19651\,
            carryout => \ADC_IAC.n19652\,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.bit_cnt_i4_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25584\,
            in2 => \_gnd_net_\,
            in3 => \N__23283\,
            lcout => \ADC_IAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19652\,
            carryout => \ADC_IAC.n19653\,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.bit_cnt_i5_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25611\,
            in2 => \_gnd_net_\,
            in3 => \N__23280\,
            lcout => \ADC_IAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19653\,
            carryout => \ADC_IAC.n19654\,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.bit_cnt_i6_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25436\,
            in2 => \_gnd_net_\,
            in3 => \N__23526\,
            lcout => \ADC_IAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19654\,
            carryout => \ADC_IAC.n19655\,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.bit_cnt_i7_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25559\,
            in2 => \_gnd_net_\,
            in3 => \N__23523\,
            lcout => \ADC_IAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54411\,
            ce => \N__25878\,
            sr => \N__23520\
        );

    \ADC_IAC.adc_state_i0_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__35402\,
            in1 => \N__29890\,
            in2 => \N__29996\,
            in3 => \N__25542\,
            lcout => adc_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54420\,
            ce => \N__25635\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.i30_4_lut_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001010001"
        )
    port map (
            in0 => \N__29967\,
            in1 => \N__29899\,
            in2 => \N__25922\,
            in3 => \N__25392\,
            lcout => OPEN,
            ltout => \ADC_IAC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19367_2_lut_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23508\,
            in3 => \N__35401\,
            lcout => \ADC_IAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i8_4_lut_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23498\,
            in1 => \N__23486\,
            in2 => \N__23475\,
            in3 => \N__23459\,
            lcout => \ADC_VDC.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i9_4_lut_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__23441\,
            in1 => \N__23429\,
            in2 => \N__23418\,
            in3 => \N__23402\,
            lcout => \ADC_VDC.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i16_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25685\,
            in1 => \N__48797\,
            in2 => \N__23363\,
            in3 => \N__23385\,
            lcout => buf_adcdata_vdc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_21_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011100000"
        )
    port map (
            in0 => \N__48563\,
            in1 => \N__47367\,
            in2 => \N__48851\,
            in3 => \N__48349\,
            lcout => \ADC_VDC.n12899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i8_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48796\,
            in1 => \N__25686\,
            in2 => \N__23672\,
            in3 => \N__23694\,
            lcout => buf_adcdata_vdc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__48564\,
            in1 => \N__23579\,
            in2 => \N__24161\,
            in3 => \N__23807\,
            lcout => cmd_rdadctmp_5_adj_1474,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25687\,
            in1 => \N__48846\,
            in2 => \N__32864\,
            in3 => \N__23655\,
            lcout => buf_adcdata_vdc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i2_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48845\,
            in1 => \N__25688\,
            in2 => \N__28226\,
            in3 => \N__23643\,
            lcout => buf_adcdata_vdc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__48565\,
            in1 => \N__23557\,
            in2 => \N__24012\,
            in3 => \N__23814\,
            lcout => cmd_rdadctmp_9_adj_1470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__23944\,
            in1 => \N__23631\,
            in2 => \N__23839\,
            in3 => \N__48566\,
            lcout => cmd_rdadctmp_15_adj_1464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i4_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__23578\,
            in1 => \N__23600\,
            in2 => \N__23840\,
            in3 => \N__48567\,
            lcout => cmd_rdadctmp_4_adj_1475,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__24107\,
            in1 => \N__23558\,
            in2 => \N__23894\,
            in3 => \N__48579\,
            lcout => cmd_rdadctmp_8_adj_1471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i7_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__23538\,
            in1 => \N__24308\,
            in2 => \N__25752\,
            in3 => \N__48834\,
            lcout => buf_adcdata_vdc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i6_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__24127\,
            in1 => \N__24162\,
            in2 => \N__23893\,
            in3 => \N__48578\,
            lcout => cmd_rdadctmp_6_adj_1473,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i7_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__48576\,
            in1 => \N__24108\,
            in2 => \N__24135\,
            in3 => \N__23880\,
            lcout => cmd_rdadctmp_7_adj_1472,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48832\,
            in1 => \N__25736\,
            in2 => \N__24080\,
            in3 => \N__24093\,
            lcout => buf_adcdata_vdc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i13_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__48575\,
            in1 => \N__24063\,
            in2 => \N__24039\,
            in3 => \N__23876\,
            lcout => cmd_rdadctmp_13_adj_1466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i10_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__23983\,
            in1 => \N__24010\,
            in2 => \N__23892\,
            in3 => \N__48577\,
            lcout => cmd_rdadctmp_10_adj_1469,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i3_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25735\,
            in1 => \N__48833\,
            in2 => \N__27866\,
            in3 => \N__23964\,
            lcout => buf_adcdata_vdc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i16_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__23921\,
            in1 => \N__23949\,
            in2 => \N__23895\,
            in3 => \N__48591\,
            lcout => cmd_rdadctmp_16_adj_1463,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i19_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48590\,
            in1 => \N__23887\,
            in2 => \N__23735\,
            in3 => \N__23766\,
            lcout => cmd_rdadctmp_19_adj_1460,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i14_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__23709\,
            in1 => \N__46364\,
            in2 => \N__48872\,
            in3 => \N__25742\,
            lcout => buf_adcdata_vdc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i13_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25741\,
            in1 => \N__48854\,
            in2 => \N__24965\,
            in3 => \N__24366\,
            lcout => buf_adcdata_vdc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i6_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__24354\,
            in1 => \N__24332\,
            in2 => \N__48873\,
            in3 => \N__25743\,
            lcout => buf_adcdata_vdc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i12_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25740\,
            in1 => \N__48853\,
            in2 => \N__24608\,
            in3 => \N__24321\,
            lcout => buf_adcdata_vdc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i19_3_lut_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24309\,
            in1 => \N__57699\,
            in2 => \_gnd_net_\,
            in3 => \N__24293\,
            lcout => n19_adj_1623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i9_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25744\,
            in1 => \N__48855\,
            in2 => \N__34958\,
            in3 => \N__24270\,
            lcout => buf_adcdata_vdc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i11_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25745\,
            in1 => \N__48865\,
            in2 => \N__50939\,
            in3 => \N__24258\,
            lcout => buf_adcdata_vdc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i17_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48862\,
            in1 => \N__25746\,
            in2 => \N__24453\,
            in3 => \N__24246\,
            lcout => buf_adcdata_vdc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i23_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25751\,
            in1 => \N__48868\,
            in2 => \N__24207\,
            in3 => \N__24234\,
            lcout => buf_adcdata_vdc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16192_3_lut_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24206\,
            in1 => \N__24185\,
            in2 => \_gnd_net_\,
            in3 => \N__57776\,
            lcout => n19_adj_1527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i21_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25750\,
            in1 => \N__48867\,
            in2 => \N__24569\,
            in3 => \N__24585\,
            lcout => buf_adcdata_vdc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i20_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48864\,
            in1 => \N__25749\,
            in2 => \N__25058\,
            in3 => \N__24552\,
            lcout => buf_adcdata_vdc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i19_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25748\,
            in1 => \N__48866\,
            in2 => \N__25235\,
            in3 => \N__24540\,
            lcout => buf_adcdata_vdc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i18_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48863\,
            in1 => \N__25747\,
            in2 => \N__27101\,
            in3 => \N__24528\,
            lcout => buf_adcdata_vdc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i15_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33345\,
            in1 => \N__33673\,
            in2 => \N__24516\,
            in3 => \N__50201\,
            lcout => buf_adcdata_vac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i18_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33672\,
            in1 => \N__33347\,
            in2 => \N__24489\,
            in3 => \N__27080\,
            lcout => buf_adcdata_vac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22441_bdd_4_lut_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__24379\,
            in1 => \N__24452\,
            in2 => \N__24438\,
            in3 => \N__55175\,
            lcout => n22444,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i17_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33671\,
            in1 => \N__33346\,
            in2 => \N__24423\,
            in3 => \N__24380\,
            lcout => buf_adcdata_vac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i7_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__28098\,
            in1 => \N__27045\,
            in2 => \N__24743\,
            in3 => \N__35579\,
            lcout => cmd_rdadctmp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i22_3_lut_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53777\,
            in1 => \N__24833\,
            in2 => \_gnd_net_\,
            in3 => \N__24804\,
            lcout => OPEN,
            ltout => \n22_adj_1624_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i30_3_lut_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__54706\,
            in1 => \N__24795\,
            in2 => \N__24780\,
            in3 => \_gnd_net_\,
            lcout => n30_adj_1625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101000000"
        )
    port map (
            in0 => \N__34610\,
            in1 => \N__34463\,
            in2 => \N__34797\,
            in3 => \N__24763\,
            lcout => bit_cnt_0_adj_1456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15170_2_lut_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51905\,
            in2 => \_gnd_net_\,
            in3 => \N__49493\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__26867\,
            in1 => \N__28093\,
            in2 => \N__24747\,
            in3 => \N__35616\,
            lcout => cmd_rdadctmp_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.MOSI_31_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34776\,
            in1 => \_gnd_net_\,
            in2 => \N__27228\,
            in3 => \N__24707\,
            lcout => \DDS_MOSI1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19783_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__24678\,
            in1 => \N__55169\,
            in2 => \N__24636\,
            in3 => \N__57642\,
            lcout => n22435,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i8_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__27200\,
            in1 => \N__40669\,
            in2 => \N__43835\,
            in3 => \N__44975\,
            lcout => buf_dds1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i19_3_lut_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57668\,
            in1 => \N__24850\,
            in2 => \_gnd_net_\,
            in3 => \N__24612\,
            lcout => n19_adj_1511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33477\,
            in1 => \N__31515\,
            in2 => \N__24879\,
            in3 => \N__31686\,
            lcout => cmd_rdadctmp_20_adj_1430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i14_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__28606\,
            in1 => \N__40670\,
            in2 => \N__45339\,
            in3 => \N__44976\,
            lcout => buf_dds1_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i19_3_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24969\,
            in1 => \N__24916\,
            in2 => \_gnd_net_\,
            in3 => \N__57667\,
            lcout => n19_adj_1497,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i21_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__31687\,
            in1 => \N__24877\,
            in2 => \N__24947\,
            in3 => \N__33480\,
            lcout => cmd_rdadctmp_21_adj_1429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i9_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__33478\,
            in1 => \N__33733\,
            in2 => \N__26930\,
            in3 => \N__31688\,
            lcout => cmd_rdadctmp_9_adj_1441,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i13_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__24917\,
            in1 => \N__33658\,
            in2 => \N__24948\,
            in3 => \N__33479\,
            lcout => buf_adcdata_vac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i14_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__33476\,
            in1 => \N__24901\,
            in2 => \N__33679\,
            in3 => \N__46342\,
            lcout => buf_adcdata_vac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i12_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35776\,
            in1 => \N__35557\,
            in2 => \N__25041\,
            in3 => \N__46255\,
            lcout => buf_adcdata_iac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i12_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__33456\,
            in1 => \N__24878\,
            in2 => \N__33674\,
            in3 => \N__24854\,
            lcout => buf_adcdata_vac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i7_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__56552\,
            in1 => \N__27264\,
            in2 => \N__31280\,
            in3 => \N__42803\,
            lcout => \buf_cfgRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35555\,
            in1 => \N__25131\,
            in2 => \N__27374\,
            in3 => \N__28114\,
            lcout => cmd_rdadctmp_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i27_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35556\,
            in1 => \N__27321\,
            in2 => \N__27590\,
            in3 => \N__28115\,
            lcout => cmd_rdadctmp_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22417_bdd_4_lut_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__25104\,
            in1 => \N__25090\,
            in2 => \N__25062\,
            in3 => \N__55173\,
            lcout => n22420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i21_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35554\,
            in1 => \N__25037\,
            in2 => \N__35233\,
            in3 => \N__28113\,
            lcout => cmd_rdadctmp_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18528_3_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27201\,
            in1 => \N__32036\,
            in2 => \_gnd_net_\,
            in3 => \N__57796\,
            lcout => OPEN,
            ltout => \n21138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22291_bdd_4_lut_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__25017\,
            in1 => \N__25011\,
            in2 => \N__25005\,
            in3 => \N__53781\,
            lcout => n22294,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i21_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__35757\,
            in1 => \N__35529\,
            in2 => \N__24998\,
            in3 => \N__25201\,
            lcout => buf_adcdata_iac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i29_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__35527\,
            in1 => \N__28116\,
            in2 => \N__25205\,
            in3 => \N__27551\,
            lcout => cmd_rdadctmp_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i22_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__35758\,
            in1 => \N__25183\,
            in2 => \N__31933\,
            in3 => \N__35530\,
            lcout => buf_adcdata_iac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i31_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__35528\,
            in1 => \N__28117\,
            in2 => \N__25185\,
            in3 => \N__25217\,
            lcout => cmd_rdadctmp_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22435_bdd_4_lut_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__25286\,
            in1 => \N__25251\,
            in2 => \N__25242\,
            in3 => \N__55174\,
            lcout => n21076,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i23_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__35526\,
            in1 => \N__35759\,
            in2 => \N__25157\,
            in3 => \N__25218\,
            lcout => buf_adcdata_iac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i19_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35805\,
            in1 => \N__35553\,
            in2 => \N__27591\,
            in3 => \N__43216\,
            lcout => buf_adcdata_iac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i30_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35552\,
            in1 => \N__25206\,
            in2 => \N__25184\,
            in3 => \N__28092\,
            lcout => cmd_rdadctmp_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i15_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__27479\,
            in1 => \N__44977\,
            in2 => \N__40674\,
            in3 => \N__42810\,
            lcout => buf_dds1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i17_3_lut_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25150\,
            in1 => \N__25351\,
            in2 => \_gnd_net_\,
            in3 => \N__57792\,
            lcout => n17_adj_1526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_6_i16_3_lut_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28607\,
            in1 => \N__29428\,
            in2 => \_gnd_net_\,
            in3 => \N__57793\,
            lcout => n16_adj_1534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i14_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__29429\,
            in1 => \N__56498\,
            in2 => \N__45363\,
            in3 => \N__47986\,
            lcout => buf_dds0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i8_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56497\,
            in1 => \N__44860\,
            in2 => \N__42815\,
            in3 => \N__25352\,
            lcout => \VAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.bit_cnt_i0_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25485\,
            in2 => \_gnd_net_\,
            in3 => \N__25338\,
            lcout => \ADC_VAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \ADC_VAC.n19656\,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_VAC.bit_cnt_i1_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25511\,
            in2 => \_gnd_net_\,
            in3 => \N__25335\,
            lcout => \ADC_VAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19656\,
            carryout => \ADC_VAC.n19657\,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_VAC.bit_cnt_i2_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25497\,
            in2 => \_gnd_net_\,
            in3 => \N__25332\,
            lcout => \ADC_VAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19657\,
            carryout => \ADC_VAC.n19658\,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_VAC.bit_cnt_i3_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25524\,
            in2 => \_gnd_net_\,
            in3 => \N__25329\,
            lcout => \ADC_VAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19658\,
            carryout => \ADC_VAC.n19659\,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_VAC.bit_cnt_i4_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25536\,
            in2 => \_gnd_net_\,
            in3 => \N__25326\,
            lcout => \ADC_VAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19659\,
            carryout => \ADC_VAC.n19660\,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_VAC.bit_cnt_i5_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25316\,
            in2 => \_gnd_net_\,
            in3 => \N__25299\,
            lcout => \ADC_VAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19660\,
            carryout => \ADC_VAC.n19661\,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_VAC.bit_cnt_i6_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25473\,
            in2 => \_gnd_net_\,
            in3 => \N__25296\,
            lcout => \ADC_VAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19661\,
            carryout => \ADC_VAC.n19662\,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_VAC.bit_cnt_i7_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25458\,
            in2 => \_gnd_net_\,
            in3 => \N__25293\,
            lcout => \ADC_VAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54383\,
            ce => \N__30749\,
            sr => \N__30639\
        );

    \ADC_IAC.i1_4_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__30001\,
            in1 => \N__35394\,
            in2 => \N__25941\,
            in3 => \N__25391\,
            lcout => OPEN,
            ltout => \ADC_IAC.n20960_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_2_lut_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25638\,
            in3 => \N__29911\,
            lcout => \ADC_IAC.n20961\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19262_4_lut_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__25622\,
            in1 => \N__25610\,
            in2 => \N__25599\,
            in3 => \N__25583\,
            lcout => OPEN,
            ltout => \ADC_IAC.n21295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19068_4_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25572\,
            in1 => \N__25560\,
            in2 => \N__25545\,
            in3 => \N__25410\,
            lcout => \ADC_IAC.n21294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i18419_4_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25535\,
            in1 => \N__25523\,
            in2 => \N__25512\,
            in3 => \N__25496\,
            lcout => OPEN,
            ltout => \ADC_VAC.n21029_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i18433_4_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25484\,
            in1 => \N__25472\,
            in2 => \N__25461\,
            in3 => \N__25457\,
            lcout => \ADC_VAC.n21043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i6_4_lut_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__35325\,
            in1 => \N__29910\,
            in2 => \N__25437\,
            in3 => \N__25421\,
            lcout => \ADC_IAC.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_trig_300_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__30308\,
            in1 => \N__30180\,
            in2 => \N__25402\,
            in3 => \N__37297\,
            lcout => acadc_trig,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_trig_300C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_adj_3_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000100"
        )
    port map (
            in0 => \N__35324\,
            in1 => \N__30000\,
            in2 => \N__25940\,
            in3 => \N__29909\,
            lcout => \ADC_IAC.n12473\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_91_2_lut_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27810\,
            in2 => \_gnd_net_\,
            in3 => \N__55831\,
            lcout => \comm_spi.iclk_N_763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19333_4_lut_4_lut_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101011"
        )
    port map (
            in0 => \N__48528\,
            in1 => \N__48338\,
            in2 => \N__48836\,
            in3 => \N__47383\,
            lcout => OPEN,
            ltout => \ADC_VDC.n11676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.SCLK_46_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__48339\,
            in1 => \N__25835\,
            in2 => \N__25854\,
            in3 => \N__27849\,
            lcout => \VDC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_12178_12179_reset_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27822\,
            lcout => \comm_spi.n14597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54270\,
            ce => 'H',
            sr => \N__25824\
        );

    \ADC_VDC.ADC_DATA_i22_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__25684\,
            in1 => \N__25812\,
            in2 => \N__40451\,
            in3 => \N__48800\,
            lcout => buf_adcdata_vdc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i0_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__25682\,
            in1 => \N__48799\,
            in2 => \N__25964\,
            in3 => \N__25791\,
            lcout => buf_adcdata_vdc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i10_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__35972\,
            in1 => \N__48804\,
            in2 => \N__25773\,
            in3 => \N__25683\,
            lcout => buf_adcdata_vdc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_adj_20_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__48538\,
            in1 => \N__48345\,
            in2 => \N__48852\,
            in3 => \N__47366\,
            lcout => n13087,
            ltout => \n13087_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i15_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__50231\,
            in1 => \N__48805\,
            in2 => \N__26076\,
            in3 => \N__26073\,
            lcout => buf_adcdata_vdc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_19_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48537\,
            in2 => \_gnd_net_\,
            in3 => \N__48798\,
            lcout => \ADC_VDC.n20656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__26055\,
            in1 => \N__48346\,
            in2 => \N__26024\,
            in3 => \N__32733\,
            lcout => \ADC_VDC.cmd_rdadctmp_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53255\,
            ce => \N__26004\,
            sr => \N__25992\
        );

    \comm_spi.i19415_4_lut_3_lut_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__55833\,
            in1 => \_gnd_net_\,
            in2 => \N__27828\,
            in3 => \N__25983\,
            lcout => \comm_spi.n22860\,
            ltout => \comm_spi.n22860_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12180_3_lut_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27780\,
            in2 => \N__25977\,
            in3 => \N__25974\,
            lcout => \comm_spi.iclk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_90_2_lut_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27824\,
            in2 => \_gnd_net_\,
            in3 => \N__55832\,
            lcout => \comm_spi.iclk_N_762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i19_3_lut_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25965\,
            in1 => \N__26893\,
            in2 => \_gnd_net_\,
            in3 => \N__57756\,
            lcout => OPEN,
            ltout => \n19_adj_1484_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i22_3_lut_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26959\,
            in2 => \N__25947\,
            in3 => \N__53771\,
            lcout => OPEN,
            ltout => \n22_adj_1483_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i30_3_lut_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54754\,
            in2 => \N__25944\,
            in3 => \N__26991\,
            lcout => n30_adj_1482,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i0_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__35815\,
            in1 => \N__26879\,
            in2 => \N__26966\,
            in3 => \N__35636\,
            lcout => buf_adcdata_iac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33675\,
            in1 => \N__33501\,
            in2 => \N__26940\,
            in3 => \N__26894\,
            lcout => buf_adcdata_vac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i9_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35635\,
            in1 => \N__28153\,
            in2 => \N__26880\,
            in3 => \N__28125\,
            lcout => cmd_rdadctmp_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.bit_cnt_3767__i3_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__28438\,
            in1 => \N__35884\,
            in2 => \N__28422\,
            in3 => \N__28458\,
            lcout => \comm_spi.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__55870\
        );

    \comm_spi.bit_cnt_3767__i2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__28457\,
            in1 => \N__28418\,
            in2 => \_gnd_net_\,
            in3 => \N__28439\,
            lcout => \comm_spi.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__55870\
        );

    \comm_spi.bit_cnt_3767__i1_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28456\,
            lcout => \comm_spi.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__55870\
        );

    \comm_spi.bit_cnt_3767__i0_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28416\,
            lcout => \comm_spi.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__55870\
        );

    \RTD.i1_3_lut_4_lut_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010010100"
        )
    port map (
            in0 => \N__26850\,
            in1 => \N__26598\,
            in2 => \N__26448\,
            in3 => \N__26264\,
            lcout => \RTD.n15065\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i12467_3_lut_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__42288\,
            in1 => \N__41334\,
            in2 => \_gnd_net_\,
            in3 => \N__43070\,
            lcout => n14884,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.SCLK_27_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000110001"
        )
    port map (
            in0 => \N__34749\,
            in1 => \N__34609\,
            in2 => \N__27119\,
            in3 => \N__34457\,
            lcout => \DDS_SCK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18471_3_lut_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27102\,
            in1 => \N__27076\,
            in2 => \_gnd_net_\,
            in3 => \N__57737\,
            lcout => n21081,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i6_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__27015\,
            in1 => \N__35570\,
            in2 => \N__28122\,
            in3 => \N__27044\,
            lcout => cmd_rdadctmp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i5_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__27033\,
            in1 => \N__28099\,
            in2 => \N__35621\,
            in3 => \N__27014\,
            lcout => cmd_rdadctmp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19404_2_lut_3_lut_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__37317\,
            in1 => \N__30309\,
            in2 => \_gnd_net_\,
            in3 => \N__40890\,
            lcout => n21037,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i4_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__35004\,
            in1 => \N__46762\,
            in2 => \N__57004\,
            in3 => \N__39530\,
            lcout => comm_buf_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i2_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__39686\,
            in1 => \N__56868\,
            in2 => \N__47223\,
            in3 => \N__35003\,
            lcout => comm_buf_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i11_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33670\,
            in1 => \N__33344\,
            in2 => \N__50920\,
            in3 => \N__31514\,
            lcout => buf_adcdata_vac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i7_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27006\,
            lcout => buf_control_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54304\,
            ce => \N__27153\,
            sr => \N__39573\
        );

    \i1_2_lut_adj_225_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__49491\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55515\,
            lcout => OPEN,
            ltout => \n11347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_262_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__57064\,
            in1 => \N__49601\,
            in2 => \N__27156\,
            in3 => \N__52011\,
            lcout => n11919,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i23_3_lut_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27147\,
            in1 => \N__57641\,
            in2 => \_gnd_net_\,
            in3 => \N__32370\,
            lcout => n23_adj_1529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15166_2_lut_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__57062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49490\,
            lcout => n17564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_309_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55513\,
            in2 => \_gnd_net_\,
            in3 => \N__57061\,
            lcout => n12219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12096_2_lut_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__57063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52010\,
            lcout => n14506,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15336_2_lut_3_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52009\,
            in1 => \N__45340\,
            in2 => \_gnd_net_\,
            in3 => \N__55514\,
            lcout => n14_adj_1576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i10_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__34612\,
            in1 => \N__34785\,
            in2 => \N__29385\,
            in3 => \N__31806\,
            lcout => \CLK_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i11_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__34780\,
            in1 => \N__34615\,
            in2 => \N__27141\,
            in3 => \N__43971\,
            lcout => \CLK_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i12_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__34613\,
            in1 => \N__34786\,
            in2 => \N__27246\,
            in3 => \N__40317\,
            lcout => \CLK_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i13_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__34781\,
            in1 => \N__34616\,
            in2 => \N__27237\,
            in3 => \N__27175\,
            lcout => \CLK_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__34611\,
            in1 => \N__34784\,
            in2 => \N__27227\,
            in3 => \N__33924\,
            lcout => \CLK_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i15_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__34782\,
            in1 => \N__34617\,
            in2 => \N__28578\,
            in3 => \N__27480\,
            lcout => tmp_buf_15_adj_1455,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i7_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__34614\,
            in1 => \N__34787\,
            in2 => \N__33855\,
            in3 => \N__28518\,
            lcout => \CLK_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i8_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__34783\,
            in1 => \N__34618\,
            in2 => \N__27210\,
            in3 => \N__27199\,
            lcout => \CLK_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54317\,
            ce => \N__34386\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i20_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35617\,
            in1 => \N__35779\,
            in2 => \N__27558\,
            in3 => \N__40369\,
            lcout => buf_adcdata_iac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i13_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111110101010"
        )
    port map (
            in0 => \N__27176\,
            in1 => \N__37728\,
            in2 => \N__57132\,
            in3 => \N__44978\,
            lcout => buf_dds1_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i12_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56550\,
            in1 => \N__40339\,
            in2 => \N__41493\,
            in3 => \N__48009\,
            lcout => buf_dds0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i18_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35778\,
            in1 => \N__35620\,
            in2 => \N__27320\,
            in3 => \N__40696\,
            lcout => buf_adcdata_iac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i7_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56551\,
            in1 => \N__32321\,
            in2 => \N__50320\,
            in3 => \N__48010\,
            lcout => buf_dds0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i16_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35777\,
            in1 => \N__35619\,
            in2 => \N__27375\,
            in3 => \N__27343\,
            lcout => buf_adcdata_iac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i26_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__35618\,
            in1 => \N__27313\,
            in2 => \N__28124\,
            in3 => \N__31963\,
            lcout => cmd_rdadctmp_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i16_3_lut_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33848\,
            in1 => \N__32317\,
            in2 => \_gnd_net_\,
            in3 => \N__57739\,
            lcout => n16_adj_1504,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i16_3_lut_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33884\,
            in1 => \N__29449\,
            in2 => \_gnd_net_\,
            in3 => \N__57665\,
            lcout => n16_adj_1496,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_252_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__57098\,
            in1 => \N__41533\,
            in2 => \N__56549\,
            in3 => \N__34116\,
            lcout => n12395,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19058_2_lut_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57666\,
            in2 => \_gnd_net_\,
            in3 => \N__36231\,
            lcout => n21285,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i11_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__43993\,
            in1 => \N__56488\,
            in2 => \N__44227\,
            in3 => \N__47995\,
            lcout => buf_dds0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i5_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__47996\,
            in1 => \N__56499\,
            in2 => \N__29454\,
            in3 => \N__51437\,
            lcout => buf_dds0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i28_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__27586\,
            in1 => \N__28064\,
            in2 => \N__35598\,
            in3 => \N__27550\,
            lcout => cmd_rdadctmp_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i2_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44849\,
            in1 => \N__56500\,
            in2 => \N__40156\,
            in3 => \N__39787\,
            lcout => \IAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54344\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19654_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__27534\,
            in1 => \N__55057\,
            in2 => \N__31242\,
            in3 => \N__53680\,
            lcout => OPEN,
            ltout => \n22279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22279_bdd_4_lut_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__53681\,
            in1 => \N__27459\,
            in2 => \N__27519\,
            in3 => \N__27516\,
            lcout => n22282,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19749_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__55058\,
            in1 => \N__53682\,
            in2 => \N__52671\,
            in3 => \N__30042\,
            lcout => OPEN,
            ltout => \n22363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22363_bdd_4_lut_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__53683\,
            in1 => \N__27510\,
            in2 => \N__27501\,
            in3 => \N__27498\,
            lcout => OPEN,
            ltout => \n22366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1553158_i1_3_lut_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27489\,
            in2 => \N__27483\,
            in3 => \N__54719\,
            lcout => n30_adj_1531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i16_3_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27475\,
            in1 => \N__32074\,
            in2 => \_gnd_net_\,
            in3 => \N__57783\,
            lcout => n16_adj_1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.DTRIG_39_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__30729\,
            in1 => \N__27453\,
            in2 => \N__33457\,
            in3 => \N__32211\,
            lcout => acadc_dtrig_v,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i9_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56480\,
            in1 => \N__39727\,
            in2 => \N__40160\,
            in3 => \N__47969\,
            lcout => buf_dds0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__43831\,
            in1 => \N__44856\,
            in2 => \N__27625\,
            in3 => \N__56484\,
            lcout => \IAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i15_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56479\,
            in1 => \N__32078\,
            in2 => \N__42814\,
            in3 => \N__47967\,
            lcout => buf_dds0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i8_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__47968\,
            in1 => \N__56482\,
            in2 => \N__43836\,
            in3 => \N__32035\,
            lcout => buf_dds0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_327_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44787\,
            in1 => \N__36254\,
            in2 => \_gnd_net_\,
            in3 => \N__40884\,
            lcout => acadc_rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i4_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__41494\,
            in1 => \N__41861\,
            in2 => \N__31849\,
            in3 => \N__56483\,
            lcout => \VDC_RNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_247_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__56478\,
            in1 => \N__30195\,
            in2 => \_gnd_net_\,
            in3 => \N__57096\,
            lcout => n12367,
            ltout => \n12367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i1_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__37448\,
            in1 => \N__56481\,
            in2 => \N__27597\,
            in3 => \N__32134\,
            lcout => buf_dds0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14145_4_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110111"
        )
    port map (
            in0 => \N__43910\,
            in1 => \N__30018\,
            in2 => \N__34041\,
            in3 => \N__30285\,
            lcout => OPEN,
            ltout => \n16563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i0_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000010001"
        )
    port map (
            in0 => \N__30286\,
            in1 => \N__30118\,
            in2 => \N__27594\,
            in3 => \N__27765\,
            lcout => eis_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__30075\,
            sr => \N__40891\
        );

    \eis_state_1__bdd_4_lut_4_lut_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100011111000"
        )
    port map (
            in0 => \N__30116\,
            in1 => \N__30036\,
            in2 => \N__37300\,
            in3 => \N__29798\,
            lcout => n22255,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3787_3_lut_3_lut_4_lut_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30117\,
            in1 => \N__40864\,
            in2 => \N__37299\,
            in3 => \N__29799\,
            lcout => \iac_raw_buf_N_734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19371_4_lut_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__40863\,
            in1 => \N__37272\,
            in2 => \N__30302\,
            in3 => \N__30114\,
            lcout => n11654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_260_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__30115\,
            in1 => \N__30281\,
            in2 => \N__37298\,
            in3 => \N__40862\,
            lcout => n13457,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i1_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__30127\,
            in1 => \N__29787\,
            in2 => \N__37309\,
            in3 => \N__30171\,
            lcout => eis_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__30075\,
            sr => \N__40891\
        );

    \data_index_i4_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__47640\,
            in1 => \N__56504\,
            in2 => \N__57144\,
            in3 => \N__47622\,
            lcout => data_index_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_start_329_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43830\,
            in1 => \N__36258\,
            in2 => \_gnd_net_\,
            in3 => \N__43905\,
            lcout => eis_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i1_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56505\,
            in1 => \N__44328\,
            in2 => \N__37455\,
            in3 => \N__37115\,
            lcout => \acadc_skipCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_280_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100001011"
        )
    port map (
            in0 => \N__49602\,
            in1 => \N__30191\,
            in2 => \N__56553\,
            in3 => \N__57139\,
            lcout => n11396,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_200_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43904\,
            in2 => \_gnd_net_\,
            in3 => \N__30017\,
            lcout => n16571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19342_2_lut_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48759\,
            in2 => \_gnd_net_\,
            in3 => \N__48457\,
            lcout => \ADC_VDC.n21952\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.MISO_48_12186_12187_reset_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31422\,
            in1 => \N__30765\,
            in2 => \_gnd_net_\,
            in3 => \N__35176\,
            lcout => \comm_spi.n14605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12186_12187_resetC_net\,
            ce => 'H',
            sr => \N__35107\
        );

    \clk_cnt_3761_3762__i1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30606\,
            in2 => \_gnd_net_\,
            in3 => \N__27843\,
            lcout => clk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => n19746,
            clk => \N__38741\,
            ce => 'H',
            sr => \N__30543\
        );

    \clk_cnt_3761_3762__i2_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30569\,
            in2 => \_gnd_net_\,
            in3 => \N__27840\,
            lcout => clk_cnt_1,
            ltout => OPEN,
            carryin => n19746,
            carryout => n19747,
            clk => \N__38741\,
            ce => 'H',
            sr => \N__30543\
        );

    \clk_cnt_3761_3762__i3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30582\,
            in2 => \_gnd_net_\,
            in3 => \N__27837\,
            lcout => clk_cnt_2,
            ltout => OPEN,
            carryin => n19747,
            carryout => n19748,
            clk => \N__38741\,
            ce => 'H',
            sr => \N__30543\
        );

    \clk_cnt_3761_3762__i4_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30555\,
            in2 => \_gnd_net_\,
            in3 => \N__27834\,
            lcout => clk_cnt_3,
            ltout => OPEN,
            carryin => n19748,
            carryout => n19749,
            clk => \N__38741\,
            ce => 'H',
            sr => \N__30543\
        );

    \clk_cnt_3761_3762__i5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30594\,
            in2 => \_gnd_net_\,
            in3 => \N__27831\,
            lcout => clk_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38741\,
            ce => 'H',
            sr => \N__30543\
        );

    \comm_spi.iclk_40_12178_12179_set_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54272\,
            ce => 'H',
            sr => \N__27774\
        );

    \ADC_IAC.ADC_DATA_i1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__35626\,
            in1 => \N__32842\,
            in2 => \N__35816\,
            in3 => \N__28155\,
            lcout => buf_adcdata_iac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i19_3_lut_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28230\,
            in1 => \N__27886\,
            in2 => \_gnd_net_\,
            in3 => \N__57755\,
            lcout => OPEN,
            ltout => \n19_adj_1639_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i22_3_lut_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28171\,
            in2 => \N__28209\,
            in3 => \N__53722\,
            lcout => n22_adj_1640,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i30_3_lut_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28206\,
            in1 => \N__28194\,
            in2 => \_gnd_net_\,
            in3 => \N__54755\,
            lcout => n30_adj_1631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__35627\,
            in1 => \N__28172\,
            in2 => \N__35817\,
            in3 => \N__28139\,
            lcout => buf_adcdata_iac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__28154\,
            in1 => \N__28066\,
            in2 => \N__28140\,
            in3 => \N__35629\,
            lcout => cmd_rdadctmp_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i11_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__35628\,
            in1 => \N__28138\,
            in2 => \N__28108\,
            in3 => \N__28387\,
            lcout => cmd_rdadctmp_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i2_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__33676\,
            in1 => \N__27887\,
            in2 => \N__33507\,
            in3 => \N__28347\,
            lcout => buf_adcdata_vac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i19_3_lut_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27870\,
            in1 => \N__28360\,
            in2 => \_gnd_net_\,
            in3 => \N__57698\,
            lcout => n19_adj_1636,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i9_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33502\,
            in1 => \N__33663\,
            in2 => \N__34933\,
            in3 => \N__31721\,
            lcout => buf_adcdata_vac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i2_3_lut_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__28455\,
            in1 => \_gnd_net_\,
            in2 => \N__28440\,
            in3 => \N__28415\,
            lcout => \comm_spi.n17036\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i3_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35808\,
            in1 => \N__35630\,
            in2 => \N__28397\,
            in3 => \N__31039\,
            lcout => buf_adcdata_iac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33662\,
            in1 => \N__33504\,
            in2 => \N__28314\,
            in3 => \N__28361\,
            lcout => buf_adcdata_vac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i11_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__33503\,
            in1 => \N__28306\,
            in2 => \N__28346\,
            in3 => \N__31691\,
            lcout => cmd_rdadctmp_11_adj_1439,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i12_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__31692\,
            in1 => \N__28282\,
            in2 => \N__28313\,
            in3 => \N__33505\,
            lcout => cmd_rdadctmp_12_adj_1438,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i30_3_lut_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28260\,
            in1 => \N__28254\,
            in2 => \_gnd_net_\,
            in3 => \N__54756\,
            lcout => n30_adj_1641,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secclk_cnt_3765_3766__i1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31107\,
            in2 => \_gnd_net_\,
            in3 => \N__28239\,
            lcout => secclk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => n19750,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30878\,
            in2 => \_gnd_net_\,
            in3 => \N__28236\,
            lcout => secclk_cnt_1,
            ltout => OPEN,
            carryin => n19750,
            carryout => n19751,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31214\,
            in2 => \_gnd_net_\,
            in3 => \N__28233\,
            lcout => secclk_cnt_2,
            ltout => OPEN,
            carryin => n19751,
            carryout => n19752,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30915\,
            in2 => \_gnd_net_\,
            in3 => \N__28485\,
            lcout => secclk_cnt_3,
            ltout => OPEN,
            carryin => n19752,
            carryout => n19753,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i5_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31068\,
            in2 => \_gnd_net_\,
            in3 => \N__28482\,
            lcout => secclk_cnt_4,
            ltout => OPEN,
            carryin => n19753,
            carryout => n19754,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30864\,
            in2 => \_gnd_net_\,
            in3 => \N__28479\,
            lcout => secclk_cnt_5,
            ltout => OPEN,
            carryin => n19754,
            carryout => n19755,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i7_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30954\,
            in2 => \_gnd_net_\,
            in3 => \N__28476\,
            lcout => secclk_cnt_6,
            ltout => OPEN,
            carryin => n19755,
            carryout => n19756,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i8_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31199\,
            in2 => \_gnd_net_\,
            in3 => \N__28473\,
            lcout => secclk_cnt_7,
            ltout => OPEN,
            carryin => n19756,
            carryout => n19757,
            clk => \N__38746\,
            ce => 'H',
            sr => \N__31145\
        );

    \secclk_cnt_3765_3766__i9_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30891\,
            in2 => \_gnd_net_\,
            in3 => \N__28470\,
            lcout => secclk_cnt_8,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => n19758,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i10_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30996\,
            in2 => \_gnd_net_\,
            in3 => \N__28467\,
            lcout => secclk_cnt_9,
            ltout => OPEN,
            carryin => n19758,
            carryout => n19759,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i11_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30929\,
            in2 => \_gnd_net_\,
            in3 => \N__28464\,
            lcout => secclk_cnt_10,
            ltout => OPEN,
            carryin => n19759,
            carryout => n19760,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i12_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31082\,
            in2 => \_gnd_net_\,
            in3 => \N__28461\,
            lcout => secclk_cnt_11,
            ltout => OPEN,
            carryin => n19760,
            carryout => n19761,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i13_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31457\,
            in2 => \_gnd_net_\,
            in3 => \N__28512\,
            lcout => secclk_cnt_12,
            ltout => OPEN,
            carryin => n19761,
            carryout => n19762,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31188\,
            in2 => \_gnd_net_\,
            in3 => \N__28509\,
            lcout => secclk_cnt_13,
            ltout => OPEN,
            carryin => n19762,
            carryout => n19763,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i15_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30942\,
            in2 => \_gnd_net_\,
            in3 => \N__28506\,
            lcout => secclk_cnt_14,
            ltout => OPEN,
            carryin => n19763,
            carryout => n19764,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i16_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30903\,
            in2 => \_gnd_net_\,
            in3 => \N__28503\,
            lcout => secclk_cnt_15,
            ltout => OPEN,
            carryin => n19764,
            carryout => n19765,
            clk => \N__38747\,
            ce => 'H',
            sr => \N__31138\
        );

    \secclk_cnt_3765_3766__i17_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31227\,
            in2 => \_gnd_net_\,
            in3 => \N__28500\,
            lcout => secclk_cnt_16,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => n19766,
            clk => \N__38748\,
            ce => 'H',
            sr => \N__31146\
        );

    \secclk_cnt_3765_3766__i18_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31008\,
            in2 => \_gnd_net_\,
            in3 => \N__28497\,
            lcout => secclk_cnt_17,
            ltout => OPEN,
            carryin => n19766,
            carryout => n19767,
            clk => \N__38748\,
            ce => 'H',
            sr => \N__31146\
        );

    \secclk_cnt_3765_3766__i19_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31095\,
            in2 => \_gnd_net_\,
            in3 => \N__28494\,
            lcout => secclk_cnt_18,
            ltout => OPEN,
            carryin => n19767,
            carryout => n19768,
            clk => \N__38748\,
            ce => 'H',
            sr => \N__31146\
        );

    \secclk_cnt_3765_3766__i20_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31470\,
            in2 => \_gnd_net_\,
            in3 => \N__28491\,
            lcout => secclk_cnt_19,
            ltout => OPEN,
            carryin => n19768,
            carryout => n19769,
            clk => \N__38748\,
            ce => 'H',
            sr => \N__31146\
        );

    \secclk_cnt_3765_3766__i21_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31158\,
            in2 => \_gnd_net_\,
            in3 => \N__28488\,
            lcout => secclk_cnt_20,
            ltout => OPEN,
            carryin => n19769,
            carryout => n19770,
            clk => \N__38748\,
            ce => 'H',
            sr => \N__31146\
        );

    \secclk_cnt_3765_3766__i22_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31482\,
            in2 => \_gnd_net_\,
            in3 => \N__28620\,
            lcout => secclk_cnt_21,
            ltout => OPEN,
            carryin => n19770,
            carryout => n19771,
            clk => \N__38748\,
            ce => 'H',
            sr => \N__31146\
        );

    \secclk_cnt_3765_3766__i23_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31443\,
            in2 => \_gnd_net_\,
            in3 => \N__28617\,
            lcout => secclk_cnt_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38748\,
            ce => 'H',
            sr => \N__31146\
        );

    \CLK_DDS.tmp_buf_i14_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__34596\,
            in1 => \N__34791\,
            in2 => \N__28614\,
            in3 => \N__28584\,
            lcout => \CLK_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__34788\,
            in1 => \N__34601\,
            in2 => \N__33762\,
            in3 => \N__28569\,
            lcout => \CLK_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__34597\,
            in1 => \N__34792\,
            in2 => \N__28563\,
            in3 => \N__46893\,
            lcout => \CLK_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__46956\,
            in1 => \N__34795\,
            in2 => \N__28554\,
            in3 => \N__34602\,
            lcout => \CLK_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__34598\,
            in1 => \N__34793\,
            in2 => \N__28545\,
            in3 => \N__33999\,
            lcout => \CLK_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__34789\,
            in1 => \N__34600\,
            in2 => \N__28536\,
            in3 => \N__33885\,
            lcout => \CLK_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__34599\,
            in1 => \N__34794\,
            in2 => \N__28527\,
            in3 => \N__40761\,
            lcout => \CLK_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i9_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__34790\,
            in1 => \N__40241\,
            in2 => \N__34619\,
            in3 => \N__29391\,
            lcout => \CLK_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54305\,
            ce => \N__34382\,
            sr => \_gnd_net_\
        );

    \data_count_i0_i0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37953\,
            in2 => \N__29293\,
            in3 => \_gnd_net_\,
            lcout => data_count_0,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => n19586,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29179\,
            in2 => \_gnd_net_\,
            in3 => \N__29160\,
            lcout => data_count_1,
            ltout => OPEN,
            carryin => n19586,
            carryout => n19587,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29074\,
            in2 => \_gnd_net_\,
            in3 => \N__29052\,
            lcout => data_count_2,
            ltout => OPEN,
            carryin => n19587,
            carryout => n19588,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28969\,
            in2 => \_gnd_net_\,
            in3 => \N__28947\,
            lcout => data_count_3,
            ltout => OPEN,
            carryin => n19588,
            carryout => n19589,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28858\,
            in2 => \_gnd_net_\,
            in3 => \N__28836\,
            lcout => data_count_4,
            ltout => OPEN,
            carryin => n19589,
            carryout => n19590,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28753\,
            in2 => \_gnd_net_\,
            in3 => \N__28728\,
            lcout => data_count_5,
            ltout => OPEN,
            carryin => n19590,
            carryout => n19591,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28645\,
            in2 => \_gnd_net_\,
            in3 => \N__28623\,
            lcout => data_count_6,
            ltout => OPEN,
            carryin => n19591,
            carryout => n19592,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i7_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29701\,
            in2 => \_gnd_net_\,
            in3 => \N__29682\,
            lcout => data_count_7,
            ltout => OPEN,
            carryin => n19592,
            carryout => n19593,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38558\,
            sr => \N__38482\
        );

    \data_count_i0_i8_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29593\,
            in2 => \_gnd_net_\,
            in3 => \N__29574\,
            lcout => data_count_8,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => n19594,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__38552\,
            sr => \N__38496\
        );

    \data_count_i0_i9_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29482\,
            in2 => \_gnd_net_\,
            in3 => \N__29571\,
            lcout => data_count_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__38552\,
            sr => \N__38496\
        );

    \SIG_DDS.tmp_buf_i10_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__42268\,
            in1 => \N__43066\,
            in2 => \N__29817\,
            in3 => \N__40980\,
            lcout => \SIG_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i11_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43062\,
            in1 => \N__42272\,
            in2 => \N__29463\,
            in3 => \N__44000\,
            lcout => \SIG_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i5_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__42270\,
            in1 => \N__43068\,
            in2 => \N__32052\,
            in3 => \N__29453\,
            lcout => \SIG_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i13_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43064\,
            in1 => \N__42274\,
            in2 => \N__29400\,
            in3 => \N__41631\,
            lcout => \SIG_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i14_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__42269\,
            in1 => \N__43067\,
            in2 => \N__29436\,
            in3 => \N__29415\,
            lcout => \SIG_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i12_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43063\,
            in1 => \N__42273\,
            in2 => \N__29409\,
            in3 => \N__40346\,
            lcout => \SIG_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i9_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__42271\,
            in1 => \N__43069\,
            in2 => \N__32013\,
            in3 => \N__39728\,
            lcout => \SIG_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i6_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43065\,
            in1 => \N__42275\,
            in2 => \N__29808\,
            in3 => \N__40734\,
            lcout => \SIG_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54345\,
            ce => \N__42090\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_217_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__32177\,
            in1 => \N__30296\,
            in2 => \_gnd_net_\,
            in3 => \N__32207\,
            lcout => n16554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_168_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32439\,
            in1 => \N__32478\,
            in2 => \N__32274\,
            in3 => \N__32290\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_238_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__56519\,
            in1 => \N__57097\,
            in2 => \N__33111\,
            in3 => \N__41778\,
            lcout => n11915,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32176\,
            lcout => \iac_raw_buf_N_736\,
            ltout => \iac_raw_buf_N_736_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011100100"
        )
    port map (
            in0 => \N__30306\,
            in1 => \N__30122\,
            in2 => \N__29790\,
            in3 => \N__37292\,
            lcout => n17_adj_1622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19331_4_lut_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010011"
        )
    port map (
            in0 => \N__37293\,
            in1 => \N__30307\,
            in2 => \N__30135\,
            in3 => \N__32151\,
            lcout => OPEN,
            ltout => \n20826_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_end_299_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__30051\,
            in1 => \N__30297\,
            in2 => \N__29781\,
            in3 => \N__40877\,
            lcout => eis_end,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_end_299C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i26_3_lut_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38004\,
            in1 => \N__57823\,
            in2 => \_gnd_net_\,
            in3 => \N__30050\,
            lcout => n26_adj_1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18989_2_lut_3_lut_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__30295\,
            in1 => \N__32213\,
            in2 => \_gnd_net_\,
            in3 => \N__32174\,
            lcout => n21234,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32376\,
            in1 => \N__41565\,
            in2 => \N__30030\,
            in3 => \N__32382\,
            lcout => OPEN,
            ltout => \n30_adj_1604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29823\,
            in1 => \N__38412\,
            in2 => \N__30021\,
            in3 => \N__29829\,
            lcout => n31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.DTRIG_39_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010101000"
        )
    port map (
            in0 => \N__32175\,
            in1 => \N__35569\,
            in2 => \N__30006\,
            in3 => \N__29912\,
            lcout => acadc_dtrig_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15109_2_lut_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32212\,
            in2 => \_gnd_net_\,
            in3 => \N__32173\,
            lcout => n17507,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_61_i14_2_lut_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32715\,
            in2 => \_gnd_net_\,
            in3 => \N__32239\,
            lcout => OPEN,
            ltout => \n14_adj_1509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__32514\,
            in1 => \N__43639\,
            in2 => \N__29832\,
            in3 => \N__32223\,
            lcout => n26_adj_1508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_170_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32417\,
            in1 => \N__46837\,
            in2 => \N__32556\,
            in3 => \N__37111\,
            lcout => n18_adj_1609,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i4_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56546\,
            in1 => \N__44327\,
            in2 => \N__47801\,
            in3 => \N__46838\,
            lcout => \acadc_skipCount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__55208\,
            in1 => \N__57782\,
            in2 => \N__41540\,
            in3 => \N__53721\,
            lcout => n20915,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18376_4_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__30126\,
            in1 => \N__37291\,
            in2 => \N__30298\,
            in3 => \N__40885\,
            lcout => n20985,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i11_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56545\,
            in1 => \N__44326\,
            in2 => \N__44226\,
            in3 => \N__41926\,
            lcout => \acadc_skipCount_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i2_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__41874\,
            in1 => \N__56547\,
            in2 => \N__44788\,
            in3 => \N__31765\,
            lcout => \SELIRNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19109_2_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30139\,
            in2 => \_gnd_net_\,
            in3 => \N__34037\,
            lcout => n21337,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i34_3_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30140\,
            in1 => \N__37958\,
            in2 => \_gnd_net_\,
            in3 => \N__30170\,
            lcout => OPEN,
            ltout => \n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i2_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__37308\,
            in1 => \N__30274\,
            in2 => \N__30159\,
            in3 => \N__30156\,
            lcout => \eis_end_N_724\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i2C_net\,
            ce => \N__30074\,
            sr => \N__40889\
        );

    \i24_4_lut_adj_188_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__43906\,
            in1 => \N__30150\,
            in2 => \N__30141\,
            in3 => \N__34296\,
            lcout => OPEN,
            ltout => \n11_adj_1621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19384_3_lut_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37307\,
            in2 => \N__30078\,
            in3 => \N__30273\,
            lcout => n11744,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19350_2_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30272\,
            in2 => \_gnd_net_\,
            in3 => \N__32646\,
            lcout => n14671,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7704_3_lut_4_lut_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010010111100"
        )
    port map (
            in0 => \N__48299\,
            in1 => \N__47361\,
            in2 => \N__47490\,
            in3 => \N__34830\,
            lcout => OPEN,
            ltout => \ADC_VDC.n10119_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011111110"
        )
    port map (
            in0 => \N__48760\,
            in1 => \N__48465\,
            in2 => \N__30213\,
            in3 => \N__32568\,
            lcout => \ADC_VDC.n12807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i3_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100001000001010"
        )
    port map (
            in0 => \N__48466\,
            in1 => \N__48279\,
            in2 => \N__48772\,
            in3 => \N__47362\,
            lcout => adc_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53298\,
            ce => \N__30210\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16150_3_lut_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110101010"
        )
    port map (
            in0 => \N__47473\,
            in1 => \N__48278\,
            in2 => \_gnd_net_\,
            in3 => \N__47360\,
            lcout => \ADC_VDC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_10_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48689\,
            in2 => \_gnd_net_\,
            in3 => \N__48464\,
            lcout => \ADC_VDC.n20899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i0_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30801\,
            in2 => \_gnd_net_\,
            in3 => \N__30204\,
            lcout => dds0_mclkcnt_0,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => n19739,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i1_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30839\,
            in2 => \_gnd_net_\,
            in3 => \N__30201\,
            lcout => dds0_mclkcnt_1,
            ltout => OPEN,
            carryin => n19739,
            carryout => n19740,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i2_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30813\,
            in2 => \_gnd_net_\,
            in3 => \N__30198\,
            lcout => dds0_mclkcnt_2,
            ltout => OPEN,
            carryin => n19740,
            carryout => n19741,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i3_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30321\,
            in2 => \_gnd_net_\,
            in3 => \N__30621\,
            lcout => dds0_mclkcnt_3,
            ltout => OPEN,
            carryin => n19741,
            carryout => n19742,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i4_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30825\,
            in2 => \_gnd_net_\,
            in3 => \N__30618\,
            lcout => dds0_mclkcnt_4,
            ltout => OPEN,
            carryin => n19742,
            carryout => n19743,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i5_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30852\,
            in2 => \_gnd_net_\,
            in3 => \N__30615\,
            lcout => dds0_mclkcnt_5,
            ltout => OPEN,
            carryin => n19743,
            carryout => n19744,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i6_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30771\,
            in2 => \_gnd_net_\,
            in3 => \N__30612\,
            lcout => dds0_mclkcnt_6,
            ltout => OPEN,
            carryin => n19744,
            carryout => n19745,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i7_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30786\,
            in2 => \_gnd_net_\,
            in3 => \N__30609\,
            lcout => dds0_mclkcnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_250_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30593\,
            lcout => OPEN,
            ltout => \n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_253_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30581\,
            in1 => \N__30570\,
            in2 => \N__30558\,
            in3 => \N__30554\,
            lcout => n14714,
            ltout => \n14714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_RTD_287_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30531\,
            in3 => \N__30346\,
            lcout => \clk_RTD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30320\,
            in1 => \N__30851\,
            in2 => \N__30840\,
            in3 => \N__30824\,
            lcout => OPEN,
            ltout => \n12_adj_1480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30812\,
            in1 => \N__30800\,
            in2 => \N__30789\,
            in3 => \N__30785\,
            lcout => n20799,
            ltout => \n20799_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15251_2_lut_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30774\,
            in3 => \N__30974\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imiso_83_12192_12193_reset_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35178\,
            in1 => \N__34352\,
            in2 => \_gnd_net_\,
            in3 => \N__32882\,
            lcout => \comm_spi.n14611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12192_12193_resetC_net\,
            ce => 'H',
            sr => \N__35109\
        );

    \comm_spi.MISO_48_12186_12187_set_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31418\,
            in1 => \N__30761\,
            in2 => \_gnd_net_\,
            in3 => \N__35172\,
            lcout => \comm_spi.n14604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12186_12187_setC_net\,
            ce => 'H',
            sr => \N__35045\
        );

    \ADC_VAC.i12431_2_lut_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30750\,
            in2 => \_gnd_net_\,
            in3 => \N__30728\,
            lcout => \ADC_VAC.n14844\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_89_2_lut_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55637\,
            in2 => \_gnd_net_\,
            in3 => \N__55777\,
            lcout => \comm_spi.imosi_N_753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i7_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__35894\,
            in1 => \N__46404\,
            in2 => \_gnd_net_\,
            in3 => \N__35846\,
            lcout => comm_rx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => 'H',
            sr => \N__55869\
        );

    \comm_spi.data_rx_i6_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__35845\,
            in1 => \N__52058\,
            in2 => \_gnd_net_\,
            in3 => \N__35893\,
            lcout => comm_rx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => 'H',
            sr => \N__55869\
        );

    \comm_spi.data_rx_i5_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__35892\,
            in1 => \N__46715\,
            in2 => \_gnd_net_\,
            in3 => \N__35844\,
            lcout => comm_rx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => 'H',
            sr => \N__55869\
        );

    \comm_spi.data_rx_i4_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__35843\,
            in1 => \N__51054\,
            in2 => \_gnd_net_\,
            in3 => \N__35891\,
            lcout => comm_rx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => 'H',
            sr => \N__55869\
        );

    \comm_spi.data_rx_i3_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__35890\,
            in1 => \N__47174\,
            in2 => \_gnd_net_\,
            in3 => \N__35842\,
            lcout => comm_rx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => 'H',
            sr => \N__55869\
        );

    \comm_spi.data_rx_i2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__35841\,
            in1 => \N__45724\,
            in2 => \_gnd_net_\,
            in3 => \N__35889\,
            lcout => comm_rx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => 'H',
            sr => \N__55869\
        );

    \comm_spi.data_rx_i1_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__35888\,
            in1 => \N__35840\,
            in2 => \_gnd_net_\,
            in3 => \N__53050\,
            lcout => comm_rx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => 'H',
            sr => \N__55869\
        );

    \dds0_mclk_294_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__38690\,
            in1 => \N__30978\,
            in2 => \_gnd_net_\,
            in3 => \N__30963\,
            lcout => dds0_mclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclk_294C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i4_4_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43134\,
            in1 => \N__43150\,
            in2 => \N__43098\,
            in3 => \N__41301\,
            lcout => \SIG_DDS.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_196_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30953\,
            in1 => \N__30941\,
            in2 => \N__30930\,
            in3 => \N__30914\,
            lcout => n27_adj_1597,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30902\,
            in1 => \N__30890\,
            in2 => \N__30879\,
            in3 => \N__30863\,
            lcout => n25_adj_1574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_193_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31226\,
            in1 => \N__31215\,
            in2 => \N__31203\,
            in3 => \N__31187\,
            lcout => OPEN,
            ltout => \n26_adj_1575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_205_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31056\,
            in1 => \N__31176\,
            in2 => \N__31170\,
            in3 => \N__31167\,
            lcout => OPEN,
            ltout => \n19856_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_206_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31431\,
            in1 => \N__30984\,
            in2 => \N__31161\,
            in3 => \N__31157\,
            lcout => n14715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_189_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31106\,
            in1 => \N__31094\,
            in2 => \N__31083\,
            in3 => \N__31067\,
            lcout => n28_adj_1505,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__43157\,
            in1 => \N__43061\,
            in2 => \_gnd_net_\,
            in3 => \N__42881\,
            lcout => bit_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i22_3_lut_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__31040\,
            in1 => \N__31017\,
            in2 => \N__53795\,
            in3 => \_gnd_net_\,
            lcout => n22_adj_1637,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31007\,
            in2 => \_gnd_net_\,
            in3 => \N__30995\,
            lcout => n10_adj_1601,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_96_2_lut_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34902\,
            in2 => \_gnd_net_\,
            in3 => \N__55866\,
            lcout => \comm_spi.data_tx_7__N_770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i30_3_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31746\,
            in1 => \N__31728\,
            in2 => \_gnd_net_\,
            in3 => \N__54644\,
            lcout => n30_adj_1638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i18_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__31722\,
            in1 => \N__33494\,
            in2 => \N__33129\,
            in3 => \N__31689\,
            lcout => cmd_rdadctmp_18_adj_1432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i19_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__31690\,
            in1 => \N__31498\,
            in2 => \N__33506\,
            in3 => \N__33127\,
            lcout => cmd_rdadctmp_19_adj_1431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_197_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31481\,
            in1 => \N__31469\,
            in2 => \N__31458\,
            in3 => \N__31442\,
            lcout => n14_adj_1599,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imiso_83_12192_12193_set_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35177\,
            in1 => \N__34359\,
            in2 => \_gnd_net_\,
            in3 => \N__32889\,
            lcout => \comm_spi.n14610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12192_12193_setC_net\,
            ce => 'H',
            sr => \N__35049\
        );

    \mux_128_Mux_6_i20_3_lut_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31404\,
            in1 => \N__31371\,
            in2 => \_gnd_net_\,
            in3 => \N__57383\,
            lcout => n20_adj_1537,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i20_3_lut_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31323\,
            in1 => \N__31287\,
            in2 => \_gnd_net_\,
            in3 => \N__57381\,
            lcout => n20_adj_1528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_0_i16_3_lut_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57382\,
            in1 => \N__33919\,
            in2 => \_gnd_net_\,
            in3 => \N__33968\,
            lcout => n16_adj_1487,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i16_3_lut_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33754\,
            in1 => \N__32145\,
            in2 => \_gnd_net_\,
            in3 => \N__57384\,
            lcout => n16_adj_1521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i11_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__35803\,
            in1 => \N__52774\,
            in2 => \N__32001\,
            in3 => \N__35623\,
            lcout => buf_adcdata_iac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i17_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35622\,
            in1 => \N__35804\,
            in2 => \N__31968\,
            in3 => \N__39754\,
            lcout => buf_adcdata_iac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i13_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37717\,
            in1 => \N__41742\,
            in2 => \_gnd_net_\,
            in3 => \N__33944\,
            lcout => req_data_cnt_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_6_i17_3_lut_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57591\,
            in1 => \N__31937\,
            in2 => \_gnd_net_\,
            in3 => \N__31895\,
            lcout => n17_adj_1535,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i10_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__31802\,
            in1 => \N__40667\,
            in2 => \N__44792\,
            in3 => \N__44957\,
            lcout => buf_dds1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_4_i23_3_lut_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__57590\,
            in1 => \_gnd_net_\,
            in2 => \N__31859\,
            in3 => \N__32295\,
            lcout => n23_adj_1541,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000110011"
        )
    port map (
            in0 => \N__35997\,
            in1 => \N__41284\,
            in2 => \N__31821\,
            in3 => \N__43044\,
            lcout => dds_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54314\,
            ce => \N__36092\,
            sr => \_gnd_net_\
        );

    \i18462_3_lut_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31798\,
            in1 => \N__40976\,
            in2 => \_gnd_net_\,
            in3 => \N__57592\,
            lcout => n21072,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18477_3_lut_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31775\,
            in1 => \N__57593\,
            in2 => \_gnd_net_\,
            in3 => \N__32272\,
            lcout => n21087,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43568\,
            in1 => \N__51879\,
            in2 => \_gnd_net_\,
            in3 => \N__55547\,
            lcout => n14_adj_1583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_256_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55545\,
            in2 => \_gnd_net_\,
            in3 => \N__50052\,
            lcout => n20856,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__36773\,
            in1 => \N__43047\,
            in2 => \N__42287\,
            in3 => \N__33967\,
            lcout => \SIG_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__32144\,
            in1 => \N__32112\,
            in2 => \N__42282\,
            in3 => \N__43052\,
            lcout => \SIG_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i2_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__32106\,
            in1 => \N__42248\,
            in2 => \N__47928\,
            in3 => \N__43049\,
            lcout => \SIG_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__43045\,
            in1 => \N__32100\,
            in2 => \N__42283\,
            in3 => \N__46923\,
            lcout => \SIG_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i15_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__32094\,
            in1 => \N__43048\,
            in2 => \N__32088\,
            in3 => \N__42262\,
            lcout => tmp_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i4_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__33806\,
            in1 => \N__43051\,
            in2 => \N__42284\,
            in3 => \N__32058\,
            lcout => \SIG_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i8_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__32301\,
            in1 => \N__42249\,
            in2 => \N__32043\,
            in3 => \N__43050\,
            lcout => \SIG_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i7_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__43046\,
            in1 => \N__32331\,
            in2 => \N__42285\,
            in3 => \N__32325\,
            lcout => \SIG_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54327\,
            ce => \N__42089\,
            sr => \_gnd_net_\
        );

    \buf_dds0_i4_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56446\,
            in1 => \N__33802\,
            in2 => \N__47805\,
            in3 => \N__47997\,
            lcout => buf_dds0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i12_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56441\,
            in1 => \N__44323\,
            in2 => \N__41495\,
            in3 => \N__32294\,
            lcout => \acadc_skipCount_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i6_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__56445\,
            in1 => \N__41862\,
            in2 => \N__38675\,
            in3 => \N__45353\,
            lcout => buf_control_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i10_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__56440\,
            in1 => \N__44322\,
            in2 => \N__32273\,
            in3 => \N__44779\,
            lcout => \acadc_skipCount_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i13_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__44321\,
            in1 => \N__43589\,
            in2 => \N__56540\,
            in3 => \N__32243\,
            lcout => \acadc_skipCount_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i5_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__52811\,
            in1 => \N__51438\,
            in2 => \N__56539\,
            in3 => \N__44324\,
            lcout => \acadc_skipCount_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32538\,
            in1 => \N__32400\,
            in2 => \N__50087\,
            in3 => \N__52810\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_232_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__32217\,
            in1 => \N__32178\,
            in2 => \_gnd_net_\,
            in3 => \N__34030\,
            lcout => n4_adj_1546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32694\,
            in1 => \N__32457\,
            in2 => \N__41927\,
            in3 => \N__33820\,
            lcout => n23_adj_1501,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__32496\,
            in1 => \N__32673\,
            in2 => \N__34074\,
            in3 => \N__32359\,
            lcout => n24_adj_1642,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i8_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__43649\,
            in1 => \N__43824\,
            in2 => \N__44331\,
            in3 => \N__56471\,
            lcout => \acadc_skipCount_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15345_2_lut_3_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__51878\,
            in1 => \N__37431\,
            in2 => \_gnd_net_\,
            in3 => \N__55546\,
            lcout => n14_adj_1556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i15_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__32360\,
            in1 => \N__56467\,
            in2 => \N__42816\,
            in3 => \N__44299\,
            lcout => \acadc_skipCount_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i9_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__44297\,
            in1 => \N__40121\,
            in2 => \N__56548\,
            in3 => \N__34073\,
            lcout => \acadc_skipCount_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i14_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__33821\,
            in1 => \N__56466\,
            in2 => \N__45358\,
            in3 => \N__44298\,
            lcout => \acadc_skipCount_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37954\,
            in2 => \N__38451\,
            in3 => \_gnd_net_\,
            lcout => acadc_skipcnt_0,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => n19610,
            clk => \INVacadc_skipcnt_i0_i0C_net\,
            ce => \N__32656\,
            sr => \N__32346\
        );

    \add_73_2_THRU_CRY_0_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58608\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => n19610,
            carryout => \n19610_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_1_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__58621\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19610_THRU_CRY_0_THRU_CO\,
            carryout => \n19610_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_2_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58612\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19610_THRU_CRY_1_THRU_CO\,
            carryout => \n19610_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_3_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__58622\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19610_THRU_CRY_2_THRU_CO\,
            carryout => \n19610_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_4_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58616\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19610_THRU_CRY_3_THRU_CO\,
            carryout => \n19610_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_5_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__58623\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19610_THRU_CRY_4_THRU_CO\,
            carryout => \n19610_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_6_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58620\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19610_THRU_CRY_5_THRU_CO\,
            carryout => \n19610_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i1_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32418\,
            in2 => \_gnd_net_\,
            in3 => \N__32406\,
            lcout => acadc_skipcnt_1,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => n19611,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i2_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41579\,
            in2 => \_gnd_net_\,
            in3 => \N__32403\,
            lcout => acadc_skipcnt_2,
            ltout => OPEN,
            carryin => n19611,
            carryout => n19612,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i3_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32399\,
            in2 => \_gnd_net_\,
            in3 => \N__32385\,
            lcout => acadc_skipcnt_3,
            ltout => OPEN,
            carryin => n19612,
            carryout => n19613,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i4_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32555\,
            in2 => \_gnd_net_\,
            in3 => \N__32541\,
            lcout => acadc_skipcnt_4,
            ltout => OPEN,
            carryin => n19613,
            carryout => n19614,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i5_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32537\,
            in2 => \_gnd_net_\,
            in3 => \N__32523\,
            lcout => acadc_skipcnt_5,
            ltout => OPEN,
            carryin => n19614,
            carryout => n19615,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i6_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38426\,
            in2 => \_gnd_net_\,
            in3 => \N__32520\,
            lcout => acadc_skipcnt_6,
            ltout => OPEN,
            carryin => n19615,
            carryout => n19616,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i7_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41597\,
            in2 => \_gnd_net_\,
            in3 => \N__32517\,
            lcout => acadc_skipcnt_7,
            ltout => OPEN,
            carryin => n19616,
            carryout => n19617,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i8_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32513\,
            in2 => \_gnd_net_\,
            in3 => \N__32499\,
            lcout => acadc_skipcnt_8,
            ltout => OPEN,
            carryin => n19617,
            carryout => n19618,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32658\,
            sr => \N__32622\
        );

    \acadc_skipcnt_i0_i9_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32495\,
            in2 => \_gnd_net_\,
            in3 => \N__32481\,
            lcout => acadc_skipcnt_9,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => n19619,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32657\,
            sr => \N__32618\
        );

    \acadc_skipcnt_i0_i10_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32474\,
            in2 => \_gnd_net_\,
            in3 => \N__32460\,
            lcout => acadc_skipcnt_10,
            ltout => OPEN,
            carryin => n19619,
            carryout => n19620,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32657\,
            sr => \N__32618\
        );

    \acadc_skipcnt_i0_i11_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32456\,
            in2 => \_gnd_net_\,
            in3 => \N__32442\,
            lcout => acadc_skipcnt_11,
            ltout => OPEN,
            carryin => n19620,
            carryout => n19621,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32657\,
            sr => \N__32618\
        );

    \acadc_skipcnt_i0_i12_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32435\,
            in2 => \_gnd_net_\,
            in3 => \N__32421\,
            lcout => acadc_skipcnt_12,
            ltout => OPEN,
            carryin => n19621,
            carryout => n19622,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32657\,
            sr => \N__32618\
        );

    \acadc_skipcnt_i0_i13_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32711\,
            in2 => \_gnd_net_\,
            in3 => \N__32697\,
            lcout => acadc_skipcnt_13,
            ltout => OPEN,
            carryin => n19622,
            carryout => n19623,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32657\,
            sr => \N__32618\
        );

    \acadc_skipcnt_i0_i14_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32693\,
            in2 => \_gnd_net_\,
            in3 => \N__32679\,
            lcout => acadc_skipcnt_14,
            ltout => OPEN,
            carryin => n19623,
            carryout => n19624,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32657\,
            sr => \N__32618\
        );

    \acadc_skipcnt_i0_i15_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32672\,
            in2 => \_gnd_net_\,
            in3 => \N__32676\,
            lcout => acadc_skipcnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32657\,
            sr => \N__32618\
        );

    \ADC_VDC.i19363_4_lut_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110111"
        )
    port map (
            in0 => \N__48481\,
            in1 => \N__32567\,
            in2 => \N__48835\,
            in3 => \N__34338\,
            lcout => \ADC_VDC.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i2_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__48758\,
            in1 => \N__48277\,
            in2 => \_gnd_net_\,
            in3 => \N__47359\,
            lcout => adc_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53261\,
            ce => \N__32598\,
            sr => \N__32589\
        );

    \ADC_VDC.i19412_4_lut_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__48480\,
            in1 => \N__32577\,
            in2 => \N__48773\,
            in3 => \N__47480\,
            lcout => \ADC_VDC.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i2_2_lut_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48275\,
            in2 => \_gnd_net_\,
            in3 => \N__47358\,
            lcout => \ADC_VDC.n7_adj_1398\,
            ltout => \ADC_VDC.n7_adj_1398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_11_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32571\,
            in3 => \N__47481\,
            lcout => \ADC_VDC.n77\,
            ltout => \ADC_VDC.n77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_16_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101110"
        )
    port map (
            in0 => \N__48754\,
            in1 => \N__48479\,
            in2 => \N__32787\,
            in3 => \N__32784\,
            lcout => OPEN,
            ltout => \ADC_VDC.n72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_17_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__48276\,
            in1 => \N__32778\,
            in2 => \N__32772\,
            in3 => \N__34806\,
            lcout => \ADC_VDC.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i37_4_lut_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101001010010"
        )
    port map (
            in0 => \N__47334\,
            in1 => \N__48288\,
            in2 => \N__47491\,
            in3 => \N__32904\,
            lcout => OPEN,
            ltout => \ADC_VDC.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_13_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__48455\,
            in1 => \N__48774\,
            in2 => \N__32769\,
            in3 => \N__34323\,
            lcout => \ADC_VDC.n20811\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110001101100"
        )
    port map (
            in0 => \N__47333\,
            in1 => \N__48287\,
            in2 => \N__48844\,
            in3 => \N__32726\,
            lcout => OPEN,
            ltout => \ADC_VDC.n22195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.n22195_bdd_4_lut_4_lut_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010011110100"
        )
    port map (
            in0 => \N__48709\,
            in1 => \N__34329\,
            in2 => \N__32766\,
            in3 => \N__47335\,
            lcout => OPEN,
            ltout => \ADC_VDC.n22198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i1_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48778\,
            in1 => \N__48456\,
            in2 => \N__32763\,
            in3 => \N__32760\,
            lcout => \ADC_VDC.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53265\,
            ce => \N__32745\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_14_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36708\,
            in2 => \_gnd_net_\,
            in3 => \N__34845\,
            lcout => OPEN,
            ltout => \ADC_VDC.n6_adj_1399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_adj_15_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__36920\,
            in1 => \N__36611\,
            in2 => \N__32736\,
            in3 => \N__36645\,
            lcout => \ADC_VDC.n10536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18983_4_lut_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__36612\,
            in1 => \N__36921\,
            in2 => \N__48529\,
            in3 => \N__34311\,
            lcout => \ADC_VDC.n21229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i0_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110110"
        )
    port map (
            in0 => \N__48784\,
            in1 => \N__48530\,
            in2 => \N__47489\,
            in3 => \N__47357\,
            lcout => \ADC_VDC.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53207\,
            ce => \N__32898\,
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i7_12189_12190_reset_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37344\,
            in1 => \N__44445\,
            in2 => \_gnd_net_\,
            in3 => \N__42387\,
            lcout => \comm_spi.n14608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__35108\
        );

    \comm_buf_2__i1_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45725\,
            in1 => \N__32802\,
            in2 => \_gnd_net_\,
            in3 => \N__51800\,
            lcout => comm_buf_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54274\,
            ce => \N__33093\,
            sr => \N__33071\
        );

    \mux_130_Mux_1_i19_3_lut_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__57757\,
            in1 => \_gnd_net_\,
            in2 => \N__32871\,
            in3 => \N__33713\,
            lcout => OPEN,
            ltout => \n19_adj_1491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i22_3_lut_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32846\,
            in2 => \N__32823\,
            in3 => \N__53720\,
            lcout => OPEN,
            ltout => \n22_adj_1488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i30_3_lut_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__54707\,
            in1 => \N__32820\,
            in2 => \N__32805\,
            in3 => \_gnd_net_\,
            lcout => n30_adj_1506,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19734_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__32796\,
            in1 => \N__50658\,
            in2 => \N__45684\,
            in3 => \N__52331\,
            lcout => OPEN,
            ltout => \n22249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22249_bdd_4_lut_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52332\,
            in1 => \N__40145\,
            in2 => \N__32790\,
            in3 => \N__37447\,
            lcout => n22252,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19739_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__32967\,
            in1 => \N__50657\,
            in2 => \N__45504\,
            in3 => \N__52330\,
            lcout => n22381,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i0_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32994\,
            in1 => \N__51868\,
            in2 => \_gnd_net_\,
            in3 => \N__53038\,
            lcout => comm_buf_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54278\,
            ce => \N__33092\,
            sr => \N__33072\
        );

    \comm_buf_2__i7_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51867\,
            in1 => \N__50349\,
            in2 => \_gnd_net_\,
            in3 => \N__32982\,
            lcout => comm_buf_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54278\,
            ce => \N__33092\,
            sr => \N__33072\
        );

    \comm_buf_2__i6_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46405\,
            in1 => \N__32961\,
            in2 => \_gnd_net_\,
            in3 => \N__51871\,
            lcout => comm_buf_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54278\,
            ce => \N__33092\,
            sr => \N__33072\
        );

    \comm_buf_2__i5_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51866\,
            in1 => \N__52059\,
            in2 => \_gnd_net_\,
            in3 => \N__32946\,
            lcout => comm_buf_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54278\,
            ce => \N__33092\,
            sr => \N__33072\
        );

    \comm_buf_2__i4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46730\,
            in1 => \N__32934\,
            in2 => \_gnd_net_\,
            in3 => \N__51870\,
            lcout => comm_buf_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54278\,
            ce => \N__33092\,
            sr => \N__33072\
        );

    \comm_buf_2__i3_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51865\,
            in1 => \N__51055\,
            in2 => \_gnd_net_\,
            in3 => \N__32925\,
            lcout => comm_buf_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54278\,
            ce => \N__33092\,
            sr => \N__33072\
        );

    \comm_buf_2__i2_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32916\,
            in1 => \N__47175\,
            in2 => \_gnd_net_\,
            in3 => \N__51869\,
            lcout => comm_buf_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54278\,
            ce => \N__33092\,
            sr => \N__33072\
        );

    \mux_137_Mux_3_i4_3_lut_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39861\,
            in1 => \N__50669\,
            in2 => \_gnd_net_\,
            in3 => \N__42576\,
            lcout => OPEN,
            ltout => \n4_adj_1594_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18583_4_lut_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__52344\,
            in1 => \N__33780\,
            in2 => \N__32907\,
            in3 => \N__50688\,
            lcout => n21193,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19744_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__33024\,
            in1 => \N__50668\,
            in2 => \N__45435\,
            in3 => \N__52345\,
            lcout => OPEN,
            ltout => \n22387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22387_bdd_4_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52346\,
            in1 => \N__44222\,
            in2 => \N__33018\,
            in3 => \N__51012\,
            lcout => OPEN,
            ltout => \n22390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i3_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33015\,
            in2 => \N__33009\,
            in3 => \N__50538\,
            lcout => comm_tx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54281\,
            ce => \N__45234\,
            sr => \N__45172\
        );

    \mux_137_Mux_7_i4_3_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50670\,
            in1 => \N__39942\,
            in2 => \_gnd_net_\,
            in3 => \N__42675\,
            lcout => OPEN,
            ltout => \n4_adj_1587_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18565_4_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__33047\,
            in1 => \N__50671\,
            in2 => \N__33006\,
            in3 => \N__52347\,
            lcout => OPEN,
            ltout => \n21175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i7_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50539\,
            in1 => \_gnd_net_\,
            in2 => \N__33003\,
            in3 => \N__34221\,
            lcout => comm_tx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54281\,
            ce => \N__45234\,
            sr => \N__45172\
        );

    \i458_2_lut_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50038\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49846\,
            lcout => n2358,
            ltout => \n2358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_255_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__50753\,
            in1 => \N__52370\,
            in2 => \N__33000\,
            in3 => \N__52266\,
            lcout => n20850,
            ltout => \n20850_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i36_4_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__51799\,
            in1 => \N__45636\,
            in2 => \N__32997\,
            in3 => \N__33894\,
            lcout => OPEN,
            ltout => \n31_adj_1613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_270_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45927\,
            in2 => \N__33096\,
            in3 => \N__45881\,
            lcout => n12085,
            ltout => \n12085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12351_2_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__56863\,
            in1 => \_gnd_net_\,
            in2 => \N__33075\,
            in3 => \_gnd_net_\,
            lcout => n14764,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_214_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__49586\,
            in1 => \N__33030\,
            in2 => \_gnd_net_\,
            in3 => \N__56864\,
            lcout => n12228,
            ltout => \n12228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i7_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__56865\,
            in1 => \N__50380\,
            in2 => \N__33051\,
            in3 => \N__33048\,
            lcout => comm_buf_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i6_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__45593\,
            in1 => \N__56866\,
            in2 => \N__46448\,
            in3 => \N__34993\,
            lcout => comm_buf_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_213_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51792\,
            in1 => \N__33036\,
            in2 => \N__37671\,
            in3 => \N__55518\,
            lcout => n20852,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i4_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__46000\,
            in1 => \N__46071\,
            in2 => \N__46755\,
            in3 => \N__49776\,
            lcout => comm_cmd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i0_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__57388\,
            in1 => \N__53040\,
            in2 => \N__46082\,
            in3 => \N__45999\,
            lcout => comm_cmd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_104_2_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34897\,
            lcout => \comm_spi.data_tx_7__N_786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i5_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__34996\,
            in1 => \N__52092\,
            in2 => \N__57088\,
            in3 => \N__42446\,
            lcout => comm_buf_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i0_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__53039\,
            in1 => \N__56992\,
            in2 => \N__42317\,
            in3 => \N__34994\,
            lcout => comm_buf_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i3_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__34995\,
            in1 => \N__51071\,
            in2 => \N__57087\,
            in3 => \N__33776\,
            lcout => comm_buf_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i38_3_lut_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__54868\,
            in1 => \N__57387\,
            in2 => \_gnd_net_\,
            in3 => \N__53489\,
            lcout => n22_adj_1615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i1_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__44934\,
            in1 => \N__37440\,
            in2 => \N__40656\,
            in3 => \N__33758\,
            lcout => buf_dds1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33458\,
            in1 => \N__33678\,
            in2 => \N__33709\,
            in3 => \N__33738\,
            lcout => buf_adcdata_vac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i10_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33677\,
            in1 => \N__33459\,
            in2 => \N__35954\,
            in3 => \N__33128\,
            lcout => buf_adcdata_vac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i1_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__46001\,
            in1 => \N__46070\,
            in2 => \N__45794\,
            in3 => \N__54837\,
            lcout => comm_cmd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__54836\,
            in1 => \N__57262\,
            in2 => \_gnd_net_\,
            in3 => \N__53458\,
            lcout => n9_adj_1416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i0_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__33923\,
            in1 => \N__40631\,
            in2 => \N__43299\,
            in3 => \N__44935\,
            lcout => buf_dds1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__54835\,
            in1 => \N__57261\,
            in2 => \_gnd_net_\,
            in3 => \N__53457\,
            lcout => n10717,
            ltout => \n10717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19112_4_lut_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__49271\,
            in1 => \N__33903\,
            in2 => \N__33897\,
            in3 => \N__54569\,
            lcout => n21344,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i5_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__44931\,
            in1 => \N__33883\,
            in2 => \N__37496\,
            in3 => \N__57049\,
            lcout => buf_dds1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i3_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__46012\,
            in1 => \N__46079\,
            in2 => \N__51106\,
            in3 => \N__54601\,
            lcout => comm_cmd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i7_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__44932\,
            in1 => \N__33847\,
            in2 => \N__50321\,
            in3 => \N__40637\,
            lcout => buf_dds1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_6_i23_3_lut_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57589\,
            in1 => \N__38674\,
            in2 => \_gnd_net_\,
            in3 => \N__33828\,
            lcout => n23_adj_1538,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i16_3_lut_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33988\,
            in1 => \N__33807\,
            in2 => \_gnd_net_\,
            in3 => \N__57588\,
            lcout => n16_adj_1510,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i8_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41741\,
            in1 => \N__37851\,
            in2 => \_gnd_net_\,
            in3 => \N__43876\,
            lcout => req_data_cnt_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i6_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47832\,
            in1 => \N__41740\,
            in2 => \_gnd_net_\,
            in3 => \N__40781\,
            lcout => req_data_cnt_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i4_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__33992\,
            in1 => \N__40635\,
            in2 => \N__47784\,
            in3 => \N__44933\,
            lcout => buf_dds1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_284_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__49786\,
            in1 => \N__49732\,
            in2 => \N__49496\,
            in3 => \N__49696\,
            lcout => n20804,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i6_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__49733\,
            in1 => \N__46013\,
            in2 => \N__46464\,
            in3 => \N__46080\,
            lcout => comm_cmd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i3_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56474\,
            in1 => \N__44325\,
            in2 => \N__51020\,
            in3 => \N__50080\,
            lcout => \acadc_skipCount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i0_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__43290\,
            in1 => \N__56475\,
            in2 => \N__33972\,
            in3 => \N__48012\,
            lcout => buf_dds0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15337_2_lut_3_lut_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__55548\,
            in1 => \_gnd_net_\,
            in2 => \N__41491\,
            in3 => \N__51880\,
            lcout => n14_adj_1577,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_184_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__38127\,
            in1 => \N__41049\,
            in2 => \N__43877\,
            in3 => \N__33940\,
            lcout => n19_adj_1607,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i2_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37547\,
            in1 => \N__41729\,
            in2 => \_gnd_net_\,
            in3 => \N__46607\,
            lcout => req_data_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_312_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__49695\,
            in1 => \N__49777\,
            in2 => \_gnd_net_\,
            in3 => \N__49731\,
            lcout => n20893,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i9_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37827\,
            in1 => \N__41730\,
            in2 => \_gnd_net_\,
            in3 => \N__34265\,
            lcout => req_data_cnt_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_264_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34112\,
            in2 => \_gnd_net_\,
            in3 => \N__41764\,
            lcout => n10697,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34053\,
            in1 => \N__36066\,
            in2 => \N__36009\,
            in3 => \N__34122\,
            lcout => OPEN,
            ltout => \n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_198_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34284\,
            in2 => \N__34044\,
            in3 => \N__34005\,
            lcout => n16_adj_1603,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_stop_328_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34285\,
            in1 => \N__40135\,
            in2 => \_gnd_net_\,
            in3 => \N__36247\,
            lcout => eis_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_173_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__38088\,
            in1 => \N__41175\,
            in2 => \N__36230\,
            in3 => \N__34261\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_178_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__38148\,
            in1 => \N__41229\,
            in2 => \N__40820\,
            in3 => \N__34087\,
            lcout => OPEN,
            ltout => \n21_adj_1492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_187_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36039\,
            in1 => \N__34014\,
            in2 => \N__34008\,
            in3 => \N__36072\,
            lcout => n30_adj_1618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19084_2_lut_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57554\,
            in2 => \_gnd_net_\,
            in3 => \N__34088\,
            lcout => n21309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_306_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111101"
        )
    port map (
            in0 => \N__54602\,
            in1 => \N__37644\,
            in2 => \N__49495\,
            in3 => \_gnd_net_\,
            lcout => n20907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_179_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__50862\,
            in1 => \N__51155\,
            in2 => \N__50113\,
            in3 => \N__52840\,
            lcout => n20_adj_1617,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__41762\,
            in1 => \N__55542\,
            in2 => \N__51958\,
            in3 => \N__34111\,
            lcout => n10598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i12_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41699\,
            in1 => \N__37769\,
            in2 => \_gnd_net_\,
            in3 => \N__34089\,
            lcout => req_data_cnt_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i1_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37589\,
            in1 => \N__41700\,
            in2 => \_gnd_net_\,
            in3 => \N__37085\,
            lcout => req_data_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i3_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41701\,
            in1 => \_gnd_net_\,
            in2 => \N__50117\,
            in3 => \N__47096\,
            lcout => req_data_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22375_bdd_4_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__34245\,
            in1 => \N__55022\,
            in2 => \N__36366\,
            in3 => \N__34072\,
            lcout => n22378,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_263_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__56400\,
            in1 => \N__57126\,
            in2 => \N__44409\,
            in3 => \N__41763\,
            lcout => n12399,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15347_2_lut_3_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__51876\,
            in1 => \N__55543\,
            in2 => \_gnd_net_\,
            in3 => \N__43815\,
            lcout => n14_adj_1550,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15339_2_lut_3_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__55544\,
            in1 => \N__44749\,
            in2 => \_gnd_net_\,
            in3 => \N__51877\,
            lcout => n14_adj_1579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6449_3_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37424\,
            in1 => \N__36288\,
            in2 => \_gnd_net_\,
            in3 => \N__47683\,
            lcout => n8_adj_1573,
            ltout => \n8_adj_1573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__57133\,
            in1 => \N__56512\,
            in2 => \N__34299\,
            in3 => \N__36477\,
            lcout => data_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19754_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__57553\,
            in1 => \N__34295\,
            in2 => \N__55146\,
            in3 => \N__34266\,
            lcout => n22375,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22381_bdd_4_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__50318\,
            in1 => \N__52413\,
            in2 => \N__34239\,
            in3 => \N__42802\,
            lcout => n22384,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds0_304_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__42124\,
            in1 => \N__34206\,
            in2 => \N__56556\,
            in3 => \N__57134\,
            lcout => trig_dds0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.SCLK_27_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011101101"
        )
    port map (
            in0 => \N__42958\,
            in1 => \N__34178\,
            in2 => \N__41336\,
            in3 => \N__42189\,
            lcout => \DDS_SCK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i23_4_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110011001"
        )
    port map (
            in0 => \N__42188\,
            in1 => \N__42956\,
            in2 => \N__42120\,
            in3 => \N__41327\,
            lcout => \SIG_DDS.n9_adj_1393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i2_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__42957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42190\,
            lcout => dds_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i1_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41337\,
            in2 => \_gnd_net_\,
            in3 => \N__42197\,
            lcout => dds_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54413\,
            ce => \N__36096\,
            sr => \N__43060\
        );

    \comm_spi.i12188_3_lut_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34167\,
            in1 => \N__34155\,
            in2 => \_gnd_net_\,
            in3 => \N__35165\,
            lcout => \ICE_SPI_MISO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i40_3_lut_4_lut_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101101000011"
        )
    port map (
            in0 => \N__48298\,
            in1 => \N__47377\,
            in2 => \N__47492\,
            in3 => \N__34826\,
            lcout => \ADC_VDC.n19_adj_1401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19327_4_lut_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__36639\,
            in1 => \N__36604\,
            in2 => \N__36707\,
            in3 => \N__36668\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19100_4_lut_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__36912\,
            in1 => \N__34305\,
            in2 => \N__34332\,
            in3 => \N__47332\,
            lcout => \ADC_VDC.n21320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18357_2_lut_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47482\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48300\,
            lcout => \ADC_VDC.n20965\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_2_lut_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__42495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55810\,
            lcout => \comm_spi.data_tx_7__N_795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_adj_12_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__36638\,
            in1 => \N__36879\,
            in2 => \N__36706\,
            in3 => \N__36667\,
            lcout => OPEN,
            ltout => \ADC_VDC.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i5_3_lut_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36826\,
            in2 => \N__34314\,
            in3 => \N__36853\,
            lcout => \ADC_VDC.n20812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i2_3_lut_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__36854\,
            in1 => \N__36880\,
            in2 => \_gnd_net_\,
            in3 => \N__36827\,
            lcout => \ADC_VDC.n20784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__47348\,
            in1 => \N__48536\,
            in2 => \N__34854\,
            in3 => \N__48219\,
            lcout => \ADC_VDC.n18550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_9_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36603\,
            in2 => \_gnd_net_\,
            in3 => \N__36640\,
            lcout => \ADC_VDC.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i15111_2_lut_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48792\,
            in2 => \_gnd_net_\,
            in3 => \N__48297\,
            lcout => \ADC_VDC.n17509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_4_lut_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36825\,
            in1 => \N__36852\,
            in2 => \N__36882\,
            in3 => \N__36666\,
            lcout => \ADC_VDC.n11265\,
            ltout => \ADC_VDC.n11265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__36919\,
            in1 => \N__34839\,
            in2 => \N__34833\,
            in3 => \N__36704\,
            lcout => \ADC_VDC.n15\,
            ltout => \ADC_VDC.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18386_2_lut_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34809\,
            in3 => \N__47347\,
            lcout => \ADC_VDC.n20996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i19328_4_lut_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100111001100"
        )
    port map (
            in0 => \N__34771\,
            in1 => \N__34620\,
            in2 => \N__44059\,
            in3 => \N__34464\,
            lcout => \CLK_DDS.n12784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i7_12189_12190_set_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37343\,
            in1 => \N__44441\,
            in2 => \_gnd_net_\,
            in3 => \N__42386\,
            lcout => \comm_spi.n14607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52547\,
            ce => 'H',
            sr => \N__35044\
        );

    \comm_clear_301_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__56958\,
            in1 => \N__51761\,
            in2 => \_gnd_net_\,
            in3 => \N__49489\,
            lcout => comm_clear,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54279\,
            ce => \N__34866\,
            sr => \_gnd_net_\
        );

    \comm_index_i1_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100100000"
        )
    port map (
            in0 => \N__49876\,
            in1 => \N__49965\,
            in2 => \N__50780\,
            in3 => \N__52355\,
            lcout => comm_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54282\,
            ce => \N__36030\,
            sr => \N__39429\
        );

    \comm_index_i0_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__49964\,
            in1 => \N__50733\,
            in2 => \_gnd_net_\,
            in3 => \N__49875\,
            lcout => comm_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54282\,
            ce => \N__36030\,
            sr => \N__39429\
        );

    \comm_index_i2_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__50578\,
            in1 => \N__52354\,
            in2 => \N__50781\,
            in3 => \N__49087\,
            lcout => comm_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54282\,
            ce => \N__36030\,
            sr => \N__39429\
        );

    \i18512_4_lut_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__49171\,
            in1 => \N__52212\,
            in2 => \N__34875\,
            in3 => \N__55407\,
            lcout => OPEN,
            ltout => \n21122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i0_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__56826\,
            in1 => \_gnd_net_\,
            in2 => \N__34878\,
            in3 => \N__56544\,
            lcout => comm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54290\,
            ce => \N__36981\,
            sr => \_gnd_net_\
        );

    \i18510_3_lut_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010101"
        )
    port map (
            in0 => \N__49407\,
            in1 => \N__50008\,
            in2 => \_gnd_net_\,
            in3 => \N__51644\,
            lcout => n21120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_313_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__50012\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49404\,
            lcout => n14529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_adj_271_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__49406\,
            in1 => \N__51643\,
            in2 => \_gnd_net_\,
            in3 => \N__56825\,
            lcout => n11361,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i22_4_lut_4_lut_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001000"
        )
    port map (
            in0 => \N__51642\,
            in1 => \N__49849\,
            in2 => \N__50037\,
            in3 => \N__49405\,
            lcout => OPEN,
            ltout => \n7_adj_1616_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_219_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__49562\,
            in1 => \N__55406\,
            in2 => \N__34857\,
            in3 => \N__56824\,
            lcout => n11896,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_valid_85_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__35898\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35853\,
            lcout => comm_data_vld,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.data_valid_85C_net\,
            ce => 'H',
            sr => \N__55820\
        );

    \ADC_IAC.ADC_DATA_i13_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35807\,
            in1 => \N__35637\,
            in2 => \N__35250\,
            in3 => \N__53813\,
            lcout => buf_adcdata_iac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18514_4_lut_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__57385\,
            in1 => \N__35214\,
            in2 => \N__37698\,
            in3 => \N__54884\,
            lcout => n21124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19425_4_lut_3_lut_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35146\,
            in1 => \N__35065\,
            in2 => \_gnd_net_\,
            in3 => \N__55817\,
            lcout => \comm_spi.n14603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_100_2_lut_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55816\,
            in2 => \_gnd_net_\,
            in3 => \N__35067\,
            lcout => \comm_spi.data_tx_7__N_774\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_92_2_lut_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35066\,
            in2 => \_gnd_net_\,
            in3 => \N__55818\,
            lcout => \comm_spi.data_tx_7__N_766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i1_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__39638\,
            in1 => \N__56831\,
            in2 => \N__45791\,
            in3 => \N__34997\,
            lcout => comm_buf_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i19_3_lut_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34968\,
            in1 => \N__34937\,
            in2 => \_gnd_net_\,
            in3 => \N__57386\,
            lcout => n19_adj_1522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19445_4_lut_3_lut_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55819\,
            in1 => \N__39118\,
            in2 => \_gnd_net_\,
            in3 => \N__34901\,
            lcout => \comm_spi.n22875\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i2_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__44908\,
            in1 => \N__48084\,
            in2 => \N__46891\,
            in3 => \N__40636\,
            lcout => buf_dds1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_51_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__55522\,
            in1 => \N__51858\,
            in2 => \N__57109\,
            in3 => \N__44907\,
            lcout => n16891,
            ltout => \n16891_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i9_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__44909\,
            in1 => \N__40119\,
            in2 => \N__36000\,
            in3 => \N__40237\,
            lcout => buf_dds1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19009_2_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43188\,
            in2 => \_gnd_net_\,
            in3 => \N__42286\,
            lcout => \SIG_DDS.n21571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i19_3_lut_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35982\,
            in1 => \N__35947\,
            in2 => \_gnd_net_\,
            in3 => \N__57499\,
            lcout => n19_adj_1518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i2_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__46078\,
            in1 => \N__45998\,
            in2 => \N__47224\,
            in3 => \N__53670\,
            lcout => comm_cmd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_response_302_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100110000"
        )
    port map (
            in0 => \N__49485\,
            in1 => \N__55525\,
            in2 => \N__57028\,
            in3 => \N__51826\,
            lcout => \ICE_GPMI_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54333\,
            ce => \N__35907\,
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_292_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010000"
        )
    port map (
            in0 => \N__55524\,
            in1 => \N__56901\,
            in2 => \N__49591\,
            in3 => \N__49484\,
            lcout => n11385,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i17_3_lut_3_lut_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__49483\,
            in1 => \N__55523\,
            in2 => \_gnd_net_\,
            in3 => \N__51825\,
            lcout => OPEN,
            ltout => \n10_adj_1554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_261_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__49575\,
            in1 => \_gnd_net_\,
            in2 => \N__36033\,
            in3 => \N__56900\,
            lcout => n11850,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_241_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__54913\,
            in1 => \N__57498\,
            in2 => \N__41532\,
            in3 => \N__53548\,
            lcout => n20914,
            ltout => \n20914_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_226_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100011"
        )
    port map (
            in0 => \N__49574\,
            in1 => \N__36015\,
            in2 => \N__36018\,
            in3 => \N__56899\,
            lcout => n11819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18404_2_lut_3_lut_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__51824\,
            in1 => \N__55500\,
            in2 => \_gnd_net_\,
            in3 => \N__49482\,
            lcout => n21014,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i0_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__41723\,
            in1 => \N__37614\,
            in2 => \N__43334\,
            in3 => \_gnd_net_\,
            lcout => req_data_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15327_2_lut_3_lut_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__55550\,
            in1 => \N__51428\,
            in2 => \_gnd_net_\,
            in3 => \N__51862\,
            lcout => n14_adj_1584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_186_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__46511\,
            in1 => \N__43391\,
            in2 => \N__43333\,
            in3 => \N__40777\,
            lcout => n17_adj_1489,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15344_2_lut_3_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__55551\,
            in1 => \N__48068\,
            in2 => \_gnd_net_\,
            in3 => \N__51863\,
            lcout => n14_adj_1555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_251_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__54554\,
            in1 => \N__49481\,
            in2 => \_gnd_net_\,
            in3 => \N__37645\,
            lcout => n20912,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15346_2_lut_3_lut_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__55549\,
            in1 => \N__42770\,
            in2 => \_gnd_net_\,
            in3 => \N__51861\,
            lcout => n14_adj_1549,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i5_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__46081\,
            in1 => \N__46008\,
            in2 => \N__52125\,
            in3 => \N__49700\,
            lcout => comm_cmd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15385_2_lut_3_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__55552\,
            in1 => \N__43292\,
            in2 => \_gnd_net_\,
            in3 => \N__51864\,
            lcout => n14_adj_1533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i12_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__40309\,
            in1 => \N__40655\,
            in2 => \N__41492\,
            in3 => \N__44947\,
            lcout => buf_dds1_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19064_2_lut_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57661\,
            in2 => \_gnd_net_\,
            in3 => \N__36055\,
            lcout => n21286,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i14_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36056\,
            in1 => \N__38070\,
            in2 => \_gnd_net_\,
            in3 => \N__41725\,
            lcout => req_data_cnt_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19372_4_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__42131\,
            in1 => \N__41311\,
            in2 => \N__43059\,
            in3 => \N__42266\,
            lcout => \SIG_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i7_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46993\,
            in2 => \N__41739\,
            in3 => \N__37878\,
            lcout => req_data_cnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_174_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__47122\,
            in1 => \N__50452\,
            in2 => \N__46997\,
            in3 => \N__46603\,
            lcout => n22_adj_1499,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_182_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__37918\,
            in1 => \N__46192\,
            in2 => \N__46817\,
            in3 => \N__37081\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_177_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__38105\,
            in1 => \N__40936\,
            in2 => \N__36060\,
            in3 => \N__41020\,
            lcout => n23_adj_1614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i10_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37790\,
            in1 => \N__41702\,
            in2 => \_gnd_net_\,
            in3 => \N__40813\,
            lcout => req_data_cnt_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i11_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41703\,
            in1 => \N__44427\,
            in2 => \_gnd_net_\,
            in3 => \N__41021\,
            lcout => req_data_cnt_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_130_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__49426\,
            in1 => \N__47058\,
            in2 => \N__57108\,
            in3 => \N__36333\,
            lcout => n10520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i4_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37526\,
            in2 => \N__41724\,
            in3 => \N__46813\,
            lcout => req_data_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i15_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38028\,
            in1 => \N__41704\,
            in2 => \_gnd_net_\,
            in3 => \N__36223\,
            lcout => req_data_cnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_267_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__47690\,
            in1 => \N__57014\,
            in2 => \N__36558\,
            in3 => \N__56228\,
            lcout => n12280,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4408_3_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43283\,
            in1 => \N__36321\,
            in2 => \_gnd_net_\,
            in3 => \N__47689\,
            lcout => n8_adj_1532,
            ltout => \n8_adj_1532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__36302\,
            in1 => \N__56227\,
            in2 => \N__36204\,
            in3 => \N__57013\,
            lcout => \data_index_9_N_216_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i0_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__57015\,
            in1 => \N__36303\,
            in2 => \N__56344\,
            in3 => \N__36102\,
            lcout => data_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_310_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__57654\,
            in1 => \N__54747\,
            in2 => \_gnd_net_\,
            in3 => \N__37652\,
            lcout => n11338,
            ltout => \n11338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__49425\,
            in1 => \N__55056\,
            in2 => \N__36327\,
            in3 => \N__53679\,
            lcout => n8813,
            ltout => \n8813_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6429_3_lut_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51019\,
            in2 => \N__36324\,
            in3 => \N__41099\,
            lcout => n8_adj_1569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i5_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37497\,
            in1 => \N__41698\,
            in2 => \_gnd_net_\,
            in3 => \N__52844\,
            lcout => req_data_cnt_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_2_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36320\,
            in1 => \N__36319\,
            in2 => \N__36536\,
            in3 => \N__36291\,
            lcout => n7,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => n19625,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_3_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36287\,
            in1 => \N__36286\,
            in2 => \N__36559\,
            in3 => \N__36270\,
            lcout => n7_adj_1572,
            ltout => OPEN,
            carryin => n19625,
            carryout => n19626,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_4_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41004\,
            in1 => \N__41003\,
            in2 => \N__36537\,
            in3 => \N__36267\,
            lcout => n7_adj_1570,
            ltout => OPEN,
            carryin => n19626,
            carryout => n19627,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_5_lut_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41100\,
            in1 => \N__41098\,
            in2 => \N__36560\,
            in3 => \N__36264\,
            lcout => n7_adj_1568,
            ltout => OPEN,
            carryin => n19627,
            carryout => n19628,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_6_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47723\,
            in1 => \N__47722\,
            in2 => \N__36538\,
            in3 => \N__36261\,
            lcout => n7_adj_1566,
            ltout => OPEN,
            carryin => n19628,
            carryout => n19629,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_7_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__40569\,
            in1 => \N__40567\,
            in2 => \N__36561\,
            in3 => \N__36579\,
            lcout => n17487,
            ltout => OPEN,
            carryin => n19629,
            carryout => n19630,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_8_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38393\,
            in1 => \N__38392\,
            in2 => \N__36539\,
            in3 => \N__36576\,
            lcout => n7_adj_1564,
            ltout => OPEN,
            carryin => n19630,
            carryout => n19631,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_9_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41991\,
            in1 => \N__41990\,
            in2 => \N__36562\,
            in3 => \N__36573\,
            lcout => n7_adj_1562,
            ltout => OPEN,
            carryin => n19631,
            carryout => n19632,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_10_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42062\,
            in1 => \N__42058\,
            in2 => \N__36567\,
            in3 => \N__36570\,
            lcout => n7_adj_1560,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => n19633,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_11_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39076\,
            in1 => \N__39077\,
            in2 => \N__36566\,
            in3 => \N__36480\,
            lcout => n7_adj_1558,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i8_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__57059\,
            in1 => \N__42042\,
            in2 => \N__56473\,
            in3 => \N__38952\,
            lcout => data_index_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i3_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56357\,
            in1 => \N__41887\,
            in2 => \N__44228\,
            in3 => \N__41953\,
            lcout => \SELIRNG1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__36476\,
            in1 => \N__57090\,
            in2 => \N__56472\,
            in3 => \N__36465\,
            lcout => \data_index_9_N_216_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i1_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56356\,
            in1 => \N__41886\,
            in2 => \N__40155\,
            in3 => \N__36352\,
            lcout => \DDS_RNG_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.MOSI_31_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36780\,
            in1 => \N__36752\,
            in2 => \_gnd_net_\,
            in3 => \N__42976\,
            lcout => \DDS_MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i9_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__39060\,
            in1 => \N__57060\,
            in2 => \N__56476\,
            in3 => \N__39054\,
            lcout => data_index_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.CS_28_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__42196\,
            in1 => \N__42983\,
            in2 => \_gnd_net_\,
            in3 => \N__41335\,
            lcout => \DDS_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54421\,
            ce => \N__36720\,
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i2_12204_12205_reset_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39344\,
            in1 => \N__38573\,
            in2 => \_gnd_net_\,
            in3 => \N__38618\,
            lcout => \comm_spi.n14623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52641\,
            ce => 'H',
            sr => \N__39321\
        );

    \comm_spi.data_tx_i0_12174_12175_reset_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__58335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52639\,
            ce => 'H',
            sr => \N__36714\
        );

    \ADC_VDC.bit_cnt_3769__i0_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36705\,
            in2 => \_gnd_net_\,
            in3 => \N__36672\,
            lcout => \ADC_VDC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \ADC_VDC.n19772\,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \ADC_VDC.bit_cnt_3769__i1_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36669\,
            in2 => \_gnd_net_\,
            in3 => \N__36648\,
            lcout => \ADC_VDC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19772\,
            carryout => \ADC_VDC.n19773\,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \ADC_VDC.bit_cnt_3769__i2_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36644\,
            in2 => \_gnd_net_\,
            in3 => \N__36615\,
            lcout => \ADC_VDC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19773\,
            carryout => \ADC_VDC.n19774\,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \ADC_VDC.bit_cnt_3769__i3_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36610\,
            in2 => \_gnd_net_\,
            in3 => \N__36582\,
            lcout => \ADC_VDC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19774\,
            carryout => \ADC_VDC.n19775\,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \ADC_VDC.bit_cnt_3769__i4_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36913\,
            in2 => \_gnd_net_\,
            in3 => \N__36885\,
            lcout => \ADC_VDC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19775\,
            carryout => \ADC_VDC.n19776\,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \ADC_VDC.bit_cnt_3769__i5_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36881\,
            in2 => \_gnd_net_\,
            in3 => \N__36858\,
            lcout => \ADC_VDC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19776\,
            carryout => \ADC_VDC.n19777\,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \ADC_VDC.bit_cnt_3769__i6_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36855\,
            in2 => \_gnd_net_\,
            in3 => \N__36834\,
            lcout => \ADC_VDC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19777\,
            carryout => \ADC_VDC.n19778\,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \ADC_VDC.bit_cnt_3769__i7_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36828\,
            in2 => \_gnd_net_\,
            in3 => \N__36831\,
            lcout => \ADC_VDC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53194\,
            ce => \N__47508\,
            sr => \N__36804\
        );

    \wdtick_flag_289_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__39245\,
            in1 => \N__39225\,
            in2 => \N__39264\,
            in3 => \N__44633\,
            lcout => wdtick_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39205\,
            ce => 'H',
            sr => \N__39417\
        );

    \comm_spi.data_tx_i4_12212_12213_reset_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39131\,
            in1 => \N__39095\,
            in2 => \_gnd_net_\,
            in3 => \N__39146\,
            lcout => \comm_spi.n14631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52548\,
            ce => 'H',
            sr => \N__39492\
        );

    \comm_spi.data_tx_i3_12208_12209_reset_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39287\,
            in1 => \N__37359\,
            in2 => \_gnd_net_\,
            in3 => \N__37385\,
            lcout => \comm_spi.n14627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => 'H',
            sr => \N__36795\
        );

    \i2_3_lut_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__45861\,
            in1 => \N__36968\,
            in2 => \_gnd_net_\,
            in3 => \N__49086\,
            lcout => n19902,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_258_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__51645\,
            in1 => \N__49167\,
            in2 => \N__45878\,
            in3 => \N__49874\,
            lcout => OPEN,
            ltout => \n20944_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__49654\,
            in1 => \N__36975\,
            in2 => \N__36984\,
            in3 => \N__36954\,
            lcout => n20964,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_4_lut_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110011"
        )
    port map (
            in0 => \N__49409\,
            in1 => \N__51636\,
            in2 => \N__50031\,
            in3 => \N__49873\,
            lcout => n20962,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_317_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100101111"
        )
    port map (
            in0 => \N__49872\,
            in1 => \N__49408\,
            in2 => \N__51759\,
            in3 => \N__49994\,
            lcout => n4_adj_1586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_298_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__36969\,
            in1 => \N__49653\,
            in2 => \N__50030\,
            in3 => \N__37035\,
            lcout => n20801,
            ltout => \n20801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__49655\,
            in1 => \N__36948\,
            in2 => \N__36942\,
            in3 => \N__36939\,
            lcout => n20829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19129_2_lut_3_lut_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__49993\,
            in1 => \N__51632\,
            in2 => \_gnd_net_\,
            in3 => \N__49871\,
            lcout => n21369,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_1__bdd_4_lut_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__37626\,
            in1 => \N__51637\,
            in2 => \N__49172\,
            in3 => \N__55404\,
            lcout => n22423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__51641\,
            in1 => \N__49412\,
            in2 => \N__50047\,
            in3 => \N__37028\,
            lcout => OPEN,
            ltout => \n2_adj_1581_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22423_bdd_4_lut_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__49413\,
            in1 => \N__36933\,
            in2 => \N__36924\,
            in3 => \N__55405\,
            lcout => n22426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19296_4_lut_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__50035\,
            in1 => \N__55451\,
            in2 => \N__51760\,
            in3 => \N__49088\,
            lcout => OPEN,
            ltout => \n21370_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19388_4_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011011111"
        )
    port map (
            in0 => \N__49411\,
            in1 => \N__56822\,
            in2 => \N__37065\,
            in3 => \N__37062\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i1_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__56823\,
            in1 => \N__37017\,
            in2 => \N__56567\,
            in3 => \N__37056\,
            lcout => comm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54296\,
            ce => \N__37050\,
            sr => \_gnd_net_\
        );

    \i227_2_lut_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50036\,
            in2 => \_gnd_net_\,
            in3 => \N__49848\,
            lcout => n1264,
            ltout => \n1264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_296_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__49566\,
            in1 => \N__49410\,
            in2 => \N__37038\,
            in3 => \N__37215\,
            lcout => n4_adj_1643,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110001011"
        )
    port map (
            in0 => \N__51574\,
            in1 => \N__49402\,
            in2 => \N__37011\,
            in3 => \N__37029\,
            lcout => n8_adj_1582,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_84_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__55136\,
            in1 => \N__45666\,
            in2 => \N__40038\,
            in3 => \N__53671\,
            lcout => \comm_state_3_N_420_3\,
            ltout => \comm_state_3_N_420_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19114_2_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37002\,
            in3 => \N__49403\,
            lcout => OPEN,
            ltout => \n21435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i3_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001110101"
        )
    port map (
            in0 => \N__56830\,
            in1 => \N__56452\,
            in2 => \N__36999\,
            in3 => \N__49143\,
            lcout => comm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54308\,
            ce => \N__36996\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_275_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__51573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49401\,
            lcout => OPEN,
            ltout => \n20937_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_268_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50045\,
            in1 => \N__49847\,
            in2 => \N__37218\,
            in3 => \N__45846\,
            lcout => n20939,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_101_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__56693\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55430\,
            lcout => n20917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_311_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__55429\,
            in1 => \N__56692\,
            in2 => \_gnd_net_\,
            in3 => \N__51572\,
            lcout => n12226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19644_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__37209\,
            in1 => \N__55140\,
            in2 => \N__37203\,
            in3 => \N__53552\,
            lcout => OPEN,
            ltout => \n22261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22261_bdd_4_lut_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__53553\,
            in1 => \N__37172\,
            in2 => \N__37140\,
            in3 => \N__37137\,
            lcout => n22264,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i26_3_lut_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__57477\,
            in1 => \_gnd_net_\,
            in2 => \N__37575\,
            in3 => \N__37923\,
            lcout => OPEN,
            ltout => \n26_adj_1523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19773_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__53554\,
            in1 => \N__55059\,
            in2 => \N__37125\,
            in3 => \N__57156\,
            lcout => OPEN,
            ltout => \n22411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22411_bdd_4_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__53555\,
            in1 => \N__37122\,
            in2 => \N__37095\,
            in3 => \N__37092\,
            lcout => OPEN,
            ltout => \n22414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1553761_i1_3_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37467\,
            in2 => \N__37461\,
            in3 => \N__54745\,
            lcout => OPEN,
            ltout => \n30_adj_1524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i1_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45768\,
            in2 => \N__37458\,
            in3 => \N__51758\,
            lcout => comm_buf_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54321\,
            ce => \N__51383\,
            sr => \N__51302\
        );

    \comm_spi.data_tx_i3_12208_12209_set_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39291\,
            in1 => \N__37355\,
            in2 => \_gnd_net_\,
            in3 => \N__37389\,
            lcout => \comm_spi.n14626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52638\,
            ce => 'H',
            sr => \N__37371\
        );

    \i19037_2_lut_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__57701\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38048\,
            lcout => n21272,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19106_2_lut_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37748\,
            in2 => \_gnd_net_\,
            in3 => \N__57700\,
            lcout => n21568,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i2_12204_12205_set_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38580\,
            in1 => \N__39351\,
            in2 => \_gnd_net_\,
            in3 => \N__38628\,
            lcout => \comm_spi.n14622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52609\,
            ce => 'H',
            sr => \N__39309\
        );

    \comm_spi.i19450_4_lut_3_lut_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55874\,
            in1 => \N__44546\,
            in2 => \_gnd_net_\,
            in3 => \N__39483\,
            lcout => \comm_spi.n22872\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19460_4_lut_3_lut_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37328\,
            in1 => \N__55875\,
            in2 => \_gnd_net_\,
            in3 => \N__45270\,
            lcout => \comm_spi.n22857\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12225_2_lut_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37316\,
            in2 => \_gnd_net_\,
            in3 => \N__38556\,
            lcout => n14647,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i17178_2_lut_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50579\,
            in2 => \_gnd_net_\,
            in3 => \N__49497\,
            lcout => n19783,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_211_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__49498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50580\,
            lcout => n26_adj_1644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19281_2_lut_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49499\,
            in2 => \_gnd_net_\,
            in3 => \N__37656\,
            lcout => n21521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_idxvec_i0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37613\,
            in1 => \N__56929\,
            in2 => \N__43412\,
            in3 => \N__37602\,
            lcout => data_idxvec_0,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => n19634,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37599\,
            in1 => \N__56933\,
            in2 => \N__37574\,
            in3 => \N__37554\,
            lcout => data_idxvec_1,
            ltout => OPEN,
            carryin => n19634,
            carryout => n19635,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i2_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37551\,
            in1 => \N__56930\,
            in2 => \N__47147\,
            in3 => \N__37533\,
            lcout => data_idxvec_2,
            ltout => OPEN,
            carryin => n19635,
            carryout => n19636,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i3_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47097\,
            in1 => \N__56934\,
            in2 => \N__50882\,
            in3 => \N__37530\,
            lcout => data_idxvec_3,
            ltout => OPEN,
            carryin => n19636,
            carryout => n19637,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i4_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37527\,
            in1 => \N__56931\,
            in2 => \N__46217\,
            in3 => \N__37500\,
            lcout => data_idxvec_4,
            ltout => OPEN,
            carryin => n19637,
            carryout => n19638,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i5_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37486\,
            in1 => \N__56935\,
            in2 => \N__51176\,
            in3 => \N__37470\,
            lcout => data_idxvec_5,
            ltout => OPEN,
            carryin => n19638,
            carryout => n19639,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47828\,
            in1 => \N__56932\,
            in2 => \N__46535\,
            in3 => \N__37881\,
            lcout => data_idxvec_6,
            ltout => OPEN,
            carryin => n19639,
            carryout => n19640,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i7_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37877\,
            in1 => \N__56936\,
            in2 => \N__50477\,
            in3 => \N__37854\,
            lcout => data_idxvec_7,
            ltout => OPEN,
            carryin => n19640,
            carryout => n19641,
            clk => \N__54361\,
            ce => \N__37986\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i8_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37847\,
            in1 => \N__57021\,
            in2 => \N__41069\,
            in3 => \N__37830\,
            lcout => data_idxvec_8,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => n19642,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i9_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37823\,
            in1 => \N__56945\,
            in2 => \N__41195\,
            in3 => \N__37797\,
            lcout => data_idxvec_9,
            ltout => OPEN,
            carryin => n19642,
            carryout => n19643,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i10_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37794\,
            in1 => \N__57022\,
            in2 => \N__41244\,
            in3 => \N__37776\,
            lcout => data_idxvec_10,
            ltout => OPEN,
            carryin => n19643,
            carryout => n19644,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i11_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__44426\,
            in1 => \N__56946\,
            in2 => \N__40953\,
            in3 => \N__37773\,
            lcout => data_idxvec_11,
            ltout => OPEN,
            carryin => n19644,
            carryout => n19645,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i12_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37770\,
            in1 => \N__57023\,
            in2 => \N__37749\,
            in3 => \N__37731\,
            lcout => data_idxvec_12,
            ltout => OPEN,
            carryin => n19645,
            carryout => n19646,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i13_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37727\,
            in1 => \N__56947\,
            in2 => \N__37694\,
            in3 => \N__37674\,
            lcout => data_idxvec_13,
            ltout => OPEN,
            carryin => n19646,
            carryout => n19647,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i14_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__38069\,
            in1 => \N__57024\,
            in2 => \N__38049\,
            in3 => \N__38031\,
            lcout => data_idxvec_14,
            ltout => OPEN,
            carryin => n19647,
            carryout => n19648,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i15_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38018\,
            in1 => \N__38000\,
            in2 => \N__57095\,
            in3 => \N__38007\,
            lcout => data_idxvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54374\,
            ce => \N__37982\,
            sr => \_gnd_net_\
        );

    \data_cntvec_i0_i0_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43387\,
            in2 => \N__37962\,
            in3 => \_gnd_net_\,
            lcout => data_cntvec_0,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => n19595,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37919\,
            in2 => \_gnd_net_\,
            in3 => \N__37899\,
            lcout => data_cntvec_1,
            ltout => OPEN,
            carryin => n19595,
            carryout => n19596,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i2_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47123\,
            in2 => \_gnd_net_\,
            in3 => \N__37896\,
            lcout => data_cntvec_2,
            ltout => OPEN,
            carryin => n19596,
            carryout => n19597,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i3_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50854\,
            in2 => \_gnd_net_\,
            in3 => \N__37893\,
            lcout => data_cntvec_3,
            ltout => OPEN,
            carryin => n19597,
            carryout => n19598,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i4_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46193\,
            in2 => \_gnd_net_\,
            in3 => \N__37890\,
            lcout => data_cntvec_4,
            ltout => OPEN,
            carryin => n19598,
            carryout => n19599,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i5_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51151\,
            in2 => \_gnd_net_\,
            in3 => \N__37887\,
            lcout => data_cntvec_5,
            ltout => OPEN,
            carryin => n19599,
            carryout => n19600,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i6_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46507\,
            in2 => \_gnd_net_\,
            in3 => \N__37884\,
            lcout => data_cntvec_6,
            ltout => OPEN,
            carryin => n19600,
            carryout => n19601,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i7_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50453\,
            in2 => \_gnd_net_\,
            in3 => \N__38163\,
            lcout => data_cntvec_7,
            ltout => OPEN,
            carryin => n19601,
            carryout => n19602,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38559\,
            sr => \N__38481\
        );

    \data_cntvec_i0_i8_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41045\,
            in2 => \_gnd_net_\,
            in3 => \N__38160\,
            lcout => data_cntvec_8,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => n19603,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \data_cntvec_i0_i9_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41171\,
            in2 => \_gnd_net_\,
            in3 => \N__38157\,
            lcout => data_cntvec_9,
            ltout => OPEN,
            carryin => n19603,
            carryout => n19604,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \data_cntvec_i0_i10_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41225\,
            in2 => \_gnd_net_\,
            in3 => \N__38154\,
            lcout => data_cntvec_10,
            ltout => OPEN,
            carryin => n19604,
            carryout => n19605,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \data_cntvec_i0_i11_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40937\,
            in2 => \_gnd_net_\,
            in3 => \N__38151\,
            lcout => data_cntvec_11,
            ltout => OPEN,
            carryin => n19605,
            carryout => n19606,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \data_cntvec_i0_i12_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38144\,
            in2 => \_gnd_net_\,
            in3 => \N__38130\,
            lcout => data_cntvec_12,
            ltout => OPEN,
            carryin => n19606,
            carryout => n19607,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \data_cntvec_i0_i13_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38123\,
            in2 => \_gnd_net_\,
            in3 => \N__38109\,
            lcout => data_cntvec_13,
            ltout => OPEN,
            carryin => n19607,
            carryout => n19608,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \data_cntvec_i0_i14_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38106\,
            in2 => \_gnd_net_\,
            in3 => \N__38094\,
            lcout => data_cntvec_14,
            ltout => OPEN,
            carryin => n19608,
            carryout => n19609,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \data_cntvec_i0_i15_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38084\,
            in2 => \_gnd_net_\,
            in3 => \N__38091\,
            lcout => data_cntvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38557\,
            sr => \N__38489\
        );

    \i6389_3_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41978\,
            in1 => \N__50302\,
            in2 => \_gnd_net_\,
            in3 => \N__47681\,
            lcout => n8_adj_1563,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_171_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__38450\,
            in1 => \N__41350\,
            in2 => \N__38433\,
            in3 => \N__43357\,
            lcout => n17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6399_3_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47895\,
            in1 => \N__38394\,
            in2 => \_gnd_net_\,
            in3 => \N__47682\,
            lcout => n8_adj_1565,
            ltout => \n8_adj_1565_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i6_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56169\,
            in1 => \N__56924\,
            in2 => \N__38397\,
            in3 => \N__38268\,
            lcout => data_index_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15090_3_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51435\,
            in1 => \N__40568\,
            in2 => \_gnd_net_\,
            in3 => \N__47680\,
            lcout => n17489,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_188_i9_2_lut_3_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__55176\,
            in1 => \N__57781\,
            in2 => \_gnd_net_\,
            in3 => \N__53723\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__56923\,
            in1 => \N__56168\,
            in2 => \N__41123\,
            in3 => \N__41135\,
            lcout => \data_index_9_N_216_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__56925\,
            in1 => \N__56420\,
            in2 => \N__38280\,
            in3 => \N__38267\,
            lcout => \data_index_9_N_216_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6369_3_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39078\,
            in1 => \N__40122\,
            in2 => \_gnd_net_\,
            in3 => \N__47703\,
            lcout => n8_adj_1559,
            ltout => \n8_adj_1559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56419\,
            in1 => \N__39053\,
            in2 => \N__39042\,
            in3 => \N__56928\,
            lcout => \data_index_9_N_216_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__56927\,
            in1 => \N__38951\,
            in2 => \N__56517\,
            in3 => \N__42035\,
            lcout => \data_index_9_N_216_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__42023\,
            in1 => \N__56926\,
            in2 => \N__56516\,
            in3 => \N__42002\,
            lcout => \data_index_9_N_216_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_16MHz_I_0_3_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38766\,
            in1 => \N__38703\,
            in2 => \_gnd_net_\,
            in3 => \N__38679\,
            lcout => \DDS_MCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i1_12200_12201_reset_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38607\,
            in1 => \N__41790\,
            in2 => \_gnd_net_\,
            in3 => \N__38591\,
            lcout => \comm_spi.n14619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52626\,
            ce => 'H',
            sr => \N__39363\
        );

    \comm_spi.RESET_I_0_98_2_lut_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__39605\,
            in1 => \_gnd_net_\,
            in2 => \N__55872\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19465_4_lut_3_lut_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38606\,
            in1 => \N__42494\,
            in2 => \_gnd_net_\,
            in3 => \N__55858\,
            lcout => \comm_spi.n22884\,
            ltout => \comm_spi.n22884_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i1_12200_12201_set_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41789\,
            in1 => \_gnd_net_\,
            in2 => \N__38595\,
            in3 => \N__38592\,
            lcout => \comm_spi.n14618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52640\,
            ce => 'H',
            sr => \N__39375\
        );

    \comm_spi.RESET_I_0_106_2_lut_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39604\,
            in2 => \_gnd_net_\,
            in3 => \N__55849\,
            lcout => \comm_spi.data_tx_7__N_792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19430_4_lut_3_lut_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39606\,
            in1 => \_gnd_net_\,
            in2 => \N__55873\,
            in3 => \N__39337\,
            lcout => \comm_spi.n22881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_105_2_lut_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39658\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55848\,
            lcout => \comm_spi.data_tx_7__N_789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_97_2_lut_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55850\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39659\,
            lcout => \comm_spi.data_tx_7__N_771\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19440_4_lut_3_lut_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39660\,
            in1 => \N__39275\,
            in2 => \_gnd_net_\,
            in3 => \N__55857\,
            lcout => \comm_spi.n22878\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \wdtick_cnt_3763_3764__i1_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__39259\,
            in1 => \N__39241\,
            in2 => \_gnd_net_\,
            in3 => \N__39222\,
            lcout => wdtick_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39206\,
            ce => \N__39447\,
            sr => \N__39413\
        );

    \wdtick_cnt_3763_3764__i3_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010100000"
        )
    port map (
            in0 => \N__39224\,
            in1 => \_gnd_net_\,
            in2 => \N__39246\,
            in3 => \N__39260\,
            lcout => wdtick_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39206\,
            ce => \N__39447\,
            sr => \N__39413\
        );

    \wdtick_cnt_3763_3764__i2_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39240\,
            in2 => \_gnd_net_\,
            in3 => \N__39223\,
            lcout => wdtick_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39206\,
            ce => \N__39447\,
            sr => \N__39413\
        );

    \comm_spi.data_tx_i4_12212_12213_set_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39147\,
            in1 => \N__39135\,
            in2 => \_gnd_net_\,
            in3 => \N__39102\,
            lcout => \comm_spi.n14630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52610\,
            ce => 'H',
            sr => \N__39462\
        );

    \i46_2_lut_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__50013\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51720\,
            lcout => n23_adj_1620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9325_1_lut_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44632\,
            lcout => n11741,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_244_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__56956\,
            in1 => \N__39438\,
            in2 => \N__55512\,
            in3 => \N__49590\,
            lcout => n11390,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18382_2_lut_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__49487\,
            in1 => \_gnd_net_\,
            in2 => \N__51859\,
            in3 => \_gnd_net_\,
            lcout => n20992,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6834_2_lut_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51714\,
            in2 => \_gnd_net_\,
            in3 => \N__49486\,
            lcout => n9255,
            ltout => \n9255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_259_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__49589\,
            in1 => \N__55447\,
            in2 => \N__39432\,
            in3 => \N__56957\,
            lcout => n14737,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \flagcntwd_303_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51719\,
            in2 => \_gnd_net_\,
            in3 => \N__49488\,
            lcout => flagcntwd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54291\,
            ce => \N__39390\,
            sr => \N__39569\
        );

    \i1_4_lut_adj_279_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__49588\,
            in1 => \N__56953\,
            in2 => \N__55510\,
            in3 => \N__49619\,
            lcout => n12336,
            ltout => \n12336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12386_3_lut_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__56954\,
            in1 => \_gnd_net_\,
            in2 => \N__39378\,
            in3 => \N__52265\,
            lcout => n14799,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_63_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__51718\,
            in1 => \_gnd_net_\,
            in2 => \N__55511\,
            in3 => \N__56955\,
            lcout => n20378,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_4_i1_3_lut_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50732\,
            in1 => \N__41484\,
            in2 => \_gnd_net_\,
            in3 => \N__47783\,
            lcout => n1_adj_1591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_4_i2_3_lut_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45531\,
            in1 => \N__39546\,
            in2 => \_gnd_net_\,
            in3 => \N__50731\,
            lcout => n2_adj_1592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19294_2_lut_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39537\,
            lcout => OPEN,
            ltout => \n21538_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__39498\,
            in1 => \N__50571\,
            in2 => \N__39516\,
            in3 => \N__52386\,
            lcout => OPEN,
            ltout => \n22369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i4_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50572\,
            in1 => \N__39513\,
            in2 => \N__39507\,
            in3 => \N__39504\,
            lcout => comm_tx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54297\,
            ce => \N__45243\,
            sr => \N__45164\
        );

    \mux_137_Mux_4_i4_3_lut_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39885\,
            in1 => \N__42603\,
            in2 => \_gnd_net_\,
            in3 => \N__50729\,
            lcout => n4_adj_1593,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_103_2_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55843\,
            in2 => \_gnd_net_\,
            in3 => \N__39475\,
            lcout => \comm_spi.data_tx_7__N_783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_95_2_lut_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__39476\,
            in1 => \_gnd_net_\,
            in2 => \N__55871\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__39708\,
            in1 => \N__50754\,
            in2 => \N__45408\,
            in3 => \N__52404\,
            lcout => OPEN,
            ltout => \n22393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22393_bdd_4_lut_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52405\,
            in1 => \N__44759\,
            in2 => \N__39696\,
            in3 => \N__48080\,
            lcout => n22396,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_2_i4_3_lut_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39834\,
            in1 => \N__42546\,
            in2 => \_gnd_net_\,
            in3 => \N__50756\,
            lcout => OPEN,
            ltout => \n4_adj_1595_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18586_4_lut_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__52406\,
            in1 => \N__39693\,
            in2 => \N__39672\,
            in3 => \N__50779\,
            lcout => OPEN,
            ltout => \n21196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i2_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__50598\,
            in1 => \N__39669\,
            in2 => \N__39663\,
            in3 => \_gnd_net_\,
            lcout => comm_tx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54309\,
            ce => \N__45226\,
            sr => \N__45157\
        );

    \mux_137_Mux_1_i4_3_lut_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50755\,
            in1 => \N__39813\,
            in2 => \_gnd_net_\,
            in3 => \N__43194\,
            lcout => OPEN,
            ltout => \n4_adj_1596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18442_4_lut_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__39642\,
            in1 => \N__50757\,
            in2 => \N__39624\,
            in3 => \N__52407\,
            lcout => OPEN,
            ltout => \n21052_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i1_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39621\,
            in2 => \N__39609\,
            in3 => \N__50597\,
            lcout => comm_tx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54309\,
            ce => \N__45226\,
            sr => \N__45157\
        );

    \comm_buf_5__i0_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39588\,
            in1 => \N__51653\,
            in2 => \_gnd_net_\,
            in3 => \N__53037\,
            lcout => comm_buf_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_buf_5__i7_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51652\,
            in1 => \_gnd_net_\,
            in2 => \N__39960\,
            in3 => \N__50389\,
            lcout => comm_buf_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_buf_5__i6_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46446\,
            in1 => \N__39930\,
            in2 => \_gnd_net_\,
            in3 => \N__51656\,
            lcout => comm_buf_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_buf_5__i5_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51651\,
            in1 => \N__52111\,
            in2 => \_gnd_net_\,
            in3 => \N__39915\,
            lcout => comm_buf_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_buf_5__i4_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46776\,
            in1 => \N__39900\,
            in2 => \_gnd_net_\,
            in3 => \N__51655\,
            lcout => comm_buf_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_buf_5__i3_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51650\,
            in1 => \N__51107\,
            in2 => \_gnd_net_\,
            in3 => \N__39876\,
            lcout => comm_buf_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_buf_5__i2_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47231\,
            in1 => \N__39849\,
            in2 => \_gnd_net_\,
            in3 => \N__51654\,
            lcout => comm_buf_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_buf_5__i1_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51649\,
            in1 => \N__45792\,
            in2 => \_gnd_net_\,
            in3 => \N__39828\,
            lcout => comm_buf_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54322\,
            ce => \N__42858\,
            sr => \N__42849\
        );

    \comm_cmd_0__bdd_4_lut_19664_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__39800\,
            in1 => \N__57475\,
            in2 => \N__55211\,
            in3 => \N__39761\,
            lcout => OPEN,
            ltout => \n22237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22237_bdd_4_lut_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__55132\,
            in1 => \N__39738\,
            in2 => \N__40245\,
            in3 => \N__40242\,
            lcout => n22240,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18452_4_lut_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__57476\,
            in1 => \N__40215\,
            in2 => \N__55210\,
            in3 => \N__41151\,
            lcout => OPEN,
            ltout => \n21062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__53750\,
            in1 => \N__40206\,
            in2 => \N__40191\,
            in3 => \N__54694\,
            lcout => OPEN,
            ltout => \n22447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22447_bdd_4_lut_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__40188\,
            in1 => \N__40182\,
            in2 => \N__40167\,
            in3 => \N__54693\,
            lcout => OPEN,
            ltout => \n22450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i1_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__52026\,
            in1 => \N__45793\,
            in2 => \N__40164\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54334\,
            ce => \N__46164\,
            sr => \N__43698\
        );

    \i36_4_lut_4_lut_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100011011100"
        )
    port map (
            in0 => \N__57474\,
            in1 => \N__54692\,
            in2 => \N__55209\,
            in3 => \N__53749\,
            lcout => n30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19649_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__41829\,
            in1 => \N__54979\,
            in2 => \N__40029\,
            in3 => \N__53667\,
            lcout => OPEN,
            ltout => \n22273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22273_bdd_4_lut_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__53668\,
            in1 => \N__40020\,
            in2 => \N__40008\,
            in3 => \N__40005\,
            lcout => n22276,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22285_bdd_4_lut_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__39993\,
            in1 => \N__40392\,
            in2 => \N__39978\,
            in3 => \N__53669\,
            lcout => OPEN,
            ltout => \n22288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1552555_i1_3_lut_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54695\,
            in1 => \_gnd_net_\,
            in2 => \N__40473\,
            in3 => \N__40470\,
            lcout => OPEN,
            ltout => \n30_adj_1539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i6_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46447\,
            in2 => \N__40464\,
            in3 => \N__51872\,
            lcout => comm_buf_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54348\,
            ce => \N__46167\,
            sr => \N__43700\
        );

    \mux_128_Mux_6_i19_3_lut_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40461\,
            in1 => \N__40433\,
            in2 => \_gnd_net_\,
            in3 => \N__57736\,
            lcout => OPEN,
            ltout => \n19_adj_1536_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19659_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__40404\,
            in1 => \N__54978\,
            in2 => \N__40395\,
            in3 => \N__53666\,
            lcout => n22285,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19679_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__57624\,
            in1 => \N__41387\,
            in2 => \N__40385\,
            in3 => \N__55215\,
            lcout => OPEN,
            ltout => \n22303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22303_bdd_4_lut_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__55216\,
            in1 => \N__40347\,
            in2 => \N__40320\,
            in3 => \N__40316\,
            lcout => n22306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22243_bdd_4_lut_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__40287\,
            in1 => \N__40251\,
            in2 => \N__40275\,
            in3 => \N__53728\,
            lcout => n22246,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19634_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__41805\,
            in1 => \N__55214\,
            in2 => \N__40260\,
            in3 => \N__53727\,
            lcout => n22243,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18482_3_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53729\,
            in1 => \N__40545\,
            in2 => \_gnd_net_\,
            in3 => \N__40539\,
            lcout => OPEN,
            ltout => \n21092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1551349_i1_3_lut_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40530\,
            in2 => \N__40524\,
            in3 => \N__54631\,
            lcout => OPEN,
            ltout => \n30_adj_1542_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i4_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__51904\,
            in1 => \N__46787\,
            in2 => \N__40521\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54362\,
            ce => \N__46168\,
            sr => \N__43723\
        );

    \comm_cmd_1__bdd_4_lut_19719_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__55217\,
            in1 => \N__53763\,
            in2 => \N__53865\,
            in3 => \N__41205\,
            lcout => OPEN,
            ltout => \n22357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22357_bdd_4_lut_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__53764\,
            in1 => \N__40518\,
            in2 => \N__40509\,
            in3 => \N__40791\,
            lcout => OPEN,
            ltout => \n22360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18527_3_lut_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54691\,
            in1 => \_gnd_net_\,
            in2 => \N__40506\,
            in3 => \N__40479\,
            lcout => OPEN,
            ltout => \n21137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i2_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52032\,
            in2 => \N__40503\,
            in3 => \N__47244\,
            lcout => comm_buf_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54375\,
            ce => \N__46169\,
            sr => \N__43724\
        );

    \n22327_bdd_4_lut_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__53762\,
            in1 => \N__40680\,
            in2 => \N__40500\,
            in3 => \N__40488\,
            lcout => n22330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_6_i16_3_lut_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40750\,
            in1 => \N__40729\,
            in2 => \_gnd_net_\,
            in3 => \N__57614\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_3_i26_3_lut_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57615\,
            in1 => \N__40949\,
            in2 => \_gnd_net_\,
            in3 => \N__40938\,
            lcout => OPEN,
            ltout => \n26_adj_1544_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18475_4_lut_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__55036\,
            in1 => \N__40917\,
            in2 => \N__40902\,
            in3 => \N__57616\,
            lcout => n21085,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18478_3_lut_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57618\,
            in1 => \N__40899\,
            in2 => \_gnd_net_\,
            in3 => \N__40821\,
            lcout => n21088,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18567_3_lut_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55035\,
            in1 => \N__41357\,
            in2 => \_gnd_net_\,
            in3 => \N__40785\,
            lcout => n21177,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i6_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__40754\,
            in1 => \N__40668\,
            in2 => \N__47897\,
            in3 => \N__44971\,
            lcout => buf_dds1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i6_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56450\,
            in1 => \N__40730\,
            in2 => \N__47896\,
            in3 => \N__48027\,
            lcout => buf_dds0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18463_3_lut_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57617\,
            in1 => \N__40715\,
            in2 => \_gnd_net_\,
            in3 => \N__44678\,
            lcout => n21073,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i11_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__43966\,
            in1 => \N__40666\,
            in2 => \N__44979\,
            in3 => \N__44177\,
            lcout => buf_dds1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i5_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__57124\,
            in1 => \N__56223\,
            in2 => \N__56598\,
            in3 => \N__56030\,
            lcout => data_index_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18540_3_lut_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41240\,
            in1 => \N__57803\,
            in2 => \_gnd_net_\,
            in3 => \N__41221\,
            lcout => n21150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18450_3_lut_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__57802\,
            in1 => \_gnd_net_\,
            in2 => \N__41196\,
            in3 => \N__41167\,
            lcout => n21060,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i3_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__41142\,
            in1 => \N__57125\,
            in2 => \N__56343\,
            in3 => \N__41124\,
            lcout => data_index_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18555_3_lut_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41070\,
            in1 => \N__57801\,
            in2 => \_gnd_net_\,
            in3 => \N__41041\,
            lcout => n21165,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18474_4_lut_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__57800\,
            in1 => \N__55125\,
            in2 => \N__41904\,
            in3 => \N__41025\,
            lcout => n21084,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i2_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__46579\,
            in1 => \N__48066\,
            in2 => \N__56321\,
            in3 => \N__44316\,
            lcout => \acadc_skipCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6439_3_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47691\,
            in1 => \N__48059\,
            in2 => \_gnd_net_\,
            in3 => \N__40996\,
            lcout => n8_adj_1571,
            ltout => \n8_adj_1571_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i2_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56202\,
            in1 => \N__57094\,
            in2 => \N__41007\,
            in3 => \N__45093\,
            lcout => data_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i10_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__40969\,
            in1 => \N__56203\,
            in2 => \N__44769\,
            in3 => \N__48024\,
            lcout => buf_dds0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_304_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__41552\,
            in1 => \N__57093\,
            in2 => \N__56320\,
            in3 => \N__41777\,
            lcout => n12429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6973_2_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51959\,
            in2 => \_gnd_net_\,
            in3 => \N__55499\,
            lcout => n9306,
            ltout => \n9306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i13_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__48025\,
            in1 => \N__43593\,
            in2 => \N__41634\,
            in3 => \N__41617\,
            lcout => buf_dds0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_165_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__41601\,
            in1 => \N__41583\,
            in2 => \N__46580\,
            in3 => \N__46972\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_248_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000100"
        )
    port map (
            in0 => \N__41553\,
            in1 => \N__57122\,
            in2 => \N__41541\,
            in3 => \N__56170\,
            lcout => n12381,
            ltout => \n12381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i5_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__56175\,
            in1 => \N__41465\,
            in2 => \N__41403\,
            in3 => \N__41377\,
            lcout => \VAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i0_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__43282\,
            in1 => \N__44329\,
            in2 => \N__56291\,
            in3 => \N__43361\,
            lcout => \acadc_skipCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i6_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56174\,
            in1 => \N__44330\,
            in2 => \N__47901\,
            in3 => \N__41358\,
            lcout => \acadc_skipCount_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19329_4_lut_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000110"
        )
    port map (
            in0 => \N__41323\,
            in1 => \N__42267\,
            in2 => \N__42132\,
            in3 => \N__43020\,
            lcout => \SIG_DDS.n12722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6379_3_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43783\,
            in1 => \N__42063\,
            in2 => \_gnd_net_\,
            in3 => \N__47702\,
            lcout => n8_adj_1561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i7_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__57123\,
            in1 => \N__42024\,
            in2 => \N__42012\,
            in3 => \N__56316\,
            lcout => data_index_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_3_i23_3_lut_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41954\,
            in1 => \N__57758\,
            in2 => \_gnd_net_\,
            in3 => \N__41934\,
            lcout => n23_adj_1543,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i0_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56315\,
            in1 => \N__41892\,
            in2 => \N__43808\,
            in3 => \N__44611\,
            lcout => buf_control_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19085_2_lut_LC_17_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41838\,
            in2 => \_gnd_net_\,
            in3 => \N__57822\,
            lcout => n21273,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19092_2_lut_LC_17_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41817\,
            in2 => \_gnd_net_\,
            in3 => \N__57821\,
            lcout => n21569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12174_12175_set_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__58293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52602\,
            ce => 'H',
            sr => \N__42465\
        );

    \comm_spi.data_tx_i5_12216_12217_reset_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44528\,
            in1 => \N__44561\,
            in2 => \_gnd_net_\,
            in3 => \N__44516\,
            lcout => \comm_spi.n14635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52586\,
            ce => 'H',
            sr => \N__42360\
        );

    \comm_spi.data_tx_i6_12220_12221_reset_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44469\,
            in1 => \N__44486\,
            in2 => \_gnd_net_\,
            in3 => \N__44456\,
            lcout => \comm_spi.n14639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__42372\
        );

    \comm_spi.RESET_I_0_101_2_lut_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45260\,
            in2 => \_gnd_net_\,
            in3 => \N__55757\,
            lcout => \comm_spi.data_tx_7__N_777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_102_2_lut_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42734\,
            in2 => \_gnd_net_\,
            in3 => \N__55758\,
            lcout => \comm_spi.data_tx_7__N_780\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_6_i4_3_lut_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42348\,
            in1 => \N__42645\,
            in2 => \_gnd_net_\,
            in3 => \N__50790\,
            lcout => n4_adj_1590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19455_4_lut_3_lut_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44485\,
            in1 => \N__42735\,
            in2 => \_gnd_net_\,
            in3 => \N__55759\,
            lcout => \comm_spi.n22869\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19580_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__42324\,
            in1 => \N__50599\,
            in2 => \N__42297\,
            in3 => \N__52387\,
            lcout => OPEN,
            ltout => \n22183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i0_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50600\,
            in1 => \N__42522\,
            in2 => \N__42339\,
            in3 => \N__42501\,
            lcout => comm_tx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54310\,
            ce => \N__45236\,
            sr => \N__45171\
        );

    \mux_137_Mux_0_i4_3_lut_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42336\,
            in1 => \N__42699\,
            in2 => \_gnd_net_\,
            in3 => \N__50795\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18964_2_lut_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42318\,
            lcout => n21211,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_0_i1_3_lut_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43291\,
            in1 => \N__43825\,
            in2 => \_gnd_net_\,
            in3 => \N__50797\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_0_i2_3_lut_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50796\,
            in1 => \N__45552\,
            in2 => \_gnd_net_\,
            in3 => \N__42513\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_99_2_lut_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55847\,
            lcout => \comm_spi.data_tx_7__N_773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15080_3_lut_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42621\,
            in1 => \N__43567\,
            in2 => \_gnd_net_\,
            in3 => \N__50596\,
            lcout => OPEN,
            ltout => \n17479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i5_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__42393\,
            in1 => \N__42417\,
            in2 => \N__42450\,
            in3 => \N__50778\,
            lcout => comm_tx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54323\,
            ce => \N__45235\,
            sr => \N__45173\
        );

    \i19282_2_lut_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45450\,
            in2 => \_gnd_net_\,
            in3 => \N__50593\,
            lcout => n21212,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15081_3_lut_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50595\,
            in1 => \N__42447\,
            in2 => \_gnd_net_\,
            in3 => \N__42429\,
            lcout => n17480,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15083_3_lut_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42408\,
            in1 => \N__51436\,
            in2 => \_gnd_net_\,
            in3 => \N__50594\,
            lcout => OPEN,
            ltout => \n17482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19699_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__42402\,
            in1 => \N__50777\,
            in2 => \N__42396\,
            in3 => \N__52408\,
            lcout => n22189,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_94_2_lut_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__42728\,
            in1 => \N__55827\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_768\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__42717\,
            in1 => \N__52016\,
            in2 => \_gnd_net_\,
            in3 => \N__53036\,
            lcout => comm_buf_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \comm_buf_4__i7_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52015\,
            in1 => \N__50410\,
            in2 => \_gnd_net_\,
            in3 => \N__42690\,
            lcout => comm_buf_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \comm_buf_4__i6_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__42660\,
            in1 => \N__52017\,
            in2 => \_gnd_net_\,
            in3 => \N__46462\,
            lcout => comm_buf_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \comm_buf_4__i5_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52014\,
            in1 => \N__52113\,
            in2 => \_gnd_net_\,
            in3 => \N__42636\,
            lcout => comm_buf_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \comm_buf_4__i4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46786\,
            in1 => \N__42615\,
            in2 => \_gnd_net_\,
            in3 => \N__52019\,
            lcout => comm_buf_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \comm_buf_4__i3_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52013\,
            in1 => \N__51110\,
            in2 => \_gnd_net_\,
            in3 => \N__42591\,
            lcout => comm_buf_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \comm_buf_4__i2_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47232\,
            in1 => \N__42564\,
            in2 => \_gnd_net_\,
            in3 => \N__52018\,
            lcout => comm_buf_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \comm_buf_4__i1_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52012\,
            in1 => \N__45787\,
            in2 => \_gnd_net_\,
            in3 => \N__42540\,
            lcout => comm_buf_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54335\,
            ce => \N__45810\,
            sr => \N__42843\
        );

    \SIG_DDS.bit_cnt_i3_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__43170\,
            in1 => \N__43091\,
            in2 => \N__43127\,
            in3 => \N__43184\,
            lcout => \SIG_DDS.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54349\,
            ce => \N__43074\,
            sr => \N__42885\
        );

    \SIG_DDS.bit_cnt_i1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43116\,
            in2 => \_gnd_net_\,
            in3 => \N__43168\,
            lcout => \SIG_DDS.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54349\,
            ce => \N__43074\,
            sr => \N__42885\
        );

    \SIG_DDS.bit_cnt_i2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__43169\,
            in1 => \_gnd_net_\,
            in2 => \N__43126\,
            in3 => \N__43090\,
            lcout => \SIG_DDS.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54349\,
            ce => \N__43074\,
            sr => \N__42885\
        );

    \i1_3_lut_adj_277_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__45882\,
            in1 => \N__45916\,
            in2 => \_gnd_net_\,
            in3 => \N__46092\,
            lcout => n12220,
            ltout => \n12220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12372_2_lut_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__57069\,
            in1 => \_gnd_net_\,
            in2 => \N__42852\,
            in3 => \_gnd_net_\,
            lcout => n14785,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12337_2_lut_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57067\,
            in2 => \_gnd_net_\,
            in3 => \N__46123\,
            lcout => n14750,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12365_2_lut_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__57068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45806\,
            lcout => n14778,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i7_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52020\,
            in1 => \N__50411\,
            in2 => \_gnd_net_\,
            in3 => \N__42831\,
            lcout => comm_buf_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54363\,
            ce => \N__46165\,
            sr => \N__43699\
        );

    \comm_buf_0__i5_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52117\,
            in1 => \N__43623\,
            in2 => \_gnd_net_\,
            in3 => \N__52021\,
            lcout => comm_buf_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54363\,
            ce => \N__46165\,
            sr => \N__43699\
        );

    \n22213_bdd_4_lut_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__53755\,
            in1 => \N__43422\,
            in2 => \N__43521\,
            in3 => \N__43482\,
            lcout => n22216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19611_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__43467\,
            in1 => \N__55151\,
            in2 => \N__43449\,
            in3 => \N__53754\,
            lcout => n22213,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_0_i26_3_lut_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43416\,
            in1 => \N__57626\,
            in2 => \_gnd_net_\,
            in3 => \N__43392\,
            lcout => OPEN,
            ltout => \n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19593_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__52695\,
            in1 => \N__55152\,
            in2 => \N__43368\,
            in3 => \N__53756\,
            lcout => OPEN,
            ltout => \n22201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22201_bdd_4_lut_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__53757\,
            in1 => \N__43365\,
            in2 => \N__43341\,
            in3 => \N__43338\,
            lcout => OPEN,
            ltout => \n22204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1556173_i1_3_lut_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43311\,
            in2 => \N__43305\,
            in3 => \N__54746\,
            lcout => OPEN,
            ltout => \n30_adj_1485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i0_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__52022\,
            in1 => \_gnd_net_\,
            in2 => \N__43302\,
            in3 => \N__53051\,
            lcout => comm_buf_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54376\,
            ce => \N__51381\,
            sr => \N__51277\
        );

    \comm_cmd_0__bdd_4_lut_19669_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__44108\,
            in1 => \N__55160\,
            in2 => \N__43229\,
            in3 => \N__57625\,
            lcout => OPEN,
            ltout => \n22297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22297_bdd_4_lut_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__55161\,
            in1 => \N__44001\,
            in2 => \N__43974\,
            in3 => \N__43970\,
            lcout => n22300,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22309_bdd_4_lut_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__43941\,
            in1 => \N__54697\,
            in2 => \N__43932\,
            in3 => \N__44340\,
            lcout => OPEN,
            ltout => \n22312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i3_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__51114\,
            in1 => \_gnd_net_\,
            in2 => \N__43923\,
            in3 => \N__51993\,
            lcout => comm_buf_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54390\,
            ce => \N__46166\,
            sr => \N__43710\
        );

    \comm_cmd_0__bdd_4_lut_19616_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__55034\,
            in1 => \N__57604\,
            in2 => \N__43920\,
            in3 => \N__43881\,
            lcout => n22219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18461_3_lut_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__43854\,
            in1 => \_gnd_net_\,
            in2 => \N__44361\,
            in3 => \N__54687\,
            lcout => OPEN,
            ltout => \n21071_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i0_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51992\,
            in2 => \N__43839\,
            in3 => \N__53055\,
            lcout => comm_buf_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54402\,
            ce => \N__46173\,
            sr => \N__43725\
        );

    \i19115_4_lut_4_lut_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101101011"
        )
    port map (
            in0 => \N__57603\,
            in1 => \N__54686\,
            in2 => \N__55147\,
            in3 => \N__53672\,
            lcout => n21341,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22219_bdd_4_lut_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__43656\,
            in1 => \N__55188\,
            in2 => \N__44616\,
            in3 => \N__43650\,
            lcout => n22222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15338_2_lut_3_lut_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__44187\,
            in1 => \_gnd_net_\,
            in2 => \N__55556\,
            in3 => \N__51960\,
            lcout => n14_adj_1578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_187_i9_2_lut_3_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__53765\,
            in1 => \N__57759\,
            in2 => \_gnd_net_\,
            in3 => \N__55187\,
            lcout => n9_adj_1415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18557_4_lut_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__55189\,
            in1 => \N__57804\,
            in2 => \N__44394\,
            in3 => \N__44376\,
            lcout => OPEN,
            ltout => \n21167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18460_3_lut_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53761\,
            in2 => \N__44370\,
            in3 => \N__44367\,
            lcout => n21070,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19684_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__54696\,
            in1 => \N__44352\,
            in2 => \N__53796\,
            in3 => \N__44346\,
            lcout => n22309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i3_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56179\,
            in1 => \N__46915\,
            in2 => \N__51021\,
            in3 => \N__48026\,
            lcout => buf_dds0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i7_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56220\,
            in1 => \N__44317\,
            in2 => \N__50322\,
            in3 => \N__46976\,
            lcout => \acadc_skipCount_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i4_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56180\,
            in1 => \N__44820\,
            in2 => \N__44197\,
            in3 => \N__44104\,
            lcout => \IAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds1_305_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000110100000"
        )
    port map (
            in0 => \N__56221\,
            in1 => \N__44085\,
            in2 => \N__44032\,
            in3 => \N__57092\,
            lcout => trig_dds1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__57091\,
            in1 => \N__45099\,
            in2 => \N__56292\,
            in3 => \N__45092\,
            lcout => \data_index_9_N_216_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i3_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111110101010"
        )
    port map (
            in0 => \N__46945\,
            in1 => \N__47092\,
            in2 => \N__57143\,
            in3 => \N__44970\,
            lcout => buf_dds1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i3_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56222\,
            in1 => \N__44819\,
            in2 => \N__44786\,
            in3 => \N__44668\,
            lcout => \IAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15107_2_lut_2_lut_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__44649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44612\,
            lcout => \CONT_SD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_18_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_12182_12183_reset_LC_18_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55601\,
            lcout => \comm_spi.n14601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54283\,
            ce => 'H',
            sr => \N__44577\
        );

    \comm_spi.data_tx_i5_12216_12217_set_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44562\,
            in1 => \N__44535\,
            in2 => \_gnd_net_\,
            in3 => \N__44517\,
            lcout => \comm_spi.n14634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52587\,
            ce => 'H',
            sr => \N__44499\
        );

    \comm_spi.data_tx_i6_12220_12221_set_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44487\,
            in1 => \N__44468\,
            in2 => \_gnd_net_\,
            in3 => \N__44457\,
            lcout => \comm_spi.n14638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52531\,
            ce => 'H',
            sr => \N__45375\
        );

    \ADC_VDC.genclk.i19300_4_lut_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__48098\,
            in1 => \N__48191\,
            in2 => \N__48144\,
            in3 => \N__48206\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n21446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19039_4_lut_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45381\,
            in1 => \N__45393\,
            in2 => \N__45396\,
            in3 => \N__45387\,
            lcout => \ADC_VDC.genclk.n21444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48989\,
            in1 => \N__48902\,
            in2 => \N__48120\,
            in3 => \N__48158\,
            lcout => \ADC_VDC.genclk.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48173\,
            in1 => \N__48920\,
            in2 => \N__49008\,
            in3 => \N__48953\,
            lcout => \ADC_VDC.genclk.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_adj_8_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48935\,
            in1 => \N__49212\,
            in2 => \N__48974\,
            in3 => \N__48887\,
            lcout => \ADC_VDC.genclk.n28_adj_1397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_93_2_lut_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45259\,
            in2 => \_gnd_net_\,
            in3 => \N__55778\,
            lcout => \comm_spi.data_tx_7__N_767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_6_i1_3_lut_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45338\,
            in1 => \N__47878\,
            in2 => \_gnd_net_\,
            in3 => \N__50793\,
            lcout => OPEN,
            ltout => \n1_adj_1588_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i6_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__50604\,
            in1 => \N__45105\,
            in2 => \N__45273\,
            in3 => \N__45570\,
            lcout => comm_tx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54324\,
            ce => \N__45233\,
            sr => \N__45177\
        );

    \mux_137_Mux_6_i2_3_lut_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45474\,
            in1 => \N__45114\,
            in2 => \_gnd_net_\,
            in3 => \N__50792\,
            lcout => n2_adj_1589,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19276_2_lut_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45600\,
            in2 => \_gnd_net_\,
            in3 => \N__50791\,
            lcout => OPEN,
            ltout => \n21539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19724_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__50603\,
            in1 => \N__45579\,
            in2 => \N__45573\,
            in3 => \N__52411\,
            lcout => n22339,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i0_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45564\,
            in1 => \N__51950\,
            in2 => \_gnd_net_\,
            in3 => \N__53035\,
            lcout => comm_buf_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \comm_buf_3__i4_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51948\,
            in1 => \N__46772\,
            in2 => \_gnd_net_\,
            in3 => \N__45546\,
            lcout => comm_buf_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \comm_buf_3__i7_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50409\,
            in1 => \N__45519\,
            in2 => \_gnd_net_\,
            in3 => \N__51945\,
            lcout => comm_buf_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \comm_buf_3__i6_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51949\,
            in1 => \N__46461\,
            in2 => \_gnd_net_\,
            in3 => \N__45489\,
            lcout => comm_buf_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \comm_buf_3__i5_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52112\,
            in1 => \N__45465\,
            in2 => \_gnd_net_\,
            in3 => \N__51944\,
            lcout => comm_buf_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \comm_buf_3__i3_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51947\,
            in1 => \N__51108\,
            in2 => \_gnd_net_\,
            in3 => \N__45444\,
            lcout => comm_buf_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \comm_buf_3__i2_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47236\,
            in1 => \N__45420\,
            in2 => \_gnd_net_\,
            in3 => \N__51943\,
            lcout => comm_buf_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \comm_buf_3__i1_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51946\,
            in1 => \N__45795\,
            in2 => \_gnd_net_\,
            in3 => \N__45696\,
            lcout => comm_buf_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54336\,
            ce => \N__45651\,
            sr => \N__45642\
        );

    \i2_3_lut_adj_78_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__49793\,
            in1 => \N__49748\,
            in2 => \_gnd_net_\,
            in3 => \N__49712\,
            lcout => n20878,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19274_2_lut_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45631\,
            in2 => \_gnd_net_\,
            in3 => \N__49800\,
            lcout => OPEN,
            ltout => \n21352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011010101"
        )
    port map (
            in0 => \N__51924\,
            in1 => \N__50752\,
            in2 => \N__45657\,
            in3 => \N__45954\,
            lcout => OPEN,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_272_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45915\,
            in2 => \N__45654\,
            in3 => \N__45880\,
            lcout => n12136,
            ltout => \n12136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12358_2_lut_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45645\,
            in3 => \N__56867\,
            lcout => n14771,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_50_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__50026\,
            in1 => \N__52388\,
            in2 => \N__49877\,
            in3 => \N__52243\,
            lcout => n18991,
            ltout => \n18991_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_265_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__45632\,
            in1 => \N__50751\,
            in2 => \N__45606\,
            in3 => \N__51999\,
            lcout => OPEN,
            ltout => \n4_adj_1545_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_266_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__49665\,
            in1 => \N__45914\,
            in2 => \N__45603\,
            in3 => \N__45879\,
            lcout => n11961,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_47_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__50584\,
            in1 => \N__49503\,
            in2 => \_gnd_net_\,
            in3 => \N__49292\,
            lcout => n18993,
            ltout => \n18993_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_276_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001010101"
        )
    port map (
            in0 => \N__45953\,
            in1 => \N__50786\,
            in2 => \N__46095\,
            in3 => \N__51917\,
            lcout => n12_adj_1605,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_269_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__45876\,
            in1 => \_gnd_net_\,
            in2 => \N__45920\,
            in3 => \N__49236\,
            lcout => n11991,
            ltout => \n11991_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12344_2_lut_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__57066\,
            in1 => \_gnd_net_\,
            in2 => \N__46086\,
            in3 => \_gnd_net_\,
            lcout => n14757,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_48_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__49587\,
            in1 => \N__55408\,
            in2 => \_gnd_net_\,
            in3 => \N__57065\,
            lcout => n20843,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i7_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__46083\,
            in1 => \N__52254\,
            in2 => \N__50412\,
            in3 => \N__46014\,
            lcout => comm_cmd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_273_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__51916\,
            in1 => \N__45952\,
            in2 => \N__50798\,
            in3 => \N__45933\,
            lcout => OPEN,
            ltout => \n12_adj_1635_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_274_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45910\,
            in2 => \N__45885\,
            in3 => \N__45877\,
            lcout => n12178,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19639_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__54757\,
            in1 => \N__53611\,
            in2 => \N__46557\,
            in3 => \N__46470\,
            lcout => OPEN,
            ltout => \n22225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22225_bdd_4_lut_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__47007\,
            in1 => \N__46287\,
            in2 => \N__46539\,
            in3 => \N__54758\,
            lcout => n22228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_6_i26_3_lut_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46536\,
            in1 => \N__57805\,
            in2 => \_gnd_net_\,
            in3 => \N__46515\,
            lcout => OPEN,
            ltout => \n26_adj_1507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18568_4_lut_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__57807\,
            in1 => \N__46485\,
            in2 => \N__46473\,
            in3 => \N__55153\,
            lcout => n21178,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i6_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51860\,
            in1 => \N__46463\,
            in2 => \_gnd_net_\,
            in3 => \N__46383\,
            lcout => comm_buf_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54377\,
            ce => \N__51356\,
            sr => \N__51257\
        );

    \mux_129_Mux_6_i19_3_lut_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57806\,
            in1 => \N__46377\,
            in2 => \_gnd_net_\,
            in3 => \N__46349\,
            lcout => OPEN,
            ltout => \n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18436_3_lut_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55154\,
            in1 => \_gnd_net_\,
            in2 => \N__46320\,
            in3 => \N__46317\,
            lcout => n21046,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22231_bdd_4_lut_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__53791\,
            in1 => \N__46281\,
            in2 => \N__46269\,
            in3 => \N__46230\,
            lcout => n22234,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i26_3_lut_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46218\,
            in1 => \N__57817\,
            in2 => \_gnd_net_\,
            in3 => \N__46197\,
            lcout => OPEN,
            ltout => \n26_adj_1512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19714_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__53883\,
            in1 => \N__55157\,
            in2 => \N__46854\,
            in3 => \N__53792\,
            lcout => OPEN,
            ltout => \n22351_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22351_bdd_4_lut_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__53793\,
            in1 => \N__46851\,
            in2 => \N__46824\,
            in3 => \N__46821\,
            lcout => OPEN,
            ltout => \n22354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1555570_i1_3_lut_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46797\,
            in2 => \N__46791\,
            in3 => \N__54744\,
            lcout => OPEN,
            ltout => \n30_adj_1513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i4_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__46788\,
            in1 => \_gnd_net_\,
            in2 => \N__46689\,
            in3 => \N__52008\,
            lcout => comm_buf_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54391\,
            ce => \N__51384\,
            sr => \N__51283\
        );

    \comm_cmd_1__bdd_4_lut_19598_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__46686\,
            in1 => \N__55155\,
            in2 => \N__46674\,
            in3 => \N__53787\,
            lcout => OPEN,
            ltout => \n22207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22207_bdd_4_lut_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__53788\,
            in1 => \N__46640\,
            in2 => \N__46617\,
            in3 => \N__46863\,
            lcout => n22210,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__55156\,
            in1 => \N__47103\,
            in2 => \N__52722\,
            in3 => \N__53789\,
            lcout => OPEN,
            ltout => \n22429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22429_bdd_4_lut_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__53790\,
            in1 => \N__46614\,
            in2 => \N__46587\,
            in3 => \N__46584\,
            lcout => OPEN,
            ltout => \n22432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1554364_i1_3_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47253\,
            in2 => \N__47247\,
            in3 => \N__54764\,
            lcout => OPEN,
            ltout => \n30_adj_1520_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i2_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__51998\,
            in1 => \N__47243\,
            in2 => \N__47151\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54403\,
            ce => \N__51374\,
            sr => \N__51300\
        );

    \mux_129_Mux_2_i26_3_lut_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__47148\,
            in1 => \_gnd_net_\,
            in2 => \N__57819\,
            in3 => \N__47127\,
            lcout => n26_adj_1519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15326_2_lut_3_lut_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__50999\,
            in1 => \N__55480\,
            in2 => \_gnd_net_\,
            in3 => \N__52027\,
            lcout => n14_adj_1585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_368_i8_2_lut_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55148\,
            in2 => \_gnd_net_\,
            in3 => \N__53766\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18435_3_lut_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47039\,
            in1 => \N__47016\,
            in2 => \_gnd_net_\,
            in3 => \N__55150\,
            lcout => n21045,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18444_3_lut_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55149\,
            in1 => \N__46998\,
            in2 => \_gnd_net_\,
            in3 => \N__46977\,
            lcout => n21054,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_3_i16_3_lut_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57763\,
            in2 => \N__46952\,
            in3 => \N__46916\,
            lcout => n16_adj_1514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i16_3_lut_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46892\,
            in1 => \N__47914\,
            in2 => \_gnd_net_\,
            in3 => \N__57824\,
            lcout => n16_adj_1517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i2_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__47915\,
            in1 => \N__56451\,
            in2 => \N__48067\,
            in3 => \N__48011\,
            lcout => buf_dds0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15342_2_lut_3_lut_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__47891\,
            in1 => \N__51997\,
            in2 => \_gnd_net_\,
            in3 => \N__55541\,
            lcout => n14_adj_1552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6419_3_lut_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47763\,
            in1 => \N__47727\,
            in2 => \_gnd_net_\,
            in3 => \N__47701\,
            lcout => n8_adj_1567,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__57138\,
            in1 => \N__47633\,
            in2 => \N__56477\,
            in3 => \N__47621\,
            lcout => \data_index_9_N_216_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19407_2_lut_4_lut_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011111111111"
        )
    port map (
            in0 => \N__58010\,
            in1 => \N__53351\,
            in2 => \N__58160\,
            in3 => \N__52908\,
            lcout => \ADC_VDC.genclk.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19334_2_lut_LC_19_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52907\,
            in2 => \_gnd_net_\,
            in3 => \N__58006\,
            lcout => \ADC_VDC.genclk.n11735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16159_4_lut_LC_19_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100010111010"
        )
    port map (
            in0 => \N__48786\,
            in1 => \N__48581\,
            in2 => \N__47262\,
            in3 => \N__48356\,
            lcout => \ADC_VDC.n11750\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_LC_19_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47493\,
            in2 => \_gnd_net_\,
            in3 => \N__47363\,
            lcout => \ADC_VDC.n62\,
            ltout => \ADC_VDC.n62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i24_4_lut_LC_19_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100010111010"
        )
    port map (
            in0 => \N__48785\,
            in1 => \N__48580\,
            in2 => \N__48360\,
            in3 => \N__48355\,
            lcout => \ADC_VDC.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12196_12197_set_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52971\,
            in1 => \N__52948\,
            in2 => \_gnd_net_\,
            in3 => \N__55902\,
            lcout => \comm_spi.n14614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52570\,
            ce => 'H',
            sr => \N__52920\
        );

    \ADC_VDC.genclk.t0off_i0_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48207\,
            in2 => \_gnd_net_\,
            in3 => \N__48195\,
            lcout => \ADC_VDC.genclk.t0off_0\,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => \ADC_VDC.genclk.n19709\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i1_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48192\,
            in2 => \N__58522\,
            in3 => \N__48180\,
            lcout => \ADC_VDC.genclk.t0off_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19709\,
            carryout => \ADC_VDC.genclk.n19710\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i2_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58447\,
            in2 => \N__48177\,
            in3 => \N__48162\,
            lcout => \ADC_VDC.genclk.t0off_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19710\,
            carryout => \ADC_VDC.genclk.n19711\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i3_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48159\,
            in2 => \N__58523\,
            in3 => \N__48147\,
            lcout => \ADC_VDC.genclk.t0off_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19711\,
            carryout => \ADC_VDC.genclk.n19712\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i4_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58451\,
            in2 => \N__48143\,
            in3 => \N__48123\,
            lcout => \ADC_VDC.genclk.t0off_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19712\,
            carryout => \ADC_VDC.genclk.n19713\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i5_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48119\,
            in2 => \N__58524\,
            in3 => \N__48105\,
            lcout => \ADC_VDC.genclk.t0off_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19713\,
            carryout => \ADC_VDC.genclk.n19714\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i6_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58455\,
            in2 => \N__48102\,
            in3 => \N__48087\,
            lcout => \ADC_VDC.genclk.t0off_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19714\,
            carryout => \ADC_VDC.genclk.n19715\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i7_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49007\,
            in2 => \N__58525\,
            in3 => \N__48993\,
            lcout => \ADC_VDC.genclk.t0off_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19715\,
            carryout => \ADC_VDC.genclk.n19716\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__49197\,
            sr => \N__58243\
        );

    \ADC_VDC.genclk.t0off_i8_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48990\,
            in2 => \N__58576\,
            in3 => \N__48978\,
            lcout => \ADC_VDC.genclk.t0off_8\,
            ltout => OPEN,
            carryin => \bfn_19_8_0_\,
            carryout => \ADC_VDC.genclk.n19717\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \ADC_VDC.genclk.t0off_i9_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58541\,
            in2 => \N__48975\,
            in3 => \N__48957\,
            lcout => \ADC_VDC.genclk.t0off_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19717\,
            carryout => \ADC_VDC.genclk.n19718\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \ADC_VDC.genclk.t0off_i10_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48954\,
            in2 => \N__58573\,
            in3 => \N__48942\,
            lcout => \ADC_VDC.genclk.t0off_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19718\,
            carryout => \ADC_VDC.genclk.n19719\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \ADC_VDC.genclk.t0off_i11_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58529\,
            in2 => \N__48939\,
            in3 => \N__48924\,
            lcout => \ADC_VDC.genclk.t0off_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19719\,
            carryout => \ADC_VDC.genclk.n19720\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \ADC_VDC.genclk.t0off_i12_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48921\,
            in2 => \N__58574\,
            in3 => \N__48909\,
            lcout => \ADC_VDC.genclk.t0off_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19720\,
            carryout => \ADC_VDC.genclk.n19721\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \ADC_VDC.genclk.t0off_i13_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58533\,
            in2 => \N__48906\,
            in3 => \N__48891\,
            lcout => \ADC_VDC.genclk.t0off_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19721\,
            carryout => \ADC_VDC.genclk.n19722\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \ADC_VDC.genclk.t0off_i14_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48888\,
            in2 => \N__58575\,
            in3 => \N__48876\,
            lcout => \ADC_VDC.genclk.t0off_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19722\,
            carryout => \ADC_VDC.genclk.n19723\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \ADC_VDC.genclk.t0off_i15_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49211\,
            in1 => \N__58537\,
            in2 => \_gnd_net_\,
            in3 => \N__49215\,
            lcout => \ADC_VDC.genclk.t0off_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__49196\,
            sr => \N__58263\
        );

    \comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__55350\,
            in1 => \N__49017\,
            in2 => \N__49026\,
            in3 => \N__49176\,
            lcout => n17815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000000000"
        )
    port map (
            in0 => \N__51724\,
            in1 => \N__55351\,
            in2 => \N__50046\,
            in3 => \N__49881\,
            lcout => OPEN,
            ltout => \n21_adj_1598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19391_4_lut_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101111111111"
        )
    port map (
            in0 => \N__55352\,
            in1 => \N__49128\,
            in2 => \N__49113\,
            in3 => \N__49110\,
            lcout => n18_adj_1619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i32_4_lut_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__51725\,
            in1 => \N__55353\,
            in2 => \N__49674\,
            in3 => \N__49092\,
            lcout => OPEN,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i2_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__50058\,
            in1 => \N__49050\,
            in2 => \N__49035\,
            in3 => \N__49464\,
            lcout => comm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54350\,
            ce => \N__49032\,
            sr => \N__57118\
        );

    \i11712_2_lut_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49494\,
            in3 => \N__51721\,
            lcout => n14130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_318_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111011"
        )
    port map (
            in0 => \N__52428\,
            in1 => \N__51723\,
            in2 => \N__54459\,
            in3 => \N__52410\,
            lcout => n20880,
            ltout => \n20880_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i33_3_lut_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49463\,
            in1 => \_gnd_net_\,
            in2 => \N__49011\,
            in3 => \N__51722\,
            lcout => n12_adj_1548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__52409\,
            in1 => \N__52244\,
            in2 => \N__50051\,
            in3 => \N__49867\,
            lcout => n18984,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19308_2_lut_3_lut_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__49794\,
            in1 => \N__49749\,
            in2 => \_gnd_net_\,
            in3 => \N__49713\,
            lcout => n21546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__55348\,
            in1 => \N__56852\,
            in2 => \N__51995\,
            in3 => \N__49279\,
            lcout => n12092,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_281_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011101"
        )
    port map (
            in0 => \N__55349\,
            in1 => \N__56853\,
            in2 => \N__51996\,
            in3 => \N__49281\,
            lcout => OPEN,
            ltout => \n11853_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_121_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__49656\,
            in1 => \N__49623\,
            in2 => \N__49605\,
            in3 => \N__49585\,
            lcout => n11860,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19318_3_lut_4_lut_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__50602\,
            in1 => \N__49492\,
            in2 => \N__50799\,
            in3 => \N__49293\,
            lcout => OPEN,
            ltout => \n21339_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i42_4_lut_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__49280\,
            in1 => \N__49254\,
            in2 => \N__49239\,
            in3 => \N__51909\,
            lcout => n38_adj_1608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19674_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__54759\,
            in1 => \N__53767\,
            in2 => \N__49230\,
            in3 => \N__50418\,
            lcout => OPEN,
            ltout => \n22267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22267_bdd_4_lut_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__50160\,
            in1 => \N__52134\,
            in2 => \N__50481\,
            in3 => \N__54760\,
            lcout => n22270,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i26_3_lut_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50478\,
            in1 => \N__50457\,
            in2 => \_gnd_net_\,
            in3 => \N__57651\,
            lcout => OPEN,
            ltout => \n26_adj_1502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18445_4_lut_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__57653\,
            in1 => \N__50433\,
            in2 => \N__50421\,
            in3 => \N__55233\,
            lcout => n21055,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i7_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50408\,
            in1 => \N__52007\,
            in2 => \_gnd_net_\,
            in3 => \N__50328\,
            lcout => comm_buf_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54378\,
            ce => \N__51357\,
            sr => \N__51306\
        );

    \mux_129_Mux_7_i19_3_lut_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57652\,
            in1 => \N__50238\,
            in2 => \_gnd_net_\,
            in3 => \N__50216\,
            lcout => OPEN,
            ltout => \n19_adj_1503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18439_3_lut_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55234\,
            in1 => \_gnd_net_\,
            in2 => \N__50187\,
            in3 => \N__50184\,
            lcout => n21049,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18517_3_lut_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__50154\,
            in1 => \N__50889\,
            in2 => \N__55212\,
            in3 => \_gnd_net_\,
            lcout => n21127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18522_3_lut_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50124\,
            in1 => \N__55145\,
            in2 => \_gnd_net_\,
            in3 => \N__50088\,
            lcout => OPEN,
            ltout => \n21132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19788_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__54761\,
            in1 => \N__53612\,
            in2 => \N__51126\,
            in3 => \N__50817\,
            lcout => OPEN,
            ltout => \n22333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22333_bdd_4_lut_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__52746\,
            in1 => \N__51123\,
            in2 => \N__51117\,
            in3 => \N__54762\,
            lcout => OPEN,
            ltout => \n22336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i3_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51109\,
            in2 => \N__51024\,
            in3 => \N__51925\,
            lcout => comm_buf_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54392\,
            ce => \N__51358\,
            sr => \N__51299\
        );

    \mux_129_Mux_3_i19_3_lut_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57812\,
            in1 => \N__50949\,
            in2 => \_gnd_net_\,
            in3 => \N__50922\,
            lcout => n19_adj_1515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_3_i26_3_lut_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50883\,
            in1 => \N__57813\,
            in2 => \_gnd_net_\,
            in3 => \N__50861\,
            lcout => OPEN,
            ltout => \n26_adj_1516_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18523_4_lut_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__57814\,
            in1 => \N__50835\,
            in2 => \N__50820\,
            in3 => \N__55141\,
            lcout => n21133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19098_4_lut_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__57089\,
            in1 => \N__54653\,
            in2 => \N__52197\,
            in3 => \N__53794\,
            lcout => OPEN,
            ltout => \n21316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i2_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__53924\,
            in1 => \N__50808\,
            in2 => \N__50811\,
            in3 => \N__57754\,
            lcout => comm_length_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_315_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__50807\,
            in1 => \N__50782\,
            in2 => \N__55248\,
            in3 => \N__50601\,
            lcout => n4_adj_1600,
            ltout => \n4_adj_1600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_319_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54449\,
            in2 => \N__52416\,
            in3 => \N__52412\,
            lcout => OPEN,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19278_3_lut_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52000\,
            in2 => \N__52269\,
            in3 => \N__52258\,
            lcout => n21888,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19194_2_lut_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55421\,
            lcout => n21317,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18438_3_lut_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52187\,
            in1 => \N__52146\,
            in2 => \_gnd_net_\,
            in3 => \N__55230\,
            lcout => n21048,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i5_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__52124\,
            in1 => \N__52028\,
            in2 => \_gnd_net_\,
            in3 => \N__52794\,
            lcout => comm_buf_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54417\,
            ce => \N__51382\,
            sr => \N__51301\
        );

    \comm_cmd_1__bdd_4_lut_19759_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__51228\,
            in1 => \N__55218\,
            in2 => \N__51210\,
            in3 => \N__53782\,
            lcout => n22399,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i26_3_lut_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__51177\,
            in1 => \N__57750\,
            in2 => \_gnd_net_\,
            in3 => \N__51156\,
            lcout => OPEN,
            ltout => \n26_adj_1498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19709_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__57837\,
            in1 => \N__55219\,
            in2 => \N__51129\,
            in3 => \N__53783\,
            lcout => OPEN,
            ltout => \n22345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22345_bdd_4_lut_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__53784\,
            in1 => \N__52851\,
            in2 => \N__52824\,
            in3 => \N__52821\,
            lcout => OPEN,
            ltout => \n22348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1556776_i1_3_lut_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53358\,
            in2 => \N__52797\,
            in3 => \N__54763\,
            lcout => n30_adj_1500,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18516_3_lut_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52787\,
            in1 => \N__52752\,
            in2 => \_gnd_net_\,
            in3 => \N__55232\,
            lcout => n21126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19322_2_lut_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52734\,
            in2 => \_gnd_net_\,
            in3 => \N__57749\,
            lcout => n21564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18970_2_lut_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52707\,
            in2 => \_gnd_net_\,
            in3 => \N__57748\,
            lcout => n21218,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19053_2_lut_LC_20_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__52680\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57820\,
            lcout => n21364,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i1_LC_20_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52906\,
            in2 => \_gnd_net_\,
            in3 => \N__58002\,
            lcout => \ADC_VDC.genclk.div_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i1C_net\,
            ce => \N__52650\,
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12196_12197_reset_LC_20_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55901\,
            in1 => \N__52950\,
            in2 => \_gnd_net_\,
            in3 => \N__52970\,
            lcout => \comm_spi.n14615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52627\,
            ce => 'H',
            sr => \N__53334\
        );

    \ADC_VDC.genclk.div_state_i0_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__58005\,
            in1 => \N__53352\,
            in2 => \N__58161\,
            in3 => \N__52894\,
            lcout => \ADC_VDC.genclk.div_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_87_2_lut_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55765\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52875\,
            lcout => \comm_spi.DOUT_7__N_747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t_clk_24_LC_20_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__58004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VDC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12198_3_lut_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53067\,
            in1 => \N__53061\,
            in2 => \_gnd_net_\,
            in3 => \N__52862\,
            lcout => comm_rx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19420_4_lut_3_lut_LC_20_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55614\,
            in1 => \N__52969\,
            in2 => \_gnd_net_\,
            in3 => \N__55763\,
            lcout => \comm_spi.n22866\,
            ltout => \comm_spi.n22866_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12184_3_lut_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55900\,
            in2 => \N__52953\,
            in3 => \N__52949\,
            lcout => \comm_spi.imosi\,
            ltout => \comm_spi.imosi_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_86_2_lut_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52923\,
            in3 => \N__55764\,
            lcout => \comm_spi.DOUT_7__N_746\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12646_2_lut_2_lut_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__52893\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58003\,
            lcout => \ADC_VDC.genclk.n15051\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19435_4_lut_3_lut_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52863\,
            in1 => \N__55868\,
            in2 => \_gnd_net_\,
            in3 => \N__52874\,
            lcout => \comm_spi.n22863\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_12182_12183_set_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55636\,
            lcout => \comm_spi.n14600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54365\,
            ce => 'H',
            sr => \N__55572\
        );

    \comm_spi.RESET_I_0_88_2_lut_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55638\,
            lcout => \comm_spi.imosi_N_752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12237_3_lut_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__53917\,
            in1 => \N__55422\,
            in2 => \_gnd_net_\,
            in3 => \N__57000\,
            lcout => n14655,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i0_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010111000110"
        )
    port map (
            in0 => \N__54711\,
            in1 => \N__55235\,
            in2 => \N__57825\,
            in3 => \N__53614\,
            lcout => comm_length_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54405\,
            ce => \N__53925\,
            sr => \N__53901\
        );

    \comm_length_i1_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111011001111"
        )
    port map (
            in0 => \N__53613\,
            in1 => \N__57808\,
            in2 => \N__55239\,
            in3 => \N__54712\,
            lcout => comm_length_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__54405\,
            ce => \N__53925\,
            sr => \N__53901\
        );

    \i19319_2_lut_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__57779\,
            in1 => \_gnd_net_\,
            in2 => \N__53895\,
            in3 => \_gnd_net_\,
            lcout => n21451,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18978_2_lut_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53874\,
            in2 => \_gnd_net_\,
            in3 => \N__57778\,
            lcout => n21151,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22399_bdd_4_lut_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__53850\,
            in1 => \N__53838\,
            in2 => \N__53831\,
            in3 => \N__53785\,
            lcout => n22402,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19119_2_lut_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__57843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57780\,
            lcout => n21350,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19283_2_lut_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57831\,
            in2 => \_gnd_net_\,
            in3 => \N__57818\,
            lcout => n21529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15092_4_lut_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__56999\,
            in1 => \N__56594\,
            in2 => \N__56518\,
            in3 => \N__56031\,
            lcout => \data_index_9_N_216_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0on_i0_LC_22_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58176\,
            in2 => \_gnd_net_\,
            in3 => \N__55917\,
            lcout => \ADC_VDC.genclk.t0on_0\,
            ltout => OPEN,
            carryin => \bfn_22_7_0_\,
            carryout => \ADC_VDC.genclk.n19724\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i1_LC_22_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58206\,
            in2 => \N__58577\,
            in3 => \N__55914\,
            lcout => \ADC_VDC.genclk.t0on_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19724\,
            carryout => \ADC_VDC.genclk.n19725\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i2_LC_22_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58545\,
            in2 => \N__58119\,
            in3 => \N__55911\,
            lcout => \ADC_VDC.genclk.t0on_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19725\,
            carryout => \ADC_VDC.genclk.n19726\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i3_LC_22_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58071\,
            in2 => \N__58578\,
            in3 => \N__55908\,
            lcout => \ADC_VDC.genclk.t0on_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19726\,
            carryout => \ADC_VDC.genclk.n19727\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i4_LC_22_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58549\,
            in2 => \N__58194\,
            in3 => \N__55905\,
            lcout => \ADC_VDC.genclk.t0on_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19727\,
            carryout => \ADC_VDC.genclk.n19728\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i5_LC_22_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58043\,
            in2 => \N__58579\,
            in3 => \N__57870\,
            lcout => \ADC_VDC.genclk.t0on_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19728\,
            carryout => \ADC_VDC.genclk.n19729\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i6_LC_22_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58553\,
            in2 => \N__58221\,
            in3 => \N__57867\,
            lcout => \ADC_VDC.genclk.t0on_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19729\,
            carryout => \ADC_VDC.genclk.n19730\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i7_LC_22_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58103\,
            in2 => \N__58580\,
            in3 => \N__57864\,
            lcout => \ADC_VDC.genclk.t0on_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19730\,
            carryout => \ADC_VDC.genclk.n19731\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57959\,
            sr => \N__58259\
        );

    \ADC_VDC.genclk.t0on_i8_LC_22_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58029\,
            in2 => \N__58503\,
            in3 => \N__57861\,
            lcout => \ADC_VDC.genclk.t0on_8\,
            ltout => OPEN,
            carryin => \bfn_22_8_0_\,
            carryout => \ADC_VDC.genclk.n19732\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.t0on_i9_LC_22_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58420\,
            in2 => \N__57924\,
            in3 => \N__57858\,
            lcout => \ADC_VDC.genclk.t0on_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19732\,
            carryout => \ADC_VDC.genclk.n19733\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.t0on_i10_LC_22_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58089\,
            in2 => \N__58500\,
            in3 => \N__57855\,
            lcout => \ADC_VDC.genclk.t0on_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19733\,
            carryout => \ADC_VDC.genclk.n19734\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.t0on_i11_LC_22_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58408\,
            in2 => \N__57894\,
            in3 => \N__57852\,
            lcout => \ADC_VDC.genclk.t0on_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19734\,
            carryout => \ADC_VDC.genclk.n19735\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.t0on_i12_LC_22_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58131\,
            in2 => \N__58501\,
            in3 => \N__57849\,
            lcout => \ADC_VDC.genclk.t0on_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19735\,
            carryout => \ADC_VDC.genclk.n19736\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.t0on_i13_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58412\,
            in2 => \N__58059\,
            in3 => \N__57846\,
            lcout => \ADC_VDC.genclk.t0on_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19736\,
            carryout => \ADC_VDC.genclk.n19737\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.t0on_i14_LC_22_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57936\,
            in2 => \N__58502\,
            in3 => \N__58626\,
            lcout => \ADC_VDC.genclk.t0on_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19737\,
            carryout => \ADC_VDC.genclk.n19738\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.t0on_i15_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57908\,
            in1 => \N__58416\,
            in2 => \_gnd_net_\,
            in3 => \N__58266\,
            lcout => \ADC_VDC.genclk.t0on_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57963\,
            sr => \N__58258\
        );

    \ADC_VDC.genclk.i19049_4_lut_LC_23_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__58217\,
            in1 => \N__58205\,
            in2 => \N__58193\,
            in3 => \N__58175\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n21449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19183_4_lut_LC_23_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57879\,
            in1 => \N__58017\,
            in2 => \N__58164\,
            in3 => \N__58077\,
            lcout => \ADC_VDC.genclk.n21443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_adj_7_LC_23_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__58130\,
            in1 => \N__58115\,
            in2 => \N__58104\,
            in3 => \N__58088\,
            lcout => \ADC_VDC.genclk.n27_adj_1396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_adj_6_LC_23_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__58070\,
            in1 => \N__58055\,
            in2 => \N__58044\,
            in3 => \N__58028\,
            lcout => \ADC_VDC.genclk.n26_adj_1395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_23_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58011\,
            lcout => \ADC_VDC.genclk.div_state_1__N_1274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_LC_23_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57935\,
            in1 => \N__57920\,
            in2 => \N__57909\,
            in3 => \N__57890\,
            lcout => \ADC_VDC.genclk.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
